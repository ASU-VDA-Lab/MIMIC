module real_aes_8038_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g546 ( .A1(n_0), .A2(n_177), .B(n_547), .C(n_550), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_1), .B(n_497), .Y(n_551) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g189 ( .A(n_3), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_4), .B(n_149), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_5), .A2(n_105), .B1(n_118), .B2(n_767), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_6), .A2(n_470), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_7), .A2(n_169), .B(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_8), .A2(n_39), .B1(n_143), .B2(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_9), .B(n_169), .Y(n_178) );
AND2x6_ASAP7_75t_L g161 ( .A(n_10), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_11), .A2(n_161), .B(n_475), .C(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_12), .B(n_40), .Y(n_117) );
INVx1_ASAP7_75t_L g139 ( .A(n_13), .Y(n_139) );
INVx1_ASAP7_75t_L g182 ( .A(n_14), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_15), .B(n_147), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_16), .B(n_149), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_17), .B(n_135), .Y(n_253) );
AO32x2_ASAP7_75t_L g195 ( .A1(n_18), .A2(n_134), .A3(n_160), .B1(n_169), .B2(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_19), .B(n_143), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_20), .B(n_135), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_21), .A2(n_55), .B1(n_143), .B2(n_198), .Y(n_199) );
AOI22xp33_ASAP7_75t_SL g237 ( .A1(n_22), .A2(n_82), .B1(n_143), .B2(n_147), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_23), .B(n_143), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_24), .A2(n_160), .B(n_475), .C(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_25), .A2(n_61), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_25), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_26), .A2(n_160), .B(n_475), .C(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_27), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_28), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_29), .B(n_439), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_30), .A2(n_470), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_31), .B(n_164), .Y(n_212) );
INVx2_ASAP7_75t_L g145 ( .A(n_32), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_33), .A2(n_473), .B(n_483), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_34), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_35), .B(n_164), .Y(n_223) );
XNOR2x2_ASAP7_75t_SL g122 ( .A(n_36), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_37), .B(n_219), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_38), .A2(n_86), .B1(n_452), .B2(n_453), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_38), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_41), .B(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_42), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_43), .B(n_149), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_44), .B(n_470), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_45), .A2(n_473), .B(n_477), .C(n_483), .Y(n_472) );
OAI321xp33_ASAP7_75t_L g121 ( .A1(n_46), .A2(n_122), .A3(n_431), .B1(n_435), .B2(n_436), .C(n_438), .Y(n_121) );
INVx1_ASAP7_75t_L g435 ( .A(n_46), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_47), .B(n_143), .Y(n_172) );
INVx1_ASAP7_75t_L g548 ( .A(n_48), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_49), .A2(n_92), .B1(n_198), .B2(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g478 ( .A(n_50), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_51), .B(n_143), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_52), .B(n_143), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_53), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_54), .B(n_155), .Y(n_176) );
AOI22xp33_ASAP7_75t_SL g251 ( .A1(n_56), .A2(n_62), .B1(n_143), .B2(n_147), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_57), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_58), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_59), .B(n_143), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_60), .B(n_143), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_61), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_61), .A2(n_126), .B1(n_127), .B2(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g162 ( .A(n_63), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_64), .B(n_470), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_65), .B(n_497), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_66), .A2(n_155), .B(n_185), .C(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_67), .B(n_143), .Y(n_190) );
INVx1_ASAP7_75t_L g138 ( .A(n_68), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_69), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_70), .B(n_149), .Y(n_515) );
AO32x2_ASAP7_75t_L g233 ( .A1(n_71), .A2(n_160), .A3(n_169), .B1(n_234), .B2(n_238), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_72), .B(n_150), .Y(n_561) );
INVx1_ASAP7_75t_L g153 ( .A(n_73), .Y(n_153) );
INVx1_ASAP7_75t_L g207 ( .A(n_74), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_75), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_76), .B(n_480), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_77), .A2(n_475), .B(n_483), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_78), .B(n_147), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_79), .Y(n_492) );
INVx1_ASAP7_75t_L g110 ( .A(n_80), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_81), .B(n_479), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_83), .B(n_198), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_84), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_85), .B(n_147), .Y(n_211) );
INVx1_ASAP7_75t_L g453 ( .A(n_86), .Y(n_453) );
INVx2_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_88), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_89), .B(n_159), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_90), .B(n_147), .Y(n_173) );
INVx2_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
OR2x2_ASAP7_75t_L g434 ( .A(n_91), .B(n_114), .Y(n_434) );
OR2x2_ASAP7_75t_L g457 ( .A(n_91), .B(n_115), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_93), .A2(n_103), .B1(n_147), .B2(n_148), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_94), .B(n_470), .Y(n_511) );
INVx1_ASAP7_75t_L g514 ( .A(n_95), .Y(n_514) );
INVxp67_ASAP7_75t_L g495 ( .A(n_96), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_97), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g536 ( .A(n_99), .Y(n_536) );
INVx1_ASAP7_75t_L g557 ( .A(n_100), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_101), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_101), .Y(n_449) );
AND2x2_ASAP7_75t_L g485 ( .A(n_102), .B(n_164), .Y(n_485) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_108), .Y(n_767) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_SL g766 ( .A(n_109), .Y(n_766) );
INVx1_ASAP7_75t_SL g445 ( .A(n_111), .Y(n_445) );
INVx3_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
NOR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OR2x2_ASAP7_75t_L g462 ( .A(n_113), .B(n_115), .Y(n_462) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OA211x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_121), .B(n_442), .C(n_766), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g443 ( .A(n_120), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_122), .B(n_437), .Y(n_436) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
INVx1_ASAP7_75t_SL g459 ( .A(n_127), .Y(n_459) );
OR3x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_359), .C(n_408), .Y(n_127) );
NAND5xp2_ASAP7_75t_L g128 ( .A(n_129), .B(n_274), .C(n_302), .D(n_332), .E(n_346), .Y(n_128) );
AOI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_192), .B1(n_224), .B2(n_229), .C(n_240), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_165), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_131), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g254 ( .A(n_132), .Y(n_254) );
AND2x2_ASAP7_75t_L g262 ( .A(n_132), .B(n_168), .Y(n_262) );
AND2x2_ASAP7_75t_L g285 ( .A(n_132), .B(n_167), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_132), .B(n_179), .Y(n_300) );
OR2x2_ASAP7_75t_L g309 ( .A(n_132), .B(n_247), .Y(n_309) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_132), .Y(n_312) );
AND2x2_ASAP7_75t_L g420 ( .A(n_132), .B(n_247), .Y(n_420) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_163), .Y(n_132) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_133), .A2(n_180), .B(n_191), .Y(n_179) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_134), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_136), .B(n_137), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_152), .B(n_160), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B(n_149), .Y(n_141) );
INVx3_ASAP7_75t_L g206 ( .A(n_143), .Y(n_206) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_143), .Y(n_538) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g198 ( .A(n_144), .Y(n_198) );
BUFx3_ASAP7_75t_L g236 ( .A(n_144), .Y(n_236) );
AND2x6_ASAP7_75t_L g475 ( .A(n_144), .B(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
INVx1_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx2_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_149), .A2(n_172), .B(n_173), .Y(n_171) );
INVx2_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
O2A1O1Ixp5_ASAP7_75t_SL g205 ( .A1(n_149), .A2(n_206), .B(n_207), .C(n_208), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_149), .B(n_495), .Y(n_494) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g234 ( .A1(n_150), .A2(n_159), .B1(n_235), .B2(n_237), .Y(n_234) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVx1_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
AND2x2_ASAP7_75t_L g471 ( .A(n_151), .B(n_156), .Y(n_471) );
INVx1_ASAP7_75t_L g476 ( .A(n_151), .Y(n_476) );
O2A1O1Ixp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .C(n_158), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_154), .A2(n_177), .B(n_189), .C(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_154), .A2(n_525), .B(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_158), .A2(n_221), .B(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_159), .A2(n_177), .B1(n_197), .B2(n_199), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_159), .A2(n_177), .B1(n_250), .B2(n_251), .Y(n_249) );
INVx4_ASAP7_75t_L g549 ( .A(n_159), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g273 ( .A(n_160), .B(n_248), .C(n_249), .Y(n_273) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_161), .A2(n_171), .B(n_174), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_161), .A2(n_181), .B(n_188), .Y(n_180) );
OAI21xp5_ASAP7_75t_L g204 ( .A1(n_161), .A2(n_205), .B(n_209), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_161), .A2(n_215), .B(n_220), .Y(n_214) );
AND2x4_ASAP7_75t_L g470 ( .A(n_161), .B(n_471), .Y(n_470) );
INVx4_ASAP7_75t_SL g484 ( .A(n_161), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_161), .B(n_471), .Y(n_558) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_164), .A2(n_204), .B(n_212), .Y(n_203) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_164), .A2(n_214), .B(n_223), .Y(n_213) );
INVx2_ASAP7_75t_L g238 ( .A(n_164), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_164), .A2(n_469), .B(n_472), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_164), .A2(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g530 ( .A(n_164), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_165), .B(n_312), .Y(n_368) );
INVx2_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
OAI311xp33_ASAP7_75t_L g310 ( .A1(n_166), .A2(n_311), .A3(n_312), .B1(n_313), .C1(n_328), .Y(n_310) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_179), .Y(n_166) );
AND2x2_ASAP7_75t_L g271 ( .A(n_167), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g278 ( .A(n_167), .Y(n_278) );
AND2x2_ASAP7_75t_L g399 ( .A(n_167), .B(n_228), .Y(n_399) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_168), .B(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g255 ( .A(n_168), .B(n_179), .Y(n_255) );
AND2x2_ASAP7_75t_L g307 ( .A(n_168), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g321 ( .A(n_168), .B(n_254), .Y(n_321) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_178), .Y(n_168) );
INVx4_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_169), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_169), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .Y(n_174) );
INVx2_ASAP7_75t_L g228 ( .A(n_179), .Y(n_228) );
AND2x2_ASAP7_75t_L g270 ( .A(n_179), .B(n_254), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .C(n_185), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_183), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_183), .A2(n_561), .B(n_562), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_185), .A2(n_536), .B(n_537), .C(n_538), .Y(n_535) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_186), .A2(n_210), .B(n_211), .Y(n_209) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g480 ( .A(n_187), .Y(n_480) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_200), .Y(n_192) );
OR2x2_ASAP7_75t_L g365 ( .A(n_193), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_193), .B(n_371), .Y(n_382) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_194), .B(n_378), .Y(n_377) );
BUFx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g239 ( .A(n_195), .Y(n_239) );
AND2x2_ASAP7_75t_L g306 ( .A(n_195), .B(n_233), .Y(n_306) );
AND2x2_ASAP7_75t_L g317 ( .A(n_195), .B(n_213), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_195), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_200), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_200), .B(n_267), .Y(n_311) );
INVx2_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g298 ( .A(n_201), .B(n_257), .Y(n_298) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_213), .Y(n_201) );
INVx2_ASAP7_75t_L g231 ( .A(n_202), .Y(n_231) );
AND2x2_ASAP7_75t_L g325 ( .A(n_202), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g243 ( .A(n_203), .Y(n_243) );
OR2x2_ASAP7_75t_L g342 ( .A(n_203), .B(n_343), .Y(n_342) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_203), .Y(n_405) );
AND2x2_ASAP7_75t_L g244 ( .A(n_213), .B(n_239), .Y(n_244) );
INVx1_ASAP7_75t_L g265 ( .A(n_213), .Y(n_265) );
AND2x2_ASAP7_75t_L g286 ( .A(n_213), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g327 ( .A(n_213), .Y(n_327) );
INVx1_ASAP7_75t_L g343 ( .A(n_213), .Y(n_343) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_213), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVxp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_226), .B(n_331), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_226), .A2(n_316), .B1(n_365), .B2(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
OAI211xp5_ASAP7_75t_SL g408 ( .A1(n_227), .A2(n_409), .B(n_411), .C(n_429), .Y(n_408) );
INVx2_ASAP7_75t_L g261 ( .A(n_228), .Y(n_261) );
AND2x2_ASAP7_75t_L g319 ( .A(n_228), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g330 ( .A(n_228), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_229), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
AND2x2_ASAP7_75t_L g303 ( .A(n_230), .B(n_267), .Y(n_303) );
BUFx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g335 ( .A(n_231), .B(n_326), .Y(n_335) );
AND2x2_ASAP7_75t_L g354 ( .A(n_231), .B(n_268), .Y(n_354) );
AND2x4_ASAP7_75t_L g290 ( .A(n_232), .B(n_264), .Y(n_290) );
AND2x2_ASAP7_75t_L g428 ( .A(n_232), .B(n_404), .Y(n_428) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_239), .Y(n_232) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_233), .Y(n_257) );
INVx1_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
INVx1_ASAP7_75t_L g367 ( .A(n_233), .Y(n_367) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_236), .Y(n_482) );
INVx2_ASAP7_75t_L g550 ( .A(n_236), .Y(n_550) );
INVx1_ASAP7_75t_L g527 ( .A(n_238), .Y(n_527) );
OR2x2_ASAP7_75t_L g258 ( .A(n_239), .B(n_243), .Y(n_258) );
AND2x2_ASAP7_75t_L g267 ( .A(n_239), .B(n_268), .Y(n_267) );
NOR2xp67_ASAP7_75t_L g287 ( .A(n_239), .B(n_288), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_245), .B1(n_256), .B2(n_259), .C(n_263), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_242), .A2(n_264), .B(n_266), .C(n_269), .Y(n_263) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g288 ( .A(n_243), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_243), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_243), .B(n_265), .Y(n_371) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_243), .Y(n_378) );
AND2x2_ASAP7_75t_L g296 ( .A(n_244), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g333 ( .A(n_244), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_255), .Y(n_245) );
INVx2_ASAP7_75t_L g324 ( .A(n_246), .Y(n_324) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_246), .A2(n_257), .B1(n_374), .B2(n_376), .C1(n_377), .C2(n_379), .Y(n_373) );
AND2x2_ASAP7_75t_L g430 ( .A(n_246), .B(n_399), .Y(n_430) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_254), .Y(n_246) );
INVx1_ASAP7_75t_L g320 ( .A(n_247), .Y(n_320) );
AO21x1_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_252), .Y(n_247) );
INVx3_ASAP7_75t_L g497 ( .A(n_248), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_248), .B(n_517), .Y(n_516) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_248), .A2(n_533), .B(n_540), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_248), .B(n_541), .Y(n_540) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_248), .A2(n_556), .B(n_563), .Y(n_555) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g272 ( .A(n_253), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g358 ( .A(n_255), .B(n_292), .Y(n_358) );
AOI21xp33_ASAP7_75t_L g369 ( .A1(n_256), .A2(n_370), .B(n_372), .Y(n_369) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g297 ( .A(n_257), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_257), .B(n_264), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_257), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx3_ASAP7_75t_L g323 ( .A(n_261), .Y(n_323) );
OR2x2_ASAP7_75t_L g375 ( .A(n_261), .B(n_297), .Y(n_375) );
AND2x2_ASAP7_75t_L g291 ( .A(n_262), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g329 ( .A(n_262), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_262), .B(n_323), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_262), .B(n_319), .Y(n_345) );
AND2x2_ASAP7_75t_L g349 ( .A(n_262), .B(n_331), .Y(n_349) );
INVxp67_ASAP7_75t_L g281 ( .A(n_264), .Y(n_281) );
BUFx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_266), .A2(n_339), .B1(n_344), .B2(n_345), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_266), .B(n_371), .Y(n_401) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g387 ( .A(n_267), .B(n_378), .Y(n_387) );
AND2x2_ASAP7_75t_L g416 ( .A(n_267), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g421 ( .A(n_267), .B(n_371), .Y(n_421) );
INVx1_ASAP7_75t_L g334 ( .A(n_268), .Y(n_334) );
BUFx2_ASAP7_75t_L g340 ( .A(n_268), .Y(n_340) );
INVx1_ASAP7_75t_L g425 ( .A(n_269), .Y(n_425) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_270), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g301 ( .A(n_271), .Y(n_301) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_272), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g284 ( .A(n_272), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g293 ( .A(n_272), .Y(n_293) );
INVx3_ASAP7_75t_L g331 ( .A(n_272), .Y(n_331) );
OR2x2_ASAP7_75t_L g397 ( .A(n_272), .B(n_398), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B(n_282), .C(n_294), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_275), .A2(n_412), .B1(n_419), .B2(n_421), .C(n_422), .Y(n_411) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_283), .B(n_289), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_285), .B(n_323), .Y(n_337) );
AND2x2_ASAP7_75t_L g379 ( .A(n_285), .B(n_319), .Y(n_379) );
INVx1_ASAP7_75t_SL g392 ( .A(n_286), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_286), .B(n_340), .Y(n_395) );
INVx1_ASAP7_75t_L g413 ( .A(n_287), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_291), .A2(n_381), .B1(n_383), .B2(n_387), .C(n_388), .Y(n_380) );
AND2x2_ASAP7_75t_L g407 ( .A(n_292), .B(n_399), .Y(n_407) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g391 ( .A(n_293), .Y(n_391) );
AOI21xp33_ASAP7_75t_SL g294 ( .A1(n_295), .A2(n_298), .B(n_299), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g362 ( .A(n_297), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
INVx1_ASAP7_75t_L g376 ( .A(n_299), .Y(n_376) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_307), .C(n_310), .Y(n_302) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_303), .A2(n_341), .A3(n_428), .B(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g403 ( .A(n_306), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g424 ( .A(n_306), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_308), .B(n_323), .Y(n_351) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g426 ( .A(n_309), .B(n_323), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B1(n_322), .B2(n_325), .Y(n_313) );
NAND2xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_317), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g353 ( .A(n_317), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g356 ( .A(n_317), .B(n_340), .Y(n_356) );
AND2x2_ASAP7_75t_L g410 ( .A(n_317), .B(n_405), .Y(n_410) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g385 ( .A(n_321), .Y(n_385) );
NOR2xp67_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OAI32xp33_ASAP7_75t_L g388 ( .A1(n_323), .A2(n_357), .A3(n_389), .B1(n_391), .B2(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g363 ( .A(n_326), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_326), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g386 ( .A(n_330), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_336), .C(n_338), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_334), .B(n_371), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_335), .A2(n_347), .B1(n_348), .B2(n_349), .C(n_350), .Y(n_346) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g347 ( .A(n_345), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B1(n_355), .B2(n_357), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND4xp25_ASAP7_75t_SL g412 ( .A(n_355), .B(n_413), .C(n_414), .D(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NAND4xp25_ASAP7_75t_SL g359 ( .A(n_360), .B(n_373), .C(n_380), .D(n_393), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B(n_368), .C(n_369), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g390 ( .A(n_366), .Y(n_390) );
INVx2_ASAP7_75t_L g414 ( .A(n_371), .Y(n_414) );
OR2x2_ASAP7_75t_L g423 ( .A(n_378), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_400), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g419 ( .A(n_399), .B(n_420), .Y(n_419) );
AOI21xp33_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_402), .B(n_406), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g437 ( .A(n_433), .Y(n_437) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g441 ( .A(n_434), .Y(n_441) );
NAND4xp25_ASAP7_75t_SL g442 ( .A(n_438), .B(n_443), .C(n_444), .D(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_454), .B2(n_761), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B1(n_460), .B2(n_463), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g762 ( .A(n_456), .Y(n_762) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g763 ( .A(n_458), .Y(n_763) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g764 ( .A(n_461), .Y(n_764) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx4_ASAP7_75t_L g765 ( .A(n_463), .Y(n_765) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR5x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_634), .C(n_712), .D(n_736), .E(n_753), .Y(n_464) );
OAI211xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_506), .B(n_552), .C(n_611), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_486), .Y(n_466) );
AND2x2_ASAP7_75t_L g565 ( .A(n_467), .B(n_488), .Y(n_565) );
INVx5_ASAP7_75t_SL g593 ( .A(n_467), .Y(n_593) );
AND2x2_ASAP7_75t_L g629 ( .A(n_467), .B(n_614), .Y(n_629) );
OR2x2_ASAP7_75t_L g668 ( .A(n_467), .B(n_487), .Y(n_668) );
OR2x2_ASAP7_75t_L g699 ( .A(n_467), .B(n_590), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_467), .B(n_603), .Y(n_735) );
AND2x2_ASAP7_75t_L g747 ( .A(n_467), .B(n_590), .Y(n_747) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_485), .Y(n_467) );
BUFx2_ASAP7_75t_L g522 ( .A(n_470), .Y(n_522) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_474), .A2(n_484), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g544 ( .A1(n_474), .A2(n_484), .B(n_545), .C(n_546), .Y(n_544) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_481), .C(n_482), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_479), .A2(n_482), .B(n_514), .C(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g746 ( .A(n_486), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g609 ( .A(n_487), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_498), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_488), .B(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_488), .Y(n_602) );
INVx3_ASAP7_75t_L g617 ( .A(n_488), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_488), .B(n_498), .Y(n_641) );
OR2x2_ASAP7_75t_L g650 ( .A(n_488), .B(n_593), .Y(n_650) );
AND2x2_ASAP7_75t_L g654 ( .A(n_488), .B(n_614), .Y(n_654) );
AND2x2_ASAP7_75t_L g660 ( .A(n_488), .B(n_661), .Y(n_660) );
INVxp67_ASAP7_75t_L g697 ( .A(n_488), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_488), .B(n_555), .Y(n_711) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_496), .Y(n_488) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_497), .A2(n_543), .B(n_551), .Y(n_542) );
OR2x2_ASAP7_75t_L g603 ( .A(n_498), .B(n_555), .Y(n_603) );
AND2x2_ASAP7_75t_L g614 ( .A(n_498), .B(n_590), .Y(n_614) );
AND2x2_ASAP7_75t_L g626 ( .A(n_498), .B(n_617), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_498), .B(n_555), .Y(n_649) );
INVx1_ASAP7_75t_SL g661 ( .A(n_498), .Y(n_661) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g554 ( .A(n_499), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_499), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
AND2x2_ASAP7_75t_L g574 ( .A(n_508), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_508), .B(n_531), .Y(n_578) );
AND2x2_ASAP7_75t_L g581 ( .A(n_508), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_508), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g606 ( .A(n_508), .B(n_597), .Y(n_606) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_508), .Y(n_625) );
AND2x2_ASAP7_75t_L g646 ( .A(n_508), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g656 ( .A(n_508), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g702 ( .A(n_508), .B(n_585), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_508), .B(n_608), .Y(n_729) );
INVx5_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g599 ( .A(n_509), .Y(n_599) );
AND2x2_ASAP7_75t_L g665 ( .A(n_509), .B(n_597), .Y(n_665) );
AND2x2_ASAP7_75t_L g749 ( .A(n_509), .B(n_617), .Y(n_749) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_518), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g738 ( .A(n_518), .Y(n_738) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_531), .Y(n_518) );
AND2x2_ASAP7_75t_L g568 ( .A(n_519), .B(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_L g577 ( .A(n_519), .B(n_575), .Y(n_577) );
INVx5_ASAP7_75t_L g585 ( .A(n_519), .Y(n_585) );
AND2x2_ASAP7_75t_L g608 ( .A(n_519), .B(n_542), .Y(n_608) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_519), .Y(n_645) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_528), .Y(n_519) );
AOI21xp5_ASAP7_75t_SL g520 ( .A1(n_521), .A2(n_523), .B(n_527), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g686 ( .A(n_531), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_531), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g719 ( .A(n_531), .B(n_585), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g748 ( .A1(n_531), .A2(n_642), .B(n_749), .C(n_750), .Y(n_748) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_542), .Y(n_531) );
BUFx2_ASAP7_75t_L g569 ( .A(n_532), .Y(n_569) );
INVx2_ASAP7_75t_L g573 ( .A(n_532), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_539), .Y(n_533) );
INVx2_ASAP7_75t_L g575 ( .A(n_542), .Y(n_575) );
AND2x2_ASAP7_75t_L g582 ( .A(n_542), .B(n_573), .Y(n_582) );
AND2x2_ASAP7_75t_L g673 ( .A(n_542), .B(n_585), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AOI211x1_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_566), .B(n_579), .C(n_604), .Y(n_552) );
INVx1_ASAP7_75t_L g670 ( .A(n_553), .Y(n_670) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_565), .Y(n_553) );
INVx5_ASAP7_75t_SL g590 ( .A(n_555), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_555), .B(n_660), .Y(n_659) );
AOI311xp33_ASAP7_75t_L g678 ( .A1(n_555), .A2(n_679), .A3(n_681), .B(n_682), .C(n_688), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_555), .A2(n_626), .B(n_714), .C(n_717), .Y(n_713) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_559), .Y(n_556) );
INVxp67_ASAP7_75t_L g633 ( .A(n_565), .Y(n_633) );
NAND4xp25_ASAP7_75t_SL g566 ( .A(n_567), .B(n_570), .C(n_576), .D(n_578), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_567), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g624 ( .A(n_568), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_571), .B(n_577), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_571), .B(n_584), .Y(n_704) );
BUFx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_572), .B(n_585), .Y(n_722) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g597 ( .A(n_573), .Y(n_597) );
INVxp67_ASAP7_75t_L g632 ( .A(n_574), .Y(n_632) );
AND2x4_ASAP7_75t_L g584 ( .A(n_575), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g658 ( .A(n_575), .B(n_597), .Y(n_658) );
INVx1_ASAP7_75t_L g685 ( .A(n_575), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_575), .B(n_672), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_576), .B(n_646), .Y(n_666) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_577), .B(n_599), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_577), .B(n_646), .Y(n_745) );
INVx1_ASAP7_75t_L g756 ( .A(n_578), .Y(n_756) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_583), .B(n_586), .C(n_594), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g598 ( .A(n_582), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g636 ( .A(n_582), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g618 ( .A(n_583), .Y(n_618) );
AND2x2_ASAP7_75t_L g595 ( .A(n_584), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_584), .B(n_646), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_584), .B(n_665), .Y(n_689) );
OR2x2_ASAP7_75t_L g605 ( .A(n_585), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g637 ( .A(n_585), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_585), .B(n_597), .Y(n_652) );
AND2x2_ASAP7_75t_L g709 ( .A(n_585), .B(n_665), .Y(n_709) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_585), .Y(n_716) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_587), .A2(n_599), .B1(n_721), .B2(n_723), .C(n_726), .Y(n_720) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g610 ( .A(n_590), .B(n_593), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_590), .B(n_660), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_590), .B(n_617), .Y(n_725) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g710 ( .A(n_592), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g724 ( .A(n_592), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_593), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g621 ( .A(n_593), .B(n_614), .Y(n_621) );
AND2x2_ASAP7_75t_L g691 ( .A(n_593), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_593), .B(n_640), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_593), .B(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_598), .B(n_600), .Y(n_594) );
INVx2_ASAP7_75t_L g627 ( .A(n_595), .Y(n_627) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g647 ( .A(n_597), .Y(n_647) );
OR2x2_ASAP7_75t_L g651 ( .A(n_599), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g754 ( .A(n_599), .B(n_722), .Y(n_754) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .B(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g758 ( .A(n_605), .Y(n_758) );
INVx2_ASAP7_75t_SL g672 ( .A(n_606), .Y(n_672) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_609), .A2(n_690), .B(n_754), .C(n_755), .Y(n_753) );
OAI322xp33_ASAP7_75t_SL g622 ( .A1(n_610), .A2(n_623), .A3(n_626), .B1(n_627), .B2(n_628), .C1(n_630), .C2(n_633), .Y(n_622) );
INVx2_ASAP7_75t_L g642 ( .A(n_610), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_618), .B1(n_619), .B2(n_621), .C(n_622), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI22xp33_ASAP7_75t_SL g688 ( .A1(n_613), .A2(n_689), .B1(n_690), .B2(n_693), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_614), .B(n_617), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_614), .B(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g687 ( .A(n_616), .B(n_649), .Y(n_687) );
INVx1_ASAP7_75t_L g677 ( .A(n_617), .Y(n_677) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_621), .A2(n_731), .B(n_733), .Y(n_730) );
AOI21xp33_ASAP7_75t_L g655 ( .A1(n_623), .A2(n_656), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp67_ASAP7_75t_SL g684 ( .A(n_625), .B(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_625), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g741 ( .A(n_626), .Y(n_741) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_635), .B(n_662), .C(n_678), .D(n_694), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_643), .C(n_655), .Y(n_635) );
INVx1_ASAP7_75t_L g727 ( .A(n_636), .Y(n_727) );
AND2x2_ASAP7_75t_L g675 ( .A(n_637), .B(n_658), .Y(n_675) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_642), .B(n_677), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B1(n_651), .B2(n_653), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_645), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g693 ( .A(n_646), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_646), .A2(n_685), .B(n_708), .C(n_710), .Y(n_707) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g692 ( .A(n_649), .Y(n_692) );
INVx1_ASAP7_75t_L g752 ( .A(n_650), .Y(n_752) );
NAND2xp33_ASAP7_75t_SL g742 ( .A(n_651), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g681 ( .A(n_660), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_666), .B(n_667), .C(n_669), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_674), .B2(n_676), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_672), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_677), .B(n_698), .Y(n_760) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI21xp33_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_686), .B(n_687), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_700), .B1(n_703), .B2(n_705), .C(n_707), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_710), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
NAND3xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_720), .C(n_730), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI211xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B(n_739), .C(n_748), .Y(n_736) );
INVx1_ASAP7_75t_L g757 ( .A(n_737), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_742), .B1(n_744), .B2(n_746), .Y(n_739) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_755) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI22x1_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_761) );
endmodule