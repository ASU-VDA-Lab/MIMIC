module fake_jpeg_69_n_179 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_46),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_44),
.B(n_45),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_56),
.B1(n_51),
.B2(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_79),
.B1(n_48),
.B2(n_67),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_44),
.B1(n_55),
.B2(n_50),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_46),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_49),
.B1(n_43),
.B2(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_79),
.B(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_89),
.Y(n_101)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_88),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_78),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_3),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_59),
.B(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_112),
.Y(n_121)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_94),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_110),
.B1(n_111),
.B2(n_5),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_10),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_59),
.B1(n_15),
.B2(n_17),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_4),
.Y(n_114)
);

XNOR2x1_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_4),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_123),
.Y(n_142)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_5),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_35),
.B1(n_20),
.B2(n_21),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_7),
.B(n_8),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_129),
.B(n_11),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_19),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_131),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_7),
.B(n_9),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_9),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_10),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_31),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_145),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_150),
.B1(n_24),
.B2(n_27),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_12),
.B1(n_22),
.B2(n_23),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_153),
.B(n_155),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_128),
.C(n_125),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_151),
.C(n_161),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_160),
.B1(n_161),
.B2(n_150),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_146),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_137),
.B(n_138),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_28),
.B1(n_30),
.B2(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_164),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_155),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_136),
.C(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_142),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_171),
.B(n_169),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_165),
.C(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_165),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_148),
.Y(n_179)
);


endmodule