module fake_jpeg_3323_n_40 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.C(n_20),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_19),
.B(n_16),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_16),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_14),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_SL g25 ( 
.A1(n_24),
.A2(n_20),
.B(n_17),
.C(n_18),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_14),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_27),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_17),
.C(n_15),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.C(n_31),
.Y(n_33)
);

MAJx2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_25),
.C(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_7),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_36),
.B(n_33),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_37),
.B1(n_9),
.B2(n_10),
.Y(n_40)
);


endmodule