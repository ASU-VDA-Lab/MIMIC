module fake_ibex_1694_n_5272 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_5272);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_5272;

wire n_4557;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_962;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_4569;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_2253;
wire n_4479;
wire n_3858;
wire n_4173;
wire n_5261;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_5033;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_971;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_4757;
wire n_5254;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_5252;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_5099;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_5163;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_1471;
wire n_3441;
wire n_4559;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_5157;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_2422;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_972;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_977;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2420;
wire n_2380;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1072;
wire n_2194;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_3096;
wire n_2059;
wire n_1278;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_4082;
wire n_4367;
wire n_3273;
wire n_4282;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_985;
wire n_4611;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_4895;
wire n_3354;
wire n_4069;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_2574;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_1518;
wire n_4350;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_4686;
wire n_4682;
wire n_2914;
wire n_1833;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_4733;
wire n_987;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_1012;
wire n_960;
wire n_4412;
wire n_4266;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_3857;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_2969;
wire n_3550;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_2978;
wire n_3502;
wire n_3935;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_4926;
wire n_5043;
wire n_4688;
wire n_5097;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_969;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_3484;
wire n_2485;
wire n_4477;
wire n_5177;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_3726;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4545;
wire n_2643;
wire n_4246;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5221;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4997;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_3633;
wire n_1731;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_2076;
wire n_974;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_959;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_5089;
wire n_2573;
wire n_1793;
wire n_2424;
wire n_2390;
wire n_965;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_4991;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_3703;
wire n_5116;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_954;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_998;
wire n_1729;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_3398;
wire n_3718;
wire n_4878;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_5193;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_5153;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_4636;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_1067;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4699;
wire n_4228;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_1660;
wire n_4000;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_5159;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_5096;
wire n_3712;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_5217;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_976;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_3327;
wire n_1114;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_1175;
wire n_4408;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_5167;
wire n_4565;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_956;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5076;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_5013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_2671;
wire n_3296;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_953;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_3036;
wire n_5012;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_5208;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_955;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_1640;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_5245;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_1743;
wire n_5061;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_5184;
wire n_4943;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_4159;
wire n_4372;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_4897;
wire n_963;
wire n_2139;
wire n_3693;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_5204;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_3722;
wire n_3802;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_4806;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_2564;
wire n_5110;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_2114;
wire n_1609;
wire n_3530;
wire n_1132;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_4999;
wire n_2660;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_4604;
wire n_5123;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_3282;
wire n_5144;
wire n_1003;
wire n_2708;
wire n_5164;
wire n_2748;
wire n_2224;
wire n_2233;
wire n_2499;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5147;
wire n_1553;
wire n_3542;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4681;
wire n_4253;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_2481;
wire n_4409;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_5050;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_4500;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_2414;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_3328;
wire n_2763;
wire n_994;
wire n_5136;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_961;
wire n_3735;
wire n_2127;
wire n_3028;
wire n_3228;
wire n_5079;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_1839;
wire n_5160;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2108;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_4373;
wire n_3462;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_5101;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_2894;
wire n_5249;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_975;
wire n_4900;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_2315;
wire n_3623;
wire n_2157;
wire n_3446;
wire n_5223;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_5106;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_1105;
wire n_5198;
wire n_2898;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_4982;
wire n_1769;
wire n_1060;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_4053;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_1693;
wire n_2081;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_3989;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_967;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_3430;
wire n_1685;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_5038;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_5248;
wire n_4088;
wire n_2136;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4972;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_983;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_4967;
wire n_1080;
wire n_2290;
wire n_957;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4668;
wire n_2383;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_3033;
wire n_2151;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_5211;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_1606;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_979;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_4981;
wire n_978;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_2719;
wire n_2213;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_2646;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_4156;
wire n_3754;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_1452;
wire n_4953;
wire n_4570;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_1985;
wire n_1140;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_4407;
wire n_5077;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_3680;
wire n_3624;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1566;
wire n_1464;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_1009;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2991;
wire n_2699;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_4427;
wire n_3505;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_2525;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_5105;
wire n_964;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_5187;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_3588;
wire n_5220;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1458;
wire n_1694;
wire n_2271;
wire n_2356;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_2642;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_5091;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_4860;
wire n_4438;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_993;
wire n_2581;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_958;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5118;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_5112;
wire n_3042;
wire n_2561;
wire n_2491;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_3551;
wire n_4147;
wire n_3992;
wire n_4811;
wire n_5093;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_1419;
wire n_4738;
wire n_980;
wire n_1193;
wire n_3557;
wire n_2928;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_4086;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_966;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_1791;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_1164;
wire n_3749;
wire n_4452;
wire n_3691;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_4978;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_736),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_717),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_650),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_726),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_67),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_15),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_491),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_358),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_912),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_433),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_582),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_716),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_64),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_294),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_940),
.Y(n_967)
);

BUFx10_ASAP7_75t_L g968 ( 
.A(n_586),
.Y(n_968)
);

CKINVDCx16_ASAP7_75t_R g969 ( 
.A(n_877),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_64),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_153),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_950),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_488),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_243),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_612),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_878),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_435),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_63),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_17),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_67),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_765),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_850),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_300),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_363),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_65),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_158),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_327),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_820),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_167),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_362),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_844),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_770),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_187),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_111),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_720),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_474),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_44),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_184),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_74),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_866),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_943),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_600),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_97),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_829),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_926),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_597),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_868),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_835),
.Y(n_1008)
);

BUFx5_ASAP7_75t_L g1009 ( 
.A(n_232),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_294),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_534),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_586),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_144),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_551),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_431),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_298),
.Y(n_1016)
);

BUFx10_ASAP7_75t_L g1017 ( 
.A(n_602),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_554),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_921),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_911),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_198),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_150),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_628),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_816),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_783),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_440),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_714),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_856),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_900),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_528),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_823),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_683),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_916),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_874),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_864),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_858),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_194),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_820),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_818),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_217),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_502),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_650),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_592),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_550),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_48),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_171),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_110),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_347),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_201),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_22),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_823),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_290),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_731),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_838),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_61),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_88),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_927),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_172),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_589),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_561),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_229),
.Y(n_1061)
);

CKINVDCx16_ASAP7_75t_R g1062 ( 
.A(n_139),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_892),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_264),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_742),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_123),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_121),
.Y(n_1067)
);

CKINVDCx16_ASAP7_75t_R g1068 ( 
.A(n_824),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_241),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_770),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_321),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_182),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_836),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_492),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_62),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_773),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_486),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_923),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_565),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_374),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_931),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_466),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_96),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_577),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_205),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_36),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_932),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_318),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_798),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_671),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_407),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_273),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_919),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_112),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_761),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_937),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_209),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_378),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_733),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_573),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_213),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_479),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_913),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_493),
.Y(n_1104)
);

CKINVDCx16_ASAP7_75t_R g1105 ( 
.A(n_145),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_38),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_562),
.Y(n_1107)
);

BUFx10_ASAP7_75t_L g1108 ( 
.A(n_336),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_138),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_861),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_860),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_675),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_382),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_950),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_712),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_532),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_596),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_581),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_705),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_459),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_11),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_939),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_507),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_598),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_685),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_244),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_834),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_288),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_656),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_904),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_937),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_837),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_85),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_151),
.Y(n_1134)
);

CKINVDCx16_ASAP7_75t_R g1135 ( 
.A(n_656),
.Y(n_1135)
);

INVxp33_ASAP7_75t_R g1136 ( 
.A(n_723),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_500),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_154),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_318),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_332),
.Y(n_1140)
);

CKINVDCx16_ASAP7_75t_R g1141 ( 
.A(n_161),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_582),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_220),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_21),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_928),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_940),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_939),
.Y(n_1147)
);

BUFx10_ASAP7_75t_L g1148 ( 
.A(n_902),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_485),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_77),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_133),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_122),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_641),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_639),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_453),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_22),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_404),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_530),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_90),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_227),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_573),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_349),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_867),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_480),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_273),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_359),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_410),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_803),
.Y(n_1168)
);

BUFx10_ASAP7_75t_L g1169 ( 
.A(n_773),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_665),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_639),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_243),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_855),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_829),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_907),
.Y(n_1175)
);

CKINVDCx14_ASAP7_75t_R g1176 ( 
.A(n_922),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_338),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_925),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_616),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_341),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_21),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_290),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_807),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_236),
.Y(n_1184)
);

CKINVDCx16_ASAP7_75t_R g1185 ( 
.A(n_892),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_889),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_780),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_373),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_382),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_47),
.Y(n_1190)
);

CKINVDCx16_ASAP7_75t_R g1191 ( 
.A(n_851),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_605),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_326),
.Y(n_1193)
);

BUFx5_ASAP7_75t_L g1194 ( 
.A(n_558),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_699),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_508),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_131),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_905),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_150),
.Y(n_1199)
);

BUFx10_ASAP7_75t_L g1200 ( 
.A(n_350),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_629),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_209),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_411),
.Y(n_1203)
);

CKINVDCx14_ASAP7_75t_R g1204 ( 
.A(n_952),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_293),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_583),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_637),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_831),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_450),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_564),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_321),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_161),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_25),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_819),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_886),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_593),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_443),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_522),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_457),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_886),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_765),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_156),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_100),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_934),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_490),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_871),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_822),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_599),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_258),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_20),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_839),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_95),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_779),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_603),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_53),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_869),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_403),
.Y(n_1237)
);

BUFx10_ASAP7_75t_L g1238 ( 
.A(n_743),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_808),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_421),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_840),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_934),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_859),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_289),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_790),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_936),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_325),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_67),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_397),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_552),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_675),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_862),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_360),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_797),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_802),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_777),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_872),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_903),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_898),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_683),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_514),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_885),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_340),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_581),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_693),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_882),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_48),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_917),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_588),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_435),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_903),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_925),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_618),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_924),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_427),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_901),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_854),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_666),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_385),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_865),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_131),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_84),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_640),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_468),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_711),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_557),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_762),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_814),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_492),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_782),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_810),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_941),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_651),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_50),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_592),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_749),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_335),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_776),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_929),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_908),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_734),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_400),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_462),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_343),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_93),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_904),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_841),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_162),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_493),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_897),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_909),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_174),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_355),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_603),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_481),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_689),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_784),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_930),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_705),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_665),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_484),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_736),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_37),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_659),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_184),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_848),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_888),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_230),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_532),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_821),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_845),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_377),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_245),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_337),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_463),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_202),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_740),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_475),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_407),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_469),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_168),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_743),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_640),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_848),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_37),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_641),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_512),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_841),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_625),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_111),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_511),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_884),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_817),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_214),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_888),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_15),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_420),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_558),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_935),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_238),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_637),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_363),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_164),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_269),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_357),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_893),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_808),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_828),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_475),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_405),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_314),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_529),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_229),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_826),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_4),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_851),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_895),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_825),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_642),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_933),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_270),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_314),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_870),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_847),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_315),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_842),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_443),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_781),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_467),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_788),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_671),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_130),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_648),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_830),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_862),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_405),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_859),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_915),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_112),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_843),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_486),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_285),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_301),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_114),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_282),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_883),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_896),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_406),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_568),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_677),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_14),
.Y(n_1412)
);

BUFx5_ASAP7_75t_L g1413 ( 
.A(n_411),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_853),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_16),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_494),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_703),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_894),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_824),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_628),
.Y(n_1420)
);

BUFx10_ASAP7_75t_L g1421 ( 
.A(n_910),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_846),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_359),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_797),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_449),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_342),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_566),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_938),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_306),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_837),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_296),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_375),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_440),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_769),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_906),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_809),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_37),
.Y(n_1437)
);

CKINVDCx16_ASAP7_75t_R g1438 ( 
.A(n_803),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_419),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_194),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_0),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_657),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_944),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_672),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_863),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_796),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_914),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_800),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_147),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_42),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_833),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_293),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_701),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_857),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_374),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_793),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_594),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_887),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_251),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_918),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_670),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_880),
.Y(n_1462)
);

BUFx5_ASAP7_75t_L g1463 ( 
.A(n_323),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_211),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_376),
.Y(n_1465)
);

CKINVDCx16_ASAP7_75t_R g1466 ( 
.A(n_593),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_354),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_569),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_105),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_825),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_517),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_508),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_430),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_16),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_894),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_491),
.Y(n_1476)
);

BUFx2_ASAP7_75t_SL g1477 ( 
.A(n_383),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_680),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_830),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_160),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_298),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_721),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_853),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_881),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_367),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_601),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_324),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_875),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_244),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_766),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_82),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_701),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_322),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_376),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_885),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_703),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_605),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_169),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_114),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_41),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_920),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_663),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_686),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_272),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_876),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_16),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_890),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_879),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_952),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_764),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_906),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_873),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_7),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_827),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_262),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_835),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_73),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_306),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_157),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_622),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_386),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_509),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_251),
.Y(n_1523)
);

BUFx10_ASAP7_75t_L g1524 ( 
.A(n_790),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_536),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_5),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_899),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_400),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_852),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_796),
.Y(n_1530)
);

CKINVDCx14_ASAP7_75t_R g1531 ( 
.A(n_891),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_849),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_529),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_945),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_587),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_23),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_854),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_693),
.Y(n_1538)
);

BUFx10_ASAP7_75t_L g1539 ( 
.A(n_553),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_289),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_355),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_522),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_162),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_712),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_723),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_372),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_296),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_832),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_760),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_122),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_942),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_938),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_769),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_0),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_978),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1009),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1441),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1176),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1156),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1513),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_964),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1176),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_964),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1531),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1009),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1088),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1531),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1088),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1156),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1142),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1142),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_970),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_980),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_999),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_958),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1204),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1204),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1045),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1106),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_957),
.Y(n_1580)
);

INVxp67_ASAP7_75t_SL g1581 ( 
.A(n_1230),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1009),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_965),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1086),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_993),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1133),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1009),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1181),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1235),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1009),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1323),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1400),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1405),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1412),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1415),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_979),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1469),
.Y(n_1597)
);

INVxp33_ASAP7_75t_SL g1598 ( 
.A(n_985),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1517),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1536),
.Y(n_1600)
);

INVxp33_ASAP7_75t_SL g1601 ( 
.A(n_994),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1230),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1009),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1500),
.Y(n_1604)
);

INVxp67_ASAP7_75t_SL g1605 ( 
.A(n_1500),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_971),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1056),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1437),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_997),
.Y(n_1609)
);

INVxp33_ASAP7_75t_L g1610 ( 
.A(n_973),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1194),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1491),
.Y(n_1612)
);

CKINVDCx20_ASAP7_75t_R g1613 ( 
.A(n_1094),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_993),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1003),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1065),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1065),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1073),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1047),
.Y(n_1619)
);

INVxp33_ASAP7_75t_SL g1620 ( 
.A(n_1050),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1073),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1055),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1219),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_998),
.B(n_0),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1219),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1225),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1075),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1225),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1313),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1313),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1427),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1083),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1427),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_1223),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1518),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1351),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1518),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1121),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1194),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1194),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1144),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1194),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1194),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1007),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1194),
.Y(n_1645)
);

CKINVDCx16_ASAP7_75t_R g1646 ( 
.A(n_969),
.Y(n_1646)
);

BUFx2_ASAP7_75t_SL g1647 ( 
.A(n_1413),
.Y(n_1647)
);

CKINVDCx14_ASAP7_75t_R g1648 ( 
.A(n_1063),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1413),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1042),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1077),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1413),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1259),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1413),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1150),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1413),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1413),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_991),
.B(n_1286),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1463),
.Y(n_1659)
);

INVxp33_ASAP7_75t_L g1660 ( 
.A(n_1385),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1474),
.Y(n_1661)
);

INVxp67_ASAP7_75t_SL g1662 ( 
.A(n_1411),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1523),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1463),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1463),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1159),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1096),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1463),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1463),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1463),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1190),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1033),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1034),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1052),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1087),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1213),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1062),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1173),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1231),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1232),
.B(n_1),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1310),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1068),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1333),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1554),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_1105),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1347),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1135),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1141),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_974),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1585),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1650),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1658),
.B(n_1165),
.Y(n_1692)
);

INVxp33_ASAP7_75t_SL g1693 ( 
.A(n_1580),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1614),
.Y(n_1694)
);

INVx5_ASAP7_75t_L g1695 ( 
.A(n_1667),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1616),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1610),
.B(n_1185),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1559),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1667),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1689),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1556),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1559),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1660),
.B(n_1191),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1558),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1565),
.Y(n_1705)
);

CKINVDCx6p67_ASAP7_75t_R g1706 ( 
.A(n_1646),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1689),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1569),
.B(n_1248),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1569),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1671),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1617),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1575),
.A2(n_955),
.B1(n_976),
.B2(n_962),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1689),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1582),
.Y(n_1714)
);

INVx4_ASAP7_75t_L g1715 ( 
.A(n_1562),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1587),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1606),
.B(n_1139),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1590),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1622),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1639),
.A2(n_1399),
.B(n_1348),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1658),
.B(n_1263),
.Y(n_1721)
);

CKINVDCx20_ASAP7_75t_R g1722 ( 
.A(n_1584),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1606),
.B(n_1189),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1663),
.B(n_1438),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1581),
.B(n_1602),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1648),
.A2(n_1282),
.B1(n_1294),
.B2(n_1267),
.Y(n_1726)
);

OAI22x1_ASAP7_75t_L g1727 ( 
.A1(n_1613),
.A2(n_1136),
.B1(n_1345),
.B2(n_1305),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1605),
.B(n_1349),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1618),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1561),
.Y(n_1730)
);

NOR2x1_ASAP7_75t_L g1731 ( 
.A(n_1555),
.B(n_1207),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1604),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1603),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1611),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1621),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1623),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1664),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1640),
.Y(n_1738)
);

BUFx12f_ASAP7_75t_L g1739 ( 
.A(n_1564),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1607),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1634),
.A2(n_1661),
.B1(n_1636),
.B2(n_1014),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1642),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1625),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1643),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1608),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1626),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1628),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1645),
.Y(n_1748)
);

CKINVDCx16_ASAP7_75t_R g1749 ( 
.A(n_1677),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1598),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1649),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1601),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1652),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1653),
.A2(n_1376),
.B1(n_1450),
.B2(n_1357),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1682),
.A2(n_1020),
.B1(n_1026),
.B2(n_1011),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1654),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1656),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1657),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1659),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1629),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1665),
.Y(n_1761)
);

OA21x2_ASAP7_75t_L g1762 ( 
.A1(n_1668),
.A2(n_1670),
.B(n_1669),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1557),
.B(n_1383),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1622),
.B(n_1499),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1612),
.B(n_1506),
.Y(n_1765)
);

AND2x6_ASAP7_75t_L g1766 ( 
.A(n_1563),
.B(n_974),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1672),
.Y(n_1767)
);

AND2x6_ASAP7_75t_L g1768 ( 
.A(n_1566),
.B(n_974),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1630),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1620),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1673),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1631),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1583),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1633),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1674),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1635),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1637),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1675),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1596),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1560),
.B(n_1414),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1609),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1572),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1678),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1573),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1574),
.Y(n_1785)
);

OA21x2_ASAP7_75t_L g1786 ( 
.A1(n_1578),
.A2(n_956),
.B(n_954),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1579),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1615),
.Y(n_1788)
);

NAND2xp33_ASAP7_75t_R g1789 ( 
.A(n_1619),
.B(n_1526),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1568),
.B(n_1466),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1679),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_L g1792 ( 
.A(n_1570),
.B(n_1422),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1681),
.Y(n_1793)
);

BUFx3_ASAP7_75t_L g1794 ( 
.A(n_1627),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1683),
.Y(n_1795)
);

OA21x2_ASAP7_75t_L g1796 ( 
.A1(n_1586),
.A2(n_967),
.B(n_961),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1632),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1567),
.B(n_1276),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1571),
.B(n_953),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1686),
.Y(n_1800)
);

BUFx8_ASAP7_75t_SL g1801 ( 
.A(n_1685),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1638),
.Y(n_1802)
);

BUFx8_ASAP7_75t_L g1803 ( 
.A(n_1687),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1588),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1589),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1591),
.Y(n_1806)
);

OA21x2_ASAP7_75t_L g1807 ( 
.A1(n_1592),
.A2(n_1594),
.B(n_1593),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1662),
.A2(n_1352),
.B1(n_1375),
.B2(n_1314),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1595),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1597),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1599),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1600),
.Y(n_1812)
);

OA21x2_ASAP7_75t_L g1813 ( 
.A1(n_1680),
.A2(n_1006),
.B(n_1005),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1647),
.Y(n_1814)
);

CKINVDCx11_ASAP7_75t_R g1815 ( 
.A(n_1688),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1641),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1655),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1680),
.Y(n_1818)
);

CKINVDCx8_ASAP7_75t_R g1819 ( 
.A(n_1666),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1624),
.Y(n_1820)
);

INVx5_ASAP7_75t_L g1821 ( 
.A(n_1644),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1576),
.B(n_959),
.Y(n_1822)
);

OA21x2_ASAP7_75t_L g1823 ( 
.A1(n_1676),
.A2(n_1012),
.B(n_1008),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1577),
.B(n_960),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1684),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1651),
.Y(n_1826)
);

OAI21x1_ASAP7_75t_L g1827 ( 
.A1(n_1639),
.A2(n_1472),
.B(n_1403),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1569),
.B(n_963),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1569),
.B(n_966),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1606),
.B(n_1433),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1610),
.B(n_968),
.Y(n_1831)
);

INVx5_ASAP7_75t_L g1832 ( 
.A(n_1667),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1598),
.B(n_972),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1606),
.B(n_1492),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1559),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1610),
.B(n_968),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1689),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1598),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1585),
.Y(n_1839)
);

OA21x2_ASAP7_75t_L g1840 ( 
.A1(n_1639),
.A2(n_1016),
.B(n_1015),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1559),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1650),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1598),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1559),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1585),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1606),
.B(n_1498),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1585),
.Y(n_1847)
);

OA21x2_ASAP7_75t_L g1848 ( 
.A1(n_1639),
.A2(n_1022),
.B(n_1018),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1689),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1559),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_1585),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1585),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1559),
.Y(n_1853)
);

BUFx8_ASAP7_75t_L g1854 ( 
.A(n_1663),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1585),
.Y(n_1855)
);

BUFx2_ASAP7_75t_L g1856 ( 
.A(n_1648),
.Y(n_1856)
);

INVx4_ASAP7_75t_L g1857 ( 
.A(n_1558),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1606),
.A2(n_1458),
.B1(n_1471),
.B2(n_1429),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1689),
.Y(n_1859)
);

NOR2x1_ASAP7_75t_L g1860 ( 
.A(n_1555),
.B(n_1520),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1648),
.A2(n_975),
.B1(n_981),
.B2(n_977),
.Y(n_1861)
);

INVx6_ASAP7_75t_L g1862 ( 
.A(n_1650),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1648),
.Y(n_1863)
);

CKINVDCx20_ASAP7_75t_R g1864 ( 
.A(n_1575),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1585),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1569),
.B(n_982),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1559),
.Y(n_1867)
);

OA21x2_ASAP7_75t_L g1868 ( 
.A1(n_1639),
.A2(n_1031),
.B(n_1029),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1606),
.B(n_1035),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1559),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1610),
.B(n_1017),
.Y(n_1871)
);

OA21x2_ASAP7_75t_L g1872 ( 
.A1(n_1639),
.A2(n_1037),
.B(n_1036),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1559),
.Y(n_1873)
);

INVx6_ASAP7_75t_L g1874 ( 
.A(n_1650),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1658),
.B(n_983),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1559),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1585),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1585),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1585),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1610),
.B(n_1017),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1559),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1585),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1622),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1606),
.B(n_1039),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1569),
.B(n_984),
.Y(n_1885)
);

AND2x6_ASAP7_75t_L g1886 ( 
.A(n_1561),
.B(n_974),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1689),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1569),
.B(n_986),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1585),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1648),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1606),
.B(n_1040),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1559),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1598),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1585),
.Y(n_1894)
);

INVx4_ASAP7_75t_L g1895 ( 
.A(n_1558),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1606),
.B(n_1041),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1559),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1559),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1689),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1598),
.B(n_987),
.Y(n_1900)
);

BUFx6f_ASAP7_75t_L g1901 ( 
.A(n_1689),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1606),
.A2(n_995),
.B1(n_996),
.B2(n_988),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1648),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1689),
.Y(n_1904)
);

OA21x2_ASAP7_75t_L g1905 ( 
.A1(n_1639),
.A2(n_1058),
.B(n_1049),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1559),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1689),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1559),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1650),
.Y(n_1909)
);

OAI22x1_ASAP7_75t_L g1910 ( 
.A1(n_1663),
.A2(n_1000),
.B1(n_1002),
.B2(n_1001),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1585),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1585),
.Y(n_1912)
);

HB1xp67_ASAP7_75t_L g1913 ( 
.A(n_1622),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1569),
.B(n_1004),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1585),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1801),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1720),
.Y(n_1917)
);

CKINVDCx16_ASAP7_75t_R g1918 ( 
.A(n_1749),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1818),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1815),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1803),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1722),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1864),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1818),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1720),
.Y(n_1925)
);

CKINVDCx20_ASAP7_75t_R g1926 ( 
.A(n_1856),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1750),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1883),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1752),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_SL g1930 ( 
.A(n_1913),
.B(n_1010),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1770),
.Y(n_1931)
);

CKINVDCx6p67_ASAP7_75t_R g1932 ( 
.A(n_1706),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_R g1933 ( 
.A(n_1838),
.B(n_1051),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1782),
.Y(n_1934)
);

AOI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1827),
.A2(n_1061),
.B(n_1059),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_R g1936 ( 
.A(n_1843),
.B(n_1070),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1784),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1893),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1827),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1787),
.Y(n_1940)
);

CKINVDCx20_ASAP7_75t_R g1941 ( 
.A(n_1863),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1706),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_R g1943 ( 
.A(n_1773),
.B(n_1788),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1693),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1806),
.B(n_1013),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1890),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1903),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1811),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1809),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1719),
.B(n_1066),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1789),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1854),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1711),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1819),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_R g1955 ( 
.A(n_1819),
.B(n_1079),
.Y(n_1955)
);

BUFx3_ASAP7_75t_L g1956 ( 
.A(n_1862),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1809),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1739),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1810),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1729),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1816),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1760),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_R g1963 ( 
.A(n_1781),
.B(n_1794),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1817),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1699),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1810),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1826),
.Y(n_1967)
);

CKINVDCx20_ASAP7_75t_R g1968 ( 
.A(n_1741),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1726),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1740),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1740),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1712),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_R g1973 ( 
.A(n_1825),
.B(n_1091),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1755),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1812),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1730),
.B(n_1019),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1745),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1779),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1797),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1802),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1697),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1745),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1698),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1708),
.B(n_1725),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1825),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1702),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1835),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1812),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1841),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1703),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1762),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1727),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1861),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1807),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1821),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1844),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1821),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1767),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1902),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1704),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1715),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1857),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1895),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1710),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_R g2005 ( 
.A(n_1724),
.B(n_1123),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1754),
.Y(n_2006)
);

CKINVDCx16_ASAP7_75t_R g2007 ( 
.A(n_1831),
.Y(n_2007)
);

CKINVDCx20_ASAP7_75t_R g2008 ( 
.A(n_1874),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1910),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1690),
.Y(n_2010)
);

NAND2xp33_ASAP7_75t_R g2011 ( 
.A(n_1823),
.B(n_1021),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1850),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1853),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1836),
.Y(n_2014)
);

CKINVDCx20_ASAP7_75t_R g2015 ( 
.A(n_1871),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1867),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1880),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1851),
.Y(n_2018)
);

INVx3_ASAP7_75t_L g2019 ( 
.A(n_1767),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1870),
.Y(n_2020)
);

CKINVDCx16_ASAP7_75t_R g2021 ( 
.A(n_1764),
.Y(n_2021)
);

BUFx2_ASAP7_75t_L g2022 ( 
.A(n_1869),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1833),
.Y(n_2023)
);

INVx8_ASAP7_75t_L g2024 ( 
.A(n_1763),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1858),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1808),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1873),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1875),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_R g2029 ( 
.A(n_1730),
.B(n_1128),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1884),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1771),
.Y(n_2031)
);

NOR2xp67_ASAP7_75t_L g2032 ( 
.A(n_1790),
.B(n_1799),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1891),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1896),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1876),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1900),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_R g2037 ( 
.A(n_1691),
.B(n_1138),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1798),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1881),
.Y(n_2039)
);

CKINVDCx20_ASAP7_75t_R g2040 ( 
.A(n_1822),
.Y(n_2040)
);

INVxp33_ASAP7_75t_SL g2041 ( 
.A(n_1692),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1696),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_1820),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1765),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1721),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1824),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1842),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1892),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1909),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1897),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1839),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1898),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_R g2053 ( 
.A(n_1694),
.B(n_1906),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1717),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1908),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_1728),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1813),
.Y(n_2057)
);

CKINVDCx16_ASAP7_75t_R g2058 ( 
.A(n_1723),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1830),
.Y(n_2059)
);

INVxp67_ASAP7_75t_L g2060 ( 
.A(n_1828),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1834),
.Y(n_2061)
);

CKINVDCx20_ASAP7_75t_R g2062 ( 
.A(n_1829),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_R g2063 ( 
.A(n_1709),
.B(n_1157),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_R g2064 ( 
.A(n_1866),
.B(n_1885),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1774),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_R g2066 ( 
.A(n_1888),
.B(n_1164),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1846),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_1914),
.Y(n_2068)
);

AO21x2_ASAP7_75t_L g2069 ( 
.A1(n_1785),
.A2(n_1074),
.B(n_1072),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1845),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_1780),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1847),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1852),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1855),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_R g2075 ( 
.A(n_1732),
.B(n_1211),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1865),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1776),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_R g2078 ( 
.A(n_1735),
.B(n_1254),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_1786),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_R g2080 ( 
.A(n_1736),
.B(n_1255),
.Y(n_2080)
);

INVxp33_ASAP7_75t_L g2081 ( 
.A(n_1731),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1877),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1878),
.Y(n_2083)
);

CKINVDCx20_ASAP7_75t_R g2084 ( 
.A(n_1695),
.Y(n_2084)
);

XNOR2xp5_ASAP7_75t_L g2085 ( 
.A(n_1860),
.B(n_1261),
.Y(n_2085)
);

INVx3_ASAP7_75t_L g2086 ( 
.A(n_1771),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1777),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1775),
.Y(n_2088)
);

CKINVDCx16_ASAP7_75t_R g2089 ( 
.A(n_1792),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1879),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1804),
.B(n_1023),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1882),
.Y(n_2092)
);

XNOR2xp5_ASAP7_75t_L g2093 ( 
.A(n_1796),
.B(n_1273),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1889),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1805),
.B(n_1108),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1894),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1775),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1783),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1911),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_R g2100 ( 
.A(n_1743),
.B(n_1292),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_R g2101 ( 
.A(n_1746),
.B(n_1295),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1783),
.Y(n_2102)
);

BUFx2_ASAP7_75t_L g2103 ( 
.A(n_1814),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1793),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1912),
.Y(n_2105)
);

BUFx10_ASAP7_75t_L g2106 ( 
.A(n_1747),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1915),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1695),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1832),
.Y(n_2109)
);

CKINVDCx5p33_ASAP7_75t_R g2110 ( 
.A(n_1832),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_R g2111 ( 
.A(n_1769),
.B(n_1298),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1772),
.B(n_1024),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1793),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_R g2114 ( 
.A(n_1766),
.B(n_1311),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1800),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1800),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1778),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1791),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_R g2119 ( 
.A(n_1766),
.B(n_1317),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_1840),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_1795),
.Y(n_2121)
);

INVx6_ASAP7_75t_L g2122 ( 
.A(n_1714),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_R g2123 ( 
.A(n_1766),
.B(n_1327),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_1848),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1768),
.Y(n_2125)
);

AOI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_1868),
.A2(n_1547),
.B1(n_1548),
.B2(n_1546),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_1768),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1872),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_1768),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_R g2130 ( 
.A(n_1886),
.B(n_1362),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1905),
.Y(n_2131)
);

CKINVDCx20_ASAP7_75t_R g2132 ( 
.A(n_1714),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_1886),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1886),
.Y(n_2134)
);

CKINVDCx20_ASAP7_75t_R g2135 ( 
.A(n_1718),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1718),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1738),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1734),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1734),
.Y(n_2139)
);

CKINVDCx20_ASAP7_75t_R g2140 ( 
.A(n_1737),
.Y(n_2140)
);

CKINVDCx5p33_ASAP7_75t_R g2141 ( 
.A(n_1737),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_1748),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1748),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1742),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_1756),
.Y(n_2145)
);

NAND2xp33_ASAP7_75t_R g2146 ( 
.A(n_1701),
.B(n_1025),
.Y(n_2146)
);

CKINVDCx20_ASAP7_75t_R g2147 ( 
.A(n_1756),
.Y(n_2147)
);

OAI22xp33_ASAP7_75t_L g2148 ( 
.A1(n_1744),
.A2(n_1408),
.B1(n_1428),
.B2(n_1389),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_1758),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_1758),
.Y(n_2150)
);

BUFx3_ASAP7_75t_L g2151 ( 
.A(n_1705),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1751),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_R g2153 ( 
.A(n_1716),
.B(n_1483),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1753),
.Y(n_2154)
);

XOR2xp5_ASAP7_75t_L g2155 ( 
.A(n_1757),
.B(n_1537),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1759),
.Y(n_2156)
);

BUFx2_ASAP7_75t_L g2157 ( 
.A(n_1761),
.Y(n_2157)
);

NOR2x1p5_ASAP7_75t_L g2158 ( 
.A(n_1733),
.B(n_1027),
.Y(n_2158)
);

CKINVDCx16_ASAP7_75t_R g2159 ( 
.A(n_1700),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_1700),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1707),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1707),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1713),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1713),
.Y(n_2164)
);

INVx3_ASAP7_75t_L g2165 ( 
.A(n_1837),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1837),
.Y(n_2166)
);

NAND2xp33_ASAP7_75t_R g2167 ( 
.A(n_1849),
.B(n_1028),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1849),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_1859),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1859),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_1887),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_1887),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_1899),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1899),
.Y(n_2174)
);

CKINVDCx16_ASAP7_75t_R g2175 ( 
.A(n_1901),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_R g2176 ( 
.A(n_1907),
.B(n_1514),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1901),
.Y(n_2177)
);

AOI21x1_ASAP7_75t_L g2178 ( 
.A1(n_1904),
.A2(n_1543),
.B(n_1540),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_1904),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1907),
.Y(n_2180)
);

CKINVDCx20_ASAP7_75t_R g2181 ( 
.A(n_1722),
.Y(n_2181)
);

CKINVDCx20_ASAP7_75t_R g2182 ( 
.A(n_1722),
.Y(n_2182)
);

BUFx3_ASAP7_75t_L g2183 ( 
.A(n_1862),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1801),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_1818),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_1801),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1720),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1801),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_1801),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1720),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1818),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1818),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1720),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1801),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1801),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_1801),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1801),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_1801),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_1883),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1720),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_1801),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_1818),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1720),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1720),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1818),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1801),
.Y(n_2206)
);

BUFx10_ASAP7_75t_L g2207 ( 
.A(n_1883),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_1883),
.Y(n_2208)
);

BUFx10_ASAP7_75t_L g2209 ( 
.A(n_1883),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1801),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_1801),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_1818),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_R g2213 ( 
.A(n_1750),
.B(n_1522),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1801),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_1883),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1818),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1818),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2044),
.B(n_1030),
.Y(n_2218)
);

BUFx3_ASAP7_75t_L g2219 ( 
.A(n_2008),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_1928),
.B(n_1534),
.Y(n_2220)
);

BUFx3_ASAP7_75t_L g2221 ( 
.A(n_2132),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2041),
.B(n_1038),
.Y(n_2222)
);

INVx5_ASAP7_75t_L g2223 ( 
.A(n_2207),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_2207),
.Y(n_2224)
);

OR2x2_ASAP7_75t_L g2225 ( 
.A(n_1967),
.B(n_990),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1983),
.Y(n_2226)
);

NAND2x1p5_ASAP7_75t_L g2227 ( 
.A(n_1956),
.B(n_1048),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2045),
.A2(n_2043),
.B1(n_2056),
.B2(n_2199),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_2209),
.B(n_2202),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1986),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_2021),
.B(n_1032),
.Y(n_2231)
);

AND2x4_ASAP7_75t_L g2232 ( 
.A(n_2208),
.B(n_1172),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1987),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_2209),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2004),
.B(n_1043),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2202),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1989),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_SL g2238 ( 
.A(n_2202),
.B(n_1044),
.Y(n_2238)
);

INVx4_ASAP7_75t_L g2239 ( 
.A(n_1932),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2215),
.B(n_1108),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1996),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2212),
.Y(n_2242)
);

BUFx4f_ASAP7_75t_L g2243 ( 
.A(n_2024),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2124),
.A2(n_1093),
.B(n_1081),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2212),
.Y(n_2245)
);

BUFx3_ASAP7_75t_L g2246 ( 
.A(n_2135),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1984),
.B(n_1046),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2029),
.B(n_1148),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2060),
.B(n_1053),
.Y(n_2249)
);

BUFx3_ASAP7_75t_L g2250 ( 
.A(n_2140),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2068),
.B(n_1054),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2012),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2013),
.Y(n_2253)
);

INVx3_ASAP7_75t_L g2254 ( 
.A(n_2159),
.Y(n_2254)
);

AND2x6_ASAP7_75t_L g2255 ( 
.A(n_2057),
.B(n_1095),
.Y(n_2255)
);

HB1xp67_ASAP7_75t_L g2256 ( 
.A(n_2153),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2212),
.B(n_1057),
.Y(n_2257)
);

INVx4_ASAP7_75t_L g2258 ( 
.A(n_1952),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2148),
.B(n_1257),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_1961),
.B(n_1964),
.Y(n_2260)
);

BUFx6f_ASAP7_75t_L g2261 ( 
.A(n_2183),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2032),
.B(n_1060),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2151),
.Y(n_2263)
);

NOR2x1p5_ASAP7_75t_L g2264 ( 
.A(n_1944),
.B(n_1549),
.Y(n_2264)
);

BUFx2_ASAP7_75t_L g2265 ( 
.A(n_1926),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1994),
.Y(n_2266)
);

AND2x6_ASAP7_75t_L g2267 ( 
.A(n_2016),
.B(n_1102),
.Y(n_2267)
);

INVx2_ASAP7_75t_SL g2268 ( 
.A(n_2024),
.Y(n_2268)
);

AND2x4_ASAP7_75t_L g2269 ( 
.A(n_1941),
.B(n_2095),
.Y(n_2269)
);

BUFx3_ASAP7_75t_L g2270 ( 
.A(n_1921),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1994),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2020),
.Y(n_2272)
);

BUFx10_ASAP7_75t_L g2273 ( 
.A(n_1920),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2027),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2106),
.B(n_1064),
.Y(n_2275)
);

INVx1_ASAP7_75t_SL g2276 ( 
.A(n_2176),
.Y(n_2276)
);

INVx1_ASAP7_75t_SL g2277 ( 
.A(n_2147),
.Y(n_2277)
);

OAI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_1978),
.A2(n_1553),
.B1(n_1552),
.B2(n_1069),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2035),
.Y(n_2279)
);

HB1xp67_ASAP7_75t_L g2280 ( 
.A(n_1946),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_2024),
.Y(n_2281)
);

BUFx3_ASAP7_75t_L g2282 ( 
.A(n_1916),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1935),
.Y(n_2283)
);

NOR2xp33_ASAP7_75t_SL g2284 ( 
.A(n_1979),
.B(n_1067),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2010),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_2184),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_2175),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2039),
.Y(n_2288)
);

INVx3_ASAP7_75t_L g2289 ( 
.A(n_2106),
.Y(n_2289)
);

OR2x6_ASAP7_75t_L g2290 ( 
.A(n_2022),
.B(n_1477),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2048),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_L g2292 ( 
.A(n_2007),
.B(n_1071),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_2046),
.B(n_1076),
.Y(n_2293)
);

NAND2xp33_ASAP7_75t_SL g2294 ( 
.A(n_1963),
.B(n_1535),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2050),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2052),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_1981),
.B(n_1078),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2157),
.B(n_1080),
.Y(n_2298)
);

OR2x6_ASAP7_75t_L g2299 ( 
.A(n_2185),
.B(n_1104),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2055),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1950),
.B(n_2118),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2042),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2065),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2077),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2087),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2051),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2117),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_2146),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2158),
.B(n_1301),
.Y(n_2309)
);

CKINVDCx16_ASAP7_75t_R g2310 ( 
.A(n_1955),
.Y(n_2310)
);

NAND2x1p5_ASAP7_75t_L g2311 ( 
.A(n_1919),
.B(n_1324),
.Y(n_2311)
);

BUFx2_ASAP7_75t_L g2312 ( 
.A(n_2075),
.Y(n_2312)
);

OR2x2_ASAP7_75t_L g2313 ( 
.A(n_2155),
.B(n_1342),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_1943),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2064),
.B(n_1082),
.Y(n_2315)
);

INVx3_ASAP7_75t_L g2316 ( 
.A(n_1919),
.Y(n_2316)
);

AND2x2_ASAP7_75t_SL g2317 ( 
.A(n_1918),
.B(n_1110),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2103),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_2070),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1950),
.B(n_1084),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2074),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_1980),
.B(n_1148),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2000),
.B(n_2001),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1924),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2082),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2078),
.B(n_1169),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2121),
.B(n_1085),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2191),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2058),
.B(n_1377),
.Y(n_2329)
);

INVxp67_ASAP7_75t_L g2330 ( 
.A(n_1930),
.Y(n_2330)
);

BUFx2_ASAP7_75t_L g2331 ( 
.A(n_2080),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_2028),
.B(n_1089),
.Y(n_2332)
);

INVx4_ASAP7_75t_L g2333 ( 
.A(n_2002),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2083),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_2186),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_1947),
.B(n_1387),
.Y(n_2336)
);

HB1xp67_ASAP7_75t_L g2337 ( 
.A(n_2100),
.Y(n_2337)
);

OR2x6_ASAP7_75t_L g2338 ( 
.A(n_1934),
.B(n_1937),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1976),
.B(n_1090),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2192),
.Y(n_2340)
);

BUFx10_ASAP7_75t_L g2341 ( 
.A(n_2188),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2091),
.B(n_1092),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2205),
.B(n_1097),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_SL g2344 ( 
.A(n_2053),
.B(n_1098),
.Y(n_2344)
);

BUFx3_ASAP7_75t_L g2345 ( 
.A(n_2189),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2094),
.Y(n_2346)
);

BUFx3_ASAP7_75t_L g2347 ( 
.A(n_2194),
.Y(n_2347)
);

OR2x6_ASAP7_75t_L g2348 ( 
.A(n_1940),
.B(n_1111),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2216),
.Y(n_2349)
);

BUFx10_ASAP7_75t_L g2350 ( 
.A(n_2195),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2099),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_L g2352 ( 
.A(n_2014),
.B(n_1099),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2105),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2217),
.B(n_1100),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1965),
.Y(n_2355)
);

INVx3_ASAP7_75t_L g2356 ( 
.A(n_2090),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2137),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2144),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2126),
.B(n_1101),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2152),
.Y(n_2360)
);

BUFx2_ASAP7_75t_L g2361 ( 
.A(n_2101),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_2196),
.Y(n_2362)
);

INVx8_ASAP7_75t_L g2363 ( 
.A(n_2003),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1948),
.B(n_1103),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2197),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2154),
.Y(n_2366)
);

INVx1_ASAP7_75t_SL g2367 ( 
.A(n_2111),
.Y(n_2367)
);

NAND3xp33_ASAP7_75t_L g2368 ( 
.A(n_2017),
.B(n_1109),
.C(n_1107),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2112),
.B(n_1112),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_1917),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2066),
.B(n_1169),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2142),
.B(n_1114),
.Y(n_2372)
);

INVx4_ASAP7_75t_L g2373 ( 
.A(n_1942),
.Y(n_2373)
);

OR2x6_ASAP7_75t_L g2374 ( 
.A(n_1945),
.B(n_1113),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1925),
.Y(n_2375)
);

OAI22xp33_ASAP7_75t_L g2376 ( 
.A1(n_2025),
.A2(n_1529),
.B1(n_1538),
.B2(n_1528),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2156),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_1939),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_1953),
.B(n_1117),
.Y(n_2379)
);

NAND3x1_ASAP7_75t_L g2380 ( 
.A(n_2198),
.B(n_1116),
.C(n_1115),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2187),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1960),
.Y(n_2382)
);

OR2x6_ASAP7_75t_L g2383 ( 
.A(n_2201),
.B(n_1120),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1962),
.Y(n_2384)
);

INVx5_ASAP7_75t_L g2385 ( 
.A(n_2089),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2063),
.B(n_1200),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2069),
.B(n_1118),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_1927),
.B(n_1393),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2069),
.B(n_1119),
.Y(n_2389)
);

AND2x4_ASAP7_75t_L g2390 ( 
.A(n_1985),
.B(n_1407),
.Y(n_2390)
);

AOI22xp33_ASAP7_75t_L g2391 ( 
.A1(n_2079),
.A2(n_1130),
.B1(n_1131),
.B2(n_1122),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2190),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2193),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2200),
.Y(n_2394)
);

BUFx2_ASAP7_75t_L g2395 ( 
.A(n_2037),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_1958),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2093),
.B(n_1200),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2005),
.B(n_1215),
.Y(n_2398)
);

BUFx3_ASAP7_75t_L g2399 ( 
.A(n_2214),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2072),
.B(n_1124),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_SL g2401 ( 
.A(n_1954),
.B(n_1125),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2038),
.B(n_1215),
.Y(n_2402)
);

INVx5_ASAP7_75t_L g2403 ( 
.A(n_2122),
.Y(n_2403)
);

OAI22xp5_ASAP7_75t_SL g2404 ( 
.A1(n_1923),
.A2(n_1127),
.B1(n_1129),
.B2(n_1126),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2073),
.B(n_1134),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2203),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2204),
.Y(n_2407)
);

AND2x6_ASAP7_75t_L g2408 ( 
.A(n_2128),
.B(n_1132),
.Y(n_2408)
);

INVx6_ASAP7_75t_L g2409 ( 
.A(n_2206),
.Y(n_2409)
);

INVx5_ASAP7_75t_L g2410 ( 
.A(n_2122),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2143),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2210),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_1991),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2145),
.Y(n_2414)
);

INVx1_ASAP7_75t_SL g2415 ( 
.A(n_1933),
.Y(n_2415)
);

AND2x6_ASAP7_75t_L g2416 ( 
.A(n_1998),
.B(n_1140),
.Y(n_2416)
);

OR2x6_ASAP7_75t_L g2417 ( 
.A(n_2211),
.B(n_1143),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2149),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2178),
.Y(n_2419)
);

AND2x4_ASAP7_75t_L g2420 ( 
.A(n_1929),
.B(n_1419),
.Y(n_2420)
);

AND2x6_ASAP7_75t_L g2421 ( 
.A(n_1998),
.B(n_1145),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2030),
.B(n_1137),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2033),
.B(n_1152),
.Y(n_2423)
);

BUFx3_ASAP7_75t_L g2424 ( 
.A(n_2084),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_SL g2425 ( 
.A(n_2181),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_1949),
.Y(n_2426)
);

INVx4_ASAP7_75t_L g2427 ( 
.A(n_2136),
.Y(n_2427)
);

AND2x6_ASAP7_75t_L g2428 ( 
.A(n_2019),
.B(n_1146),
.Y(n_2428)
);

INVx1_ASAP7_75t_SL g2429 ( 
.A(n_1936),
.Y(n_2429)
);

INVx4_ASAP7_75t_L g2430 ( 
.A(n_2138),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2150),
.Y(n_2431)
);

OAI22xp33_ASAP7_75t_L g2432 ( 
.A1(n_2026),
.A2(n_1521),
.B1(n_1541),
.B2(n_1519),
.Y(n_2432)
);

INVx4_ASAP7_75t_L g2433 ( 
.A(n_2139),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1970),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2076),
.B(n_1147),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2161),
.Y(n_2436)
);

XOR2x2_ASAP7_75t_SL g2437 ( 
.A(n_2213),
.B(n_1238),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_1971),
.Y(n_2438)
);

BUFx2_ASAP7_75t_L g2439 ( 
.A(n_1973),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1977),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_1957),
.Y(n_2441)
);

INVx4_ASAP7_75t_L g2442 ( 
.A(n_2141),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2092),
.B(n_1158),
.Y(n_2443)
);

AOI22xp33_ASAP7_75t_L g2444 ( 
.A1(n_2120),
.A2(n_1153),
.B1(n_1154),
.B2(n_1151),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2018),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2034),
.B(n_2006),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_1982),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2062),
.B(n_1238),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_1959),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2088),
.Y(n_2450)
);

BUFx3_ASAP7_75t_L g2451 ( 
.A(n_1931),
.Y(n_2451)
);

NAND2x1p5_ASAP7_75t_L g2452 ( 
.A(n_2019),
.B(n_1452),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2097),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2114),
.B(n_1161),
.Y(n_2454)
);

BUFx4f_ASAP7_75t_L g2455 ( 
.A(n_1938),
.Y(n_2455)
);

BUFx2_ASAP7_75t_L g2456 ( 
.A(n_1990),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2098),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2096),
.B(n_1163),
.Y(n_2458)
);

AND2x4_ASAP7_75t_L g2459 ( 
.A(n_2015),
.B(n_1459),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2102),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2104),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2107),
.B(n_1166),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2113),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2115),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_1969),
.B(n_1241),
.Y(n_2465)
);

BUFx6f_ASAP7_75t_L g2466 ( 
.A(n_2163),
.Y(n_2466)
);

AOI22xp33_ASAP7_75t_L g2467 ( 
.A1(n_2131),
.A2(n_1160),
.B1(n_1162),
.B2(n_1155),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2061),
.B(n_1171),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2031),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_1966),
.Y(n_2470)
);

AND2x6_ASAP7_75t_L g2471 ( 
.A(n_2031),
.B(n_1167),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_1975),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_1988),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2086),
.Y(n_2474)
);

OR2x2_ASAP7_75t_L g2475 ( 
.A(n_1922),
.B(n_1177),
.Y(n_2475)
);

BUFx10_ASAP7_75t_L g2476 ( 
.A(n_1995),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2086),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_2067),
.B(n_1178),
.Y(n_2478)
);

HB1xp67_ASAP7_75t_L g2479 ( 
.A(n_2167),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2116),
.Y(n_2480)
);

CKINVDCx11_ASAP7_75t_R g2481 ( 
.A(n_2182),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2108),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_L g2483 ( 
.A(n_2054),
.B(n_1179),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2160),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2109),
.Y(n_2485)
);

INVx2_ASAP7_75t_SL g2486 ( 
.A(n_2059),
.Y(n_2486)
);

AND2x4_ASAP7_75t_L g2487 ( 
.A(n_2071),
.B(n_1168),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2119),
.B(n_1182),
.Y(n_2488)
);

HB1xp67_ASAP7_75t_L g2489 ( 
.A(n_2123),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2160),
.Y(n_2490)
);

OR2x2_ASAP7_75t_L g2491 ( 
.A(n_2085),
.B(n_1186),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2110),
.Y(n_2492)
);

AND2x6_ASAP7_75t_L g2493 ( 
.A(n_2130),
.B(n_1170),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2165),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2081),
.Y(n_2495)
);

INVx5_ASAP7_75t_L g2496 ( 
.A(n_2165),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2168),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2174),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2171),
.Y(n_2499)
);

NAND2x1p5_ASAP7_75t_L g2500 ( 
.A(n_2047),
.B(n_1175),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2036),
.B(n_2049),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_1951),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2174),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_1972),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_1999),
.B(n_1241),
.Y(n_2505)
);

BUFx3_ASAP7_75t_L g2506 ( 
.A(n_2172),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2125),
.B(n_1187),
.Y(n_2507)
);

NAND2x1p5_ASAP7_75t_L g2508 ( 
.A(n_1997),
.B(n_1180),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2173),
.Y(n_2509)
);

INVx4_ASAP7_75t_L g2510 ( 
.A(n_2179),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2040),
.B(n_1193),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_1993),
.B(n_1196),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2133),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2169),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2162),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2009),
.A2(n_1184),
.B1(n_1188),
.B2(n_1183),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2127),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2129),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2134),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_1992),
.Y(n_2520)
);

BUFx10_ASAP7_75t_L g2521 ( 
.A(n_1974),
.Y(n_2521)
);

AND2x6_ASAP7_75t_L g2522 ( 
.A(n_2011),
.B(n_1192),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2023),
.B(n_1197),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_1968),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_SL g2525 ( 
.A(n_2164),
.B(n_1198),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2166),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2170),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2177),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2180),
.B(n_1309),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_1928),
.B(n_1195),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2041),
.B(n_1203),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_1983),
.Y(n_2532)
);

OR2x2_ASAP7_75t_L g2533 ( 
.A(n_1967),
.B(n_1205),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2044),
.B(n_1206),
.Y(n_2534)
);

AND2x4_ASAP7_75t_L g2535 ( 
.A(n_1928),
.B(n_1199),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_1983),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2202),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2207),
.B(n_1208),
.Y(n_2538)
);

AND2x4_ASAP7_75t_L g2539 ( 
.A(n_1928),
.B(n_1201),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2044),
.B(n_1210),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_L g2541 ( 
.A(n_2041),
.B(n_1212),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2207),
.Y(n_2542)
);

BUFx6f_ASAP7_75t_L g2543 ( 
.A(n_2202),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_1928),
.B(n_1309),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_L g2545 ( 
.A(n_2202),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_1928),
.B(n_1421),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_1967),
.B(n_1214),
.Y(n_2547)
);

INVx4_ASAP7_75t_L g2548 ( 
.A(n_1932),
.Y(n_2548)
);

INVxp67_ASAP7_75t_L g2549 ( 
.A(n_1928),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_1983),
.Y(n_2550)
);

BUFx6f_ASAP7_75t_L g2551 ( 
.A(n_2202),
.Y(n_2551)
);

INVx2_ASAP7_75t_SL g2552 ( 
.A(n_2207),
.Y(n_2552)
);

NAND3xp33_ASAP7_75t_L g2553 ( 
.A(n_2045),
.B(n_1217),
.C(n_1216),
.Y(n_2553)
);

BUFx6f_ASAP7_75t_L g2554 ( 
.A(n_2202),
.Y(n_2554)
);

OR2x2_ASAP7_75t_L g2555 ( 
.A(n_1967),
.B(n_1218),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2008),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2044),
.B(n_1221),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2202),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_1983),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_1983),
.Y(n_2560)
);

INVxp67_ASAP7_75t_L g2561 ( 
.A(n_1928),
.Y(n_2561)
);

AND2x4_ASAP7_75t_L g2562 ( 
.A(n_1928),
.B(n_1202),
.Y(n_2562)
);

AOI22xp5_ASAP7_75t_L g2563 ( 
.A1(n_2041),
.A2(n_1222),
.B1(n_1229),
.B2(n_1226),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_1983),
.Y(n_2564)
);

INVx4_ASAP7_75t_L g2565 ( 
.A(n_1932),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2044),
.B(n_1234),
.Y(n_2566)
);

BUFx6f_ASAP7_75t_L g2567 ( 
.A(n_2202),
.Y(n_2567)
);

AND2x6_ASAP7_75t_L g2568 ( 
.A(n_2057),
.B(n_1209),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2044),
.B(n_1236),
.Y(n_2569)
);

INVx4_ASAP7_75t_L g2570 ( 
.A(n_1932),
.Y(n_2570)
);

AOI21x1_ASAP7_75t_L g2571 ( 
.A1(n_1935),
.A2(n_1227),
.B(n_1224),
.Y(n_2571)
);

CKINVDCx20_ASAP7_75t_R g2572 ( 
.A(n_1926),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1983),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_SL g2574 ( 
.A(n_2207),
.B(n_1237),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_1983),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_1921),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2044),
.B(n_1243),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_1983),
.Y(n_2578)
);

BUFx3_ASAP7_75t_L g2579 ( 
.A(n_2008),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_1928),
.B(n_1421),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1983),
.Y(n_2581)
);

INVx1_ASAP7_75t_SL g2582 ( 
.A(n_2207),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2207),
.B(n_1244),
.Y(n_2583)
);

AND2x4_ASAP7_75t_L g2584 ( 
.A(n_1928),
.B(n_1228),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_1983),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2044),
.B(n_1245),
.Y(n_2586)
);

INVx4_ASAP7_75t_L g2587 ( 
.A(n_1932),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2202),
.Y(n_2588)
);

BUFx3_ASAP7_75t_L g2589 ( 
.A(n_2008),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2202),
.Y(n_2590)
);

INVxp67_ASAP7_75t_SL g2591 ( 
.A(n_1928),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2044),
.B(n_1246),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2202),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_SL g2594 ( 
.A(n_1944),
.B(n_1247),
.Y(n_2594)
);

AO22x2_ASAP7_75t_L g2595 ( 
.A1(n_2155),
.A2(n_1239),
.B1(n_1240),
.B2(n_1233),
.Y(n_2595)
);

AND2x4_ASAP7_75t_L g2596 ( 
.A(n_1928),
.B(n_1242),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2413),
.Y(n_2597)
);

INVxp67_ASAP7_75t_L g2598 ( 
.A(n_2591),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_2289),
.B(n_1249),
.Y(n_2599)
);

NAND2x1p5_ASAP7_75t_L g2600 ( 
.A(n_2223),
.B(n_989),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2226),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2230),
.Y(n_2602)
);

OR2x2_ASAP7_75t_SL g2603 ( 
.A(n_2310),
.B(n_1251),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2393),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_2481),
.Y(n_2605)
);

INVx2_ASAP7_75t_SL g2606 ( 
.A(n_2223),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2233),
.Y(n_2607)
);

OR2x2_ASAP7_75t_L g2608 ( 
.A(n_2277),
.B(n_1250),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_SL g2609 ( 
.A(n_2224),
.B(n_1550),
.Y(n_2609)
);

A2O1A1Ixp33_ASAP7_75t_L g2610 ( 
.A1(n_2244),
.A2(n_1258),
.B(n_1265),
.C(n_1253),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_SL g2611 ( 
.A(n_2582),
.B(n_1252),
.Y(n_2611)
);

NAND3x1_ASAP7_75t_L g2612 ( 
.A(n_2228),
.B(n_1525),
.C(n_1515),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2237),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2241),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2252),
.Y(n_2615)
);

NAND2x1p5_ASAP7_75t_L g2616 ( 
.A(n_2243),
.B(n_989),
.Y(n_2616)
);

NAND3xp33_ASAP7_75t_L g2617 ( 
.A(n_2332),
.B(n_992),
.C(n_989),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2552),
.B(n_1266),
.Y(n_2618)
);

OR2x6_ASAP7_75t_SL g2619 ( 
.A(n_2314),
.B(n_1256),
.Y(n_2619)
);

A2O1A1Ixp33_ASAP7_75t_L g2620 ( 
.A1(n_2253),
.A2(n_1278),
.B(n_1285),
.C(n_1268),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2284),
.B(n_1260),
.Y(n_2621)
);

AND2x4_ASAP7_75t_L g2622 ( 
.A(n_2234),
.B(n_1287),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2394),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2406),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2272),
.Y(n_2625)
);

BUFx6f_ASAP7_75t_L g2626 ( 
.A(n_2543),
.Y(n_2626)
);

BUFx3_ASAP7_75t_L g2627 ( 
.A(n_2363),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2274),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2279),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2288),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2301),
.B(n_1262),
.Y(n_2631)
);

AO22x2_ASAP7_75t_L g2632 ( 
.A1(n_2367),
.A2(n_2259),
.B1(n_2276),
.B2(n_2397),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2291),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2295),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2296),
.Y(n_2635)
);

AND2x4_ASAP7_75t_L g2636 ( 
.A(n_2542),
.B(n_1290),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2300),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2532),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2536),
.Y(n_2639)
);

OR2x2_ASAP7_75t_SL g2640 ( 
.A(n_2260),
.B(n_1296),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2247),
.B(n_1264),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2550),
.Y(n_2642)
);

AND2x4_ASAP7_75t_L g2643 ( 
.A(n_2333),
.B(n_1304),
.Y(n_2643)
);

BUFx8_ASAP7_75t_L g2644 ( 
.A(n_2425),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2407),
.Y(n_2645)
);

NAND3x1_ASAP7_75t_L g2646 ( 
.A(n_2437),
.B(n_1512),
.C(n_1511),
.Y(n_2646)
);

NAND3x1_ASAP7_75t_L g2647 ( 
.A(n_2520),
.B(n_1530),
.C(n_1527),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_SL g2648 ( 
.A(n_2549),
.B(n_1509),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2559),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2560),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2338),
.B(n_1307),
.Y(n_2651)
);

AND2x4_ASAP7_75t_L g2652 ( 
.A(n_2338),
.B(n_1312),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2564),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2573),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2575),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2578),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2267),
.B(n_1269),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2581),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2585),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2267),
.B(n_2561),
.Y(n_2660)
);

INVx6_ASAP7_75t_L g2661 ( 
.A(n_2273),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2303),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2304),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2370),
.Y(n_2664)
);

AO22x2_ASAP7_75t_L g2665 ( 
.A1(n_2415),
.A2(n_1326),
.B1(n_1328),
.B2(n_1315),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2220),
.B(n_1524),
.Y(n_2666)
);

AO22x2_ASAP7_75t_L g2667 ( 
.A1(n_2429),
.A2(n_1332),
.B1(n_1335),
.B2(n_1330),
.Y(n_2667)
);

OAI221xp5_ASAP7_75t_L g2668 ( 
.A1(n_2516),
.A2(n_1272),
.B1(n_1274),
.B2(n_1271),
.C(n_1270),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2305),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2375),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2307),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2357),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2358),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2378),
.Y(n_2674)
);

AND2x4_ASAP7_75t_L g2675 ( 
.A(n_2299),
.B(n_1337),
.Y(n_2675)
);

AND2x4_ASAP7_75t_L g2676 ( 
.A(n_2299),
.B(n_1344),
.Y(n_2676)
);

AND2x4_ASAP7_75t_L g2677 ( 
.A(n_2239),
.B(n_1346),
.Y(n_2677)
);

AOI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2222),
.A2(n_2541),
.B1(n_2531),
.B2(n_2594),
.Y(n_2678)
);

INVxp67_ASAP7_75t_L g2679 ( 
.A(n_2267),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2381),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2392),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_L g2682 ( 
.A(n_2512),
.B(n_1275),
.Y(n_2682)
);

BUFx8_ASAP7_75t_L g2683 ( 
.A(n_2265),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2360),
.Y(n_2684)
);

AOI22xp33_ASAP7_75t_L g2685 ( 
.A1(n_2522),
.A2(n_1539),
.B1(n_1524),
.B2(n_1279),
.Y(n_2685)
);

OAI21xp33_ASAP7_75t_L g2686 ( 
.A1(n_2249),
.A2(n_1280),
.B(n_1277),
.Y(n_2686)
);

NAND2x1p5_ASAP7_75t_L g2687 ( 
.A(n_2548),
.B(n_989),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2572),
.Y(n_2688)
);

AND2x4_ASAP7_75t_L g2689 ( 
.A(n_2565),
.B(n_1350),
.Y(n_2689)
);

NAND2xp33_ASAP7_75t_L g2690 ( 
.A(n_2255),
.B(n_1551),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2391),
.B(n_1281),
.Y(n_2691)
);

OAI22xp5_ASAP7_75t_SL g2692 ( 
.A1(n_2317),
.A2(n_1284),
.B1(n_1288),
.B2(n_1283),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2366),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2377),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2374),
.B(n_1289),
.Y(n_2695)
);

AND2x2_ASAP7_75t_SL g2696 ( 
.A(n_2455),
.B(n_1545),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2318),
.Y(n_2697)
);

AO22x2_ASAP7_75t_L g2698 ( 
.A1(n_2309),
.A2(n_1361),
.B1(n_1364),
.B2(n_1353),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2382),
.Y(n_2699)
);

NAND2x1p5_ASAP7_75t_L g2700 ( 
.A(n_2570),
.B(n_992),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2255),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2384),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2374),
.B(n_1291),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2266),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2355),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2285),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2444),
.B(n_1293),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_L g2708 ( 
.A(n_2511),
.B(n_1297),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2467),
.B(n_1299),
.Y(n_2709)
);

NOR3xp33_ASAP7_75t_L g2710 ( 
.A(n_2293),
.B(n_1533),
.C(n_1532),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2302),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2306),
.Y(n_2712)
);

AO22x2_ASAP7_75t_L g2713 ( 
.A1(n_2313),
.A2(n_2225),
.B1(n_2459),
.B2(n_2308),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2232),
.B(n_1302),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2271),
.Y(n_2715)
);

NAND2x1p5_ASAP7_75t_L g2716 ( 
.A(n_2587),
.B(n_992),
.Y(n_2716)
);

NAND3xp33_ASAP7_75t_L g2717 ( 
.A(n_2248),
.B(n_1149),
.C(n_992),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_2401),
.B(n_1544),
.Y(n_2718)
);

INVxp67_ASAP7_75t_L g2719 ( 
.A(n_2280),
.Y(n_2719)
);

HB1xp67_ASAP7_75t_L g2720 ( 
.A(n_2221),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2321),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2325),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2334),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2522),
.B(n_1303),
.Y(n_2724)
);

AND2x4_ASAP7_75t_L g2725 ( 
.A(n_2275),
.B(n_1367),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_L g2726 ( 
.A(n_2269),
.B(n_1306),
.Y(n_2726)
);

NAND2x1p5_ASAP7_75t_L g2727 ( 
.A(n_2385),
.B(n_2436),
.Y(n_2727)
);

INVx4_ASAP7_75t_L g2728 ( 
.A(n_2363),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2346),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2522),
.B(n_1308),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2351),
.Y(n_2731)
);

AND3x1_ASAP7_75t_L g2732 ( 
.A(n_2396),
.B(n_1382),
.C(n_1374),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2353),
.Y(n_2733)
);

AO22x2_ASAP7_75t_L g2734 ( 
.A1(n_2336),
.A2(n_1386),
.B1(n_1392),
.B2(n_1384),
.Y(n_2734)
);

AOI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2231),
.A2(n_2448),
.B1(n_2352),
.B2(n_2446),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2324),
.Y(n_2736)
);

AND2x4_ASAP7_75t_L g2737 ( 
.A(n_2445),
.B(n_1396),
.Y(n_2737)
);

INVxp67_ASAP7_75t_L g2738 ( 
.A(n_2256),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2385),
.B(n_1397),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2328),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2340),
.Y(n_2741)
);

INVx3_ASAP7_75t_L g2742 ( 
.A(n_2436),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2349),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2529),
.Y(n_2744)
);

AOI22x1_ASAP7_75t_L g2745 ( 
.A1(n_2419),
.A2(n_1416),
.B1(n_1420),
.B2(n_1406),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2263),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2255),
.B(n_1316),
.Y(n_2747)
);

BUFx4f_ASAP7_75t_L g2748 ( 
.A(n_2409),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2343),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2500),
.B(n_2595),
.Y(n_2750)
);

INVx1_ASAP7_75t_SL g2751 ( 
.A(n_2246),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2330),
.B(n_1425),
.Y(n_2752)
);

OAI22xp5_ASAP7_75t_L g2753 ( 
.A1(n_2348),
.A2(n_1319),
.B1(n_1320),
.B2(n_1318),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2595),
.B(n_1539),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2354),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2543),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_SL g2757 ( 
.A(n_2278),
.B(n_1496),
.Y(n_2757)
);

AOI22xp5_ASAP7_75t_L g2758 ( 
.A1(n_2297),
.A2(n_1325),
.B1(n_1329),
.B2(n_1322),
.Y(n_2758)
);

INVx3_ASAP7_75t_L g2759 ( 
.A(n_2466),
.Y(n_2759)
);

INVxp67_ASAP7_75t_L g2760 ( 
.A(n_2533),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2545),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2545),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2551),
.Y(n_2763)
);

CKINVDCx5p33_ASAP7_75t_R g2764 ( 
.A(n_2576),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2294),
.B(n_1503),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_R g2766 ( 
.A(n_2362),
.B(n_1331),
.Y(n_2766)
);

NAND2xp33_ASAP7_75t_L g2767 ( 
.A(n_2568),
.B(n_1508),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2551),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2554),
.Y(n_2769)
);

AND2x4_ASAP7_75t_L g2770 ( 
.A(n_2348),
.B(n_1430),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2554),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2387),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2568),
.B(n_1334),
.Y(n_2773)
);

NOR2xp33_ASAP7_75t_L g2774 ( 
.A(n_2505),
.B(n_1336),
.Y(n_2774)
);

AO22x2_ASAP7_75t_L g2775 ( 
.A1(n_2388),
.A2(n_1436),
.B1(n_1443),
.B2(n_1431),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2568),
.B(n_1338),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2218),
.B(n_1339),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_SL g2778 ( 
.A(n_2312),
.B(n_2331),
.Y(n_2778)
);

OAI221xp5_ASAP7_75t_L g2779 ( 
.A1(n_2320),
.A2(n_1343),
.B1(n_1354),
.B2(n_1341),
.C(n_1340),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2547),
.B(n_1355),
.Y(n_2780)
);

NAND2x1p5_ASAP7_75t_L g2781 ( 
.A(n_2466),
.B(n_1149),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2389),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2567),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2364),
.Y(n_2784)
);

NAND2xp33_ASAP7_75t_L g2785 ( 
.A(n_2408),
.B(n_1504),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2379),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_2361),
.B(n_1501),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2534),
.B(n_1358),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2567),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2311),
.Y(n_2790)
);

AO22x2_ASAP7_75t_L g2791 ( 
.A1(n_2491),
.A2(n_1449),
.B1(n_1451),
.B2(n_1444),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2236),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2242),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2540),
.B(n_1359),
.Y(n_2794)
);

AO22x2_ASAP7_75t_L g2795 ( 
.A1(n_2398),
.A2(n_1465),
.B1(n_1467),
.B2(n_1454),
.Y(n_2795)
);

BUFx3_ASAP7_75t_L g2796 ( 
.A(n_2261),
.Y(n_2796)
);

AO22x2_ASAP7_75t_L g2797 ( 
.A1(n_2390),
.A2(n_1478),
.B1(n_1481),
.B2(n_1475),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2452),
.Y(n_2798)
);

CKINVDCx16_ASAP7_75t_R g2799 ( 
.A(n_2270),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2434),
.Y(n_2800)
);

NOR3xp33_ASAP7_75t_L g2801 ( 
.A(n_2315),
.B(n_1507),
.C(n_1502),
.Y(n_2801)
);

BUFx2_ASAP7_75t_L g2802 ( 
.A(n_2250),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2245),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2438),
.Y(n_2804)
);

NOR3xp33_ASAP7_75t_L g2805 ( 
.A(n_2337),
.B(n_1484),
.C(n_1482),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2557),
.B(n_1360),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2440),
.Y(n_2807)
);

NOR2xp33_ASAP7_75t_L g2808 ( 
.A(n_2555),
.B(n_1363),
.Y(n_2808)
);

AND2x4_ASAP7_75t_L g2809 ( 
.A(n_2319),
.B(n_1486),
.Y(n_2809)
);

AND2x4_ASAP7_75t_L g2810 ( 
.A(n_2356),
.B(n_1489),
.Y(n_2810)
);

AND2x4_ASAP7_75t_L g2811 ( 
.A(n_2268),
.B(n_1),
.Y(n_2811)
);

INVxp67_ASAP7_75t_L g2812 ( 
.A(n_2456),
.Y(n_2812)
);

OR2x2_ASAP7_75t_L g2813 ( 
.A(n_2329),
.B(n_1365),
.Y(n_2813)
);

NAND2x1p5_ASAP7_75t_L g2814 ( 
.A(n_2254),
.B(n_1149),
.Y(n_2814)
);

INVxp67_ASAP7_75t_L g2815 ( 
.A(n_2439),
.Y(n_2815)
);

NAND3xp33_ASAP7_75t_L g2816 ( 
.A(n_2326),
.B(n_1174),
.C(n_1149),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2537),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2447),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2558),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2450),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2453),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2457),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_SL g2823 ( 
.A(n_2341),
.Y(n_2823)
);

AOI211xp5_ASAP7_75t_L g2824 ( 
.A1(n_2404),
.A2(n_1368),
.B(n_1369),
.C(n_1366),
.Y(n_2824)
);

OR2x2_ASAP7_75t_SL g2825 ( 
.A(n_2479),
.B(n_1545),
.Y(n_2825)
);

AOI22xp5_ASAP7_75t_L g2826 ( 
.A1(n_2235),
.A2(n_1371),
.B1(n_1372),
.B2(n_1370),
.Y(n_2826)
);

NAND2x1p5_ASAP7_75t_L g2827 ( 
.A(n_2287),
.B(n_1174),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2460),
.Y(n_2828)
);

INVxp67_ASAP7_75t_L g2829 ( 
.A(n_2451),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2461),
.Y(n_2830)
);

CKINVDCx20_ASAP7_75t_R g2831 ( 
.A(n_2412),
.Y(n_2831)
);

OAI22xp5_ASAP7_75t_SL g2832 ( 
.A1(n_2383),
.A2(n_1490),
.B1(n_1493),
.B2(n_1488),
.Y(n_2832)
);

INVxp67_ASAP7_75t_L g2833 ( 
.A(n_2420),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2463),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_2350),
.Y(n_2835)
);

AOI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_2530),
.A2(n_1378),
.B1(n_1379),
.B2(n_1373),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2464),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2566),
.B(n_1380),
.Y(n_2838)
);

CKINVDCx20_ASAP7_75t_R g2839 ( 
.A(n_2219),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2535),
.Y(n_2840)
);

NOR3xp33_ASAP7_75t_L g2841 ( 
.A(n_2402),
.B(n_1388),
.C(n_1381),
.Y(n_2841)
);

A2O1A1Ixp33_ASAP7_75t_L g2842 ( 
.A1(n_2369),
.A2(n_2339),
.B(n_2342),
.C(n_2359),
.Y(n_2842)
);

BUFx3_ASAP7_75t_L g2843 ( 
.A(n_2261),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2569),
.B(n_1390),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2539),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2562),
.Y(n_2846)
);

A2O1A1Ixp33_ASAP7_75t_L g2847 ( 
.A1(n_2262),
.A2(n_1220),
.B(n_1300),
.C(n_1174),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_SL g2848 ( 
.A(n_2323),
.B(n_1391),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2588),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2584),
.Y(n_2850)
);

AO22x2_ASAP7_75t_L g2851 ( 
.A1(n_2386),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_SL g2852 ( 
.A(n_2508),
.B(n_2577),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2586),
.B(n_1394),
.Y(n_2853)
);

INVxp33_ASAP7_75t_L g2854 ( 
.A(n_2292),
.Y(n_2854)
);

OR2x2_ASAP7_75t_L g2855 ( 
.A(n_2592),
.B(n_1395),
.Y(n_2855)
);

INVxp67_ASAP7_75t_L g2856 ( 
.A(n_2227),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2596),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2590),
.Y(n_2858)
);

INVxp67_ASAP7_75t_L g2859 ( 
.A(n_2493),
.Y(n_2859)
);

NAND2x1p5_ASAP7_75t_L g2860 ( 
.A(n_2427),
.B(n_1174),
.Y(n_2860)
);

AOI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2422),
.A2(n_1401),
.B1(n_1402),
.B2(n_1398),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2593),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2571),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2514),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2298),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2416),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2416),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_2432),
.B(n_2376),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2416),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2421),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2421),
.Y(n_2871)
);

INVxp67_ASAP7_75t_SL g2872 ( 
.A(n_2506),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2528),
.Y(n_2873)
);

AND2x4_ASAP7_75t_L g2874 ( 
.A(n_2281),
.B(n_2),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2251),
.B(n_1404),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2421),
.Y(n_2876)
);

AO22x2_ASAP7_75t_L g2877 ( 
.A1(n_2371),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2428),
.Y(n_2878)
);

BUFx6f_ASAP7_75t_L g2879 ( 
.A(n_2424),
.Y(n_2879)
);

CKINVDCx20_ASAP7_75t_R g2880 ( 
.A(n_2556),
.Y(n_2880)
);

INVxp67_ASAP7_75t_L g2881 ( 
.A(n_2493),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2426),
.Y(n_2882)
);

OR2x6_ASAP7_75t_L g2883 ( 
.A(n_2258),
.B(n_2290),
.Y(n_2883)
);

INVxp67_ASAP7_75t_L g2884 ( 
.A(n_2493),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2428),
.Y(n_2885)
);

AND2x2_ASAP7_75t_SL g2886 ( 
.A(n_2395),
.B(n_1545),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2428),
.Y(n_2887)
);

A2O1A1Ixp33_ASAP7_75t_L g2888 ( 
.A1(n_2283),
.A2(n_1300),
.B(n_1321),
.C(n_1220),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2441),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2471),
.Y(n_2890)
);

AND2x4_ASAP7_75t_L g2891 ( 
.A(n_2510),
.B(n_3),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2471),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2449),
.Y(n_2893)
);

AND2x4_ASAP7_75t_L g2894 ( 
.A(n_2482),
.B(n_5),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2471),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2470),
.Y(n_2896)
);

INVxp67_ASAP7_75t_L g2897 ( 
.A(n_2240),
.Y(n_2897)
);

NAND2xp33_ASAP7_75t_L g2898 ( 
.A(n_2408),
.B(n_1505),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_SL g2899 ( 
.A(n_2327),
.B(n_1497),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2472),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2473),
.Y(n_2901)
);

INVxp67_ASAP7_75t_L g2902 ( 
.A(n_2544),
.Y(n_2902)
);

NOR2xp33_ASAP7_75t_L g2903 ( 
.A(n_2465),
.B(n_1409),
.Y(n_2903)
);

NAND2x1p5_ASAP7_75t_L g2904 ( 
.A(n_2430),
.B(n_2433),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2238),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2257),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_SL g2907 ( 
.A(n_2400),
.B(n_1516),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_SL g2908 ( 
.A(n_2282),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2316),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2515),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2513),
.Y(n_2911)
);

INVxp67_ASAP7_75t_L g2912 ( 
.A(n_2546),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2408),
.B(n_1417),
.Y(n_2913)
);

AO22x2_ASAP7_75t_L g2914 ( 
.A1(n_2442),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_2914)
);

INVx3_ASAP7_75t_L g2915 ( 
.A(n_2476),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2580),
.B(n_1418),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2525),
.Y(n_2917)
);

NAND3xp33_ASAP7_75t_L g2918 ( 
.A(n_2553),
.B(n_1300),
.C(n_1220),
.Y(n_2918)
);

BUFx10_ASAP7_75t_L g2919 ( 
.A(n_2290),
.Y(n_2919)
);

AO22x2_ASAP7_75t_L g2920 ( 
.A1(n_2229),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_2920)
);

INVx5_ASAP7_75t_L g2921 ( 
.A(n_2373),
.Y(n_2921)
);

OAI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2405),
.A2(n_2443),
.B1(n_2458),
.B2(n_2435),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2527),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2469),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2495),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2322),
.B(n_1423),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2485),
.B(n_6),
.Y(n_2927)
);

INVxp67_ASAP7_75t_L g2928 ( 
.A(n_2468),
.Y(n_2928)
);

BUFx8_ASAP7_75t_L g2929 ( 
.A(n_2286),
.Y(n_2929)
);

INVx1_ASAP7_75t_SL g2930 ( 
.A(n_2579),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2474),
.Y(n_2931)
);

AO22x2_ASAP7_75t_L g2932 ( 
.A1(n_2454),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_2932)
);

AND2x2_ASAP7_75t_SL g2933 ( 
.A(n_2489),
.B(n_1470),
.Y(n_2933)
);

AOI22x1_ASAP7_75t_L g2934 ( 
.A1(n_2484),
.A2(n_2490),
.B1(n_2498),
.B2(n_2494),
.Y(n_2934)
);

INVxp67_ASAP7_75t_L g2935 ( 
.A(n_2478),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2477),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2411),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2526),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_SL g2939 ( 
.A1(n_2383),
.A2(n_1476),
.B1(n_1479),
.B2(n_1473),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2526),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2503),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2414),
.Y(n_2942)
);

AO22x2_ASAP7_75t_L g2943 ( 
.A1(n_2488),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2418),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2431),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2563),
.B(n_1424),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2423),
.B(n_1426),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2496),
.Y(n_2948)
);

NAND2x1p5_ASAP7_75t_L g2949 ( 
.A(n_2589),
.B(n_2403),
.Y(n_2949)
);

INVxp67_ASAP7_75t_L g2950 ( 
.A(n_2487),
.Y(n_2950)
);

HB1xp67_ASAP7_75t_L g2951 ( 
.A(n_2486),
.Y(n_2951)
);

AOI22x1_ASAP7_75t_L g2952 ( 
.A1(n_2517),
.A2(n_1300),
.B1(n_1321),
.B2(n_1220),
.Y(n_2952)
);

INVxp67_ASAP7_75t_L g2953 ( 
.A(n_2475),
.Y(n_2953)
);

NOR2xp33_ASAP7_75t_R g2954 ( 
.A(n_2335),
.B(n_1432),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2496),
.Y(n_2955)
);

CKINVDCx5p33_ASAP7_75t_R g2956 ( 
.A(n_2345),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2462),
.B(n_1510),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2480),
.Y(n_2958)
);

BUFx6f_ASAP7_75t_L g2959 ( 
.A(n_2347),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2403),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2483),
.B(n_2264),
.Y(n_2961)
);

NAND2x1p5_ASAP7_75t_L g2962 ( 
.A(n_2410),
.B(n_1321),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2410),
.Y(n_2963)
);

CKINVDCx5p33_ASAP7_75t_R g2964 ( 
.A(n_2365),
.Y(n_2964)
);

AND2x6_ASAP7_75t_L g2965 ( 
.A(n_2518),
.B(n_1321),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2492),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2497),
.Y(n_2967)
);

AND2x2_ASAP7_75t_SL g2968 ( 
.A(n_2524),
.B(n_1545),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2519),
.Y(n_2969)
);

INVx3_ASAP7_75t_L g2970 ( 
.A(n_2399),
.Y(n_2970)
);

INVxp67_ASAP7_75t_L g2971 ( 
.A(n_2417),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2523),
.B(n_1434),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2368),
.B(n_1435),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2499),
.Y(n_2974)
);

AOI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_2509),
.A2(n_1440),
.B1(n_1442),
.B2(n_1439),
.Y(n_2975)
);

NAND2x1p5_ASAP7_75t_L g2976 ( 
.A(n_2501),
.B(n_1356),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2538),
.B(n_1445),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2507),
.Y(n_2978)
);

INVx2_ASAP7_75t_SL g2979 ( 
.A(n_2521),
.Y(n_2979)
);

NOR2xp33_ASAP7_75t_L g2980 ( 
.A(n_2574),
.B(n_1446),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2583),
.B(n_1447),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2344),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2372),
.Y(n_2983)
);

A2O1A1Ixp33_ASAP7_75t_L g2984 ( 
.A1(n_2502),
.A2(n_1410),
.B(n_1468),
.C(n_1356),
.Y(n_2984)
);

NAND3xp33_ASAP7_75t_L g2985 ( 
.A(n_2417),
.B(n_1410),
.C(n_1356),
.Y(n_2985)
);

INVxp67_ASAP7_75t_L g2986 ( 
.A(n_2504),
.Y(n_2986)
);

AND2x4_ASAP7_75t_L g2987 ( 
.A(n_2380),
.B(n_9),
.Y(n_2987)
);

AND2x6_ASAP7_75t_L g2988 ( 
.A(n_2289),
.B(n_1356),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2226),
.Y(n_2989)
);

A2O1A1Ixp33_ASAP7_75t_L g2990 ( 
.A1(n_2244),
.A2(n_1468),
.B(n_1470),
.C(n_1410),
.Y(n_2990)
);

INVxp67_ASAP7_75t_L g2991 ( 
.A(n_2591),
.Y(n_2991)
);

AND2x4_ASAP7_75t_L g2992 ( 
.A(n_2289),
.B(n_10),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2522),
.A2(n_1448),
.B1(n_1455),
.B2(n_1453),
.Y(n_2993)
);

AO22x2_ASAP7_75t_L g2994 ( 
.A1(n_2367),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2226),
.Y(n_2995)
);

AO22x2_ASAP7_75t_L g2996 ( 
.A1(n_2367),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2413),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2413),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2247),
.B(n_1456),
.Y(n_2999)
);

NOR3xp33_ASAP7_75t_L g3000 ( 
.A(n_2222),
.B(n_1460),
.C(n_1457),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2299),
.A2(n_1461),
.B1(n_1464),
.B2(n_1462),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2247),
.B(n_1480),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2228),
.B(n_1485),
.Y(n_3003)
);

INVxp67_ASAP7_75t_L g3004 ( 
.A(n_2591),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2223),
.B(n_1542),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2247),
.B(n_1487),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2289),
.B(n_12),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2226),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2226),
.Y(n_3009)
);

AND2x4_ASAP7_75t_L g3010 ( 
.A(n_2289),
.B(n_13),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_2591),
.B(n_1494),
.Y(n_3011)
);

OR2x2_ASAP7_75t_SL g3012 ( 
.A(n_2310),
.B(n_1410),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2226),
.Y(n_3013)
);

BUFx2_ASAP7_75t_L g3014 ( 
.A(n_2255),
.Y(n_3014)
);

AO22x2_ASAP7_75t_L g3015 ( 
.A1(n_2367),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2413),
.Y(n_3016)
);

BUFx6f_ASAP7_75t_L g3017 ( 
.A(n_2543),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2413),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2226),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2247),
.B(n_1495),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2226),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2226),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2226),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2226),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2228),
.A2(n_1470),
.B1(n_1468),
.B2(n_18),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2226),
.Y(n_3026)
);

NAND2xp33_ASAP7_75t_L g3027 ( 
.A(n_2255),
.B(n_1468),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2413),
.Y(n_3028)
);

AO22x2_ASAP7_75t_L g3029 ( 
.A1(n_2367),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_3029)
);

NAND2x1p5_ASAP7_75t_L g3030 ( 
.A(n_2223),
.B(n_1470),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2413),
.Y(n_3031)
);

CKINVDCx16_ASAP7_75t_R g3032 ( 
.A(n_2572),
.Y(n_3032)
);

OAI221xp5_ASAP7_75t_L g3033 ( 
.A1(n_2301),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.C(n_21),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2591),
.B(n_19),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2226),
.Y(n_3035)
);

AO22x2_ASAP7_75t_L g3036 ( 
.A1(n_2367),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2413),
.Y(n_3037)
);

NAND2x1p5_ASAP7_75t_L g3038 ( 
.A(n_2223),
.B(n_23),
.Y(n_3038)
);

OR2x2_ASAP7_75t_L g3039 ( 
.A(n_2277),
.B(n_23),
.Y(n_3039)
);

OAI221xp5_ASAP7_75t_L g3040 ( 
.A1(n_2301),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.C(n_27),
.Y(n_3040)
);

HB1xp67_ASAP7_75t_L g3041 ( 
.A(n_2223),
.Y(n_3041)
);

OR2x2_ASAP7_75t_SL g3042 ( 
.A(n_2310),
.B(n_24),
.Y(n_3042)
);

OAI22xp5_ASAP7_75t_L g3043 ( 
.A1(n_2299),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_3043)
);

BUFx3_ASAP7_75t_L g3044 ( 
.A(n_2223),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2226),
.Y(n_3045)
);

INVx3_ASAP7_75t_L g3046 ( 
.A(n_2223),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2413),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2413),
.Y(n_3048)
);

AOI22xp33_ASAP7_75t_L g3049 ( 
.A1(n_2522),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_3049)
);

NAND2x1p5_ASAP7_75t_L g3050 ( 
.A(n_2223),
.B(n_27),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2413),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2591),
.B(n_28),
.Y(n_3052)
);

AOI22xp5_ASAP7_75t_L g3053 ( 
.A1(n_2228),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2413),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2226),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2226),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2226),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2228),
.B(n_29),
.Y(n_3058)
);

HB1xp67_ASAP7_75t_L g3059 ( 
.A(n_2223),
.Y(n_3059)
);

OR2x2_ASAP7_75t_SL g3060 ( 
.A(n_2310),
.B(n_29),
.Y(n_3060)
);

OR2x2_ASAP7_75t_L g3061 ( 
.A(n_2277),
.B(n_30),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2413),
.Y(n_3062)
);

INVx1_ASAP7_75t_SL g3063 ( 
.A(n_2277),
.Y(n_3063)
);

AO22x2_ASAP7_75t_L g3064 ( 
.A1(n_2367),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_3064)
);

HB1xp67_ASAP7_75t_L g3065 ( 
.A(n_2223),
.Y(n_3065)
);

BUFx6f_ASAP7_75t_L g3066 ( 
.A(n_2543),
.Y(n_3066)
);

A2O1A1Ixp33_ASAP7_75t_L g3067 ( 
.A1(n_2244),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_3067)
);

AOI22xp5_ASAP7_75t_L g3068 ( 
.A1(n_2228),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2226),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2413),
.Y(n_3070)
);

AND2x4_ASAP7_75t_L g3071 ( 
.A(n_2289),
.B(n_33),
.Y(n_3071)
);

NOR2xp67_ASAP7_75t_L g3072 ( 
.A(n_2223),
.B(n_34),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2247),
.B(n_34),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2223),
.B(n_35),
.Y(n_3074)
);

AO22x2_ASAP7_75t_L g3075 ( 
.A1(n_2367),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2223),
.B(n_36),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_2228),
.B(n_35),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_SL g3078 ( 
.A(n_2223),
.B(n_39),
.Y(n_3078)
);

AO22x2_ASAP7_75t_L g3079 ( 
.A1(n_2367),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_3079)
);

BUFx8_ASAP7_75t_L g3080 ( 
.A(n_2425),
.Y(n_3080)
);

BUFx3_ASAP7_75t_L g3081 ( 
.A(n_2223),
.Y(n_3081)
);

BUFx12f_ASAP7_75t_L g3082 ( 
.A(n_2481),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2226),
.Y(n_3083)
);

AOI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_2228),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_3084)
);

NAND2xp33_ASAP7_75t_L g3085 ( 
.A(n_2255),
.B(n_41),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2226),
.Y(n_3086)
);

HB1xp67_ASAP7_75t_L g3087 ( 
.A(n_2223),
.Y(n_3087)
);

CKINVDCx5p33_ASAP7_75t_R g3088 ( 
.A(n_2481),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2226),
.Y(n_3089)
);

INVxp67_ASAP7_75t_L g3090 ( 
.A(n_2591),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_L g3091 ( 
.A(n_2228),
.B(n_40),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2247),
.B(n_41),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2413),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2247),
.B(n_42),
.Y(n_3094)
);

INVxp67_ASAP7_75t_L g3095 ( 
.A(n_2591),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2226),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2413),
.Y(n_3097)
);

NAND2x1p5_ASAP7_75t_L g3098 ( 
.A(n_2223),
.B(n_42),
.Y(n_3098)
);

BUFx2_ASAP7_75t_L g3099 ( 
.A(n_2255),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2226),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2226),
.Y(n_3101)
);

HB1xp67_ASAP7_75t_L g3102 ( 
.A(n_2223),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2413),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2226),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2591),
.B(n_43),
.Y(n_3105)
);

AND2x2_ASAP7_75t_SL g3106 ( 
.A(n_2317),
.B(n_43),
.Y(n_3106)
);

NAND2x1p5_ASAP7_75t_L g3107 ( 
.A(n_2223),
.B(n_43),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2226),
.Y(n_3108)
);

OR2x6_ASAP7_75t_L g3109 ( 
.A(n_2363),
.B(n_44),
.Y(n_3109)
);

AND2x4_ASAP7_75t_L g3110 ( 
.A(n_2289),
.B(n_44),
.Y(n_3110)
);

NAND2xp33_ASAP7_75t_L g3111 ( 
.A(n_2255),
.B(n_46),
.Y(n_3111)
);

NOR2xp33_ASAP7_75t_L g3112 ( 
.A(n_2228),
.B(n_45),
.Y(n_3112)
);

AO22x2_ASAP7_75t_L g3113 ( 
.A1(n_2367),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_2522),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2413),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2226),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2226),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2247),
.B(n_48),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2413),
.Y(n_3119)
);

AOI22xp33_ASAP7_75t_L g3120 ( 
.A1(n_2522),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2226),
.Y(n_3121)
);

AOI22xp33_ASAP7_75t_L g3122 ( 
.A1(n_2522),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2591),
.B(n_49),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2226),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2247),
.B(n_51),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2226),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2247),
.B(n_52),
.Y(n_3127)
);

AND2x4_ASAP7_75t_L g3128 ( 
.A(n_2289),
.B(n_52),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2226),
.Y(n_3129)
);

INVx2_ASAP7_75t_L g3130 ( 
.A(n_2413),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2226),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2226),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2226),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2413),
.Y(n_3134)
);

A2O1A1Ixp33_ASAP7_75t_L g3135 ( 
.A1(n_2244),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2413),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2247),
.B(n_53),
.Y(n_3137)
);

AND2x4_ASAP7_75t_L g3138 ( 
.A(n_2289),
.B(n_54),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2413),
.Y(n_3139)
);

NAND2x1p5_ASAP7_75t_L g3140 ( 
.A(n_2223),
.B(n_54),
.Y(n_3140)
);

AO22x2_ASAP7_75t_L g3141 ( 
.A1(n_2367),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2413),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2413),
.Y(n_3143)
);

CKINVDCx5p33_ASAP7_75t_R g3144 ( 
.A(n_2481),
.Y(n_3144)
);

AO22x2_ASAP7_75t_L g3145 ( 
.A1(n_2367),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_3145)
);

O2A1O1Ixp33_ASAP7_75t_L g3146 ( 
.A1(n_2301),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2413),
.Y(n_3147)
);

INVxp33_ASAP7_75t_L g3148 ( 
.A(n_2284),
.Y(n_3148)
);

AOI22xp33_ASAP7_75t_L g3149 ( 
.A1(n_2522),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_3149)
);

HB1xp67_ASAP7_75t_L g3150 ( 
.A(n_2223),
.Y(n_3150)
);

INVxp67_ASAP7_75t_L g3151 ( 
.A(n_2591),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2228),
.B(n_58),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2226),
.Y(n_3153)
);

INVx4_ASAP7_75t_L g3154 ( 
.A(n_2223),
.Y(n_3154)
);

NAND2x1p5_ASAP7_75t_L g3155 ( 
.A(n_2223),
.B(n_58),
.Y(n_3155)
);

HB1xp67_ASAP7_75t_L g3156 ( 
.A(n_2223),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2591),
.B(n_59),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2226),
.Y(n_3158)
);

AO22x2_ASAP7_75t_L g3159 ( 
.A1(n_2367),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_3159)
);

INVx2_ASAP7_75t_SL g3160 ( 
.A(n_2223),
.Y(n_3160)
);

INVx8_ASAP7_75t_L g3161 ( 
.A(n_2363),
.Y(n_3161)
);

AND2x4_ASAP7_75t_L g3162 ( 
.A(n_2289),
.B(n_60),
.Y(n_3162)
);

NOR2xp67_ASAP7_75t_L g3163 ( 
.A(n_2223),
.B(n_61),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2226),
.Y(n_3164)
);

AO22x2_ASAP7_75t_L g3165 ( 
.A1(n_2367),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2413),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2226),
.Y(n_3167)
);

INVxp67_ASAP7_75t_L g3168 ( 
.A(n_2591),
.Y(n_3168)
);

BUFx3_ASAP7_75t_L g3169 ( 
.A(n_2223),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2226),
.Y(n_3170)
);

AOI22xp5_ASAP7_75t_L g3171 ( 
.A1(n_2228),
.A2(n_65),
.B1(n_62),
.B2(n_63),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2413),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_SL g3173 ( 
.A(n_2223),
.B(n_66),
.Y(n_3173)
);

NAND2xp33_ASAP7_75t_L g3174 ( 
.A(n_2255),
.B(n_66),
.Y(n_3174)
);

INVxp67_ASAP7_75t_SL g3175 ( 
.A(n_2549),
.Y(n_3175)
);

AOI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_2228),
.A2(n_68),
.B1(n_65),
.B2(n_66),
.Y(n_3176)
);

OR2x2_ASAP7_75t_SL g3177 ( 
.A(n_2310),
.B(n_68),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2413),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2226),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2226),
.Y(n_3180)
);

AND2x2_ASAP7_75t_L g3181 ( 
.A(n_2591),
.B(n_68),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2247),
.B(n_69),
.Y(n_3182)
);

BUFx4f_ASAP7_75t_L g3183 ( 
.A(n_2363),
.Y(n_3183)
);

INVx3_ASAP7_75t_L g3184 ( 
.A(n_2223),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2247),
.B(n_69),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2413),
.Y(n_3186)
);

AND2x4_ASAP7_75t_L g3187 ( 
.A(n_2289),
.B(n_69),
.Y(n_3187)
);

HB1xp67_ASAP7_75t_L g3188 ( 
.A(n_2223),
.Y(n_3188)
);

INVxp33_ASAP7_75t_L g3189 ( 
.A(n_2284),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2413),
.Y(n_3190)
);

INVxp67_ASAP7_75t_L g3191 ( 
.A(n_2591),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2413),
.Y(n_3192)
);

CKINVDCx5p33_ASAP7_75t_R g3193 ( 
.A(n_2481),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2413),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2413),
.Y(n_3195)
);

AOI22xp5_ASAP7_75t_SL g3196 ( 
.A1(n_2572),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3196)
);

NAND2x1p5_ASAP7_75t_L g3197 ( 
.A(n_2223),
.B(n_70),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2413),
.Y(n_3198)
);

NOR2xp33_ASAP7_75t_L g3199 ( 
.A(n_2228),
.B(n_70),
.Y(n_3199)
);

AO22x2_ASAP7_75t_L g3200 ( 
.A1(n_2367),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2413),
.Y(n_3201)
);

INVxp67_ASAP7_75t_L g3202 ( 
.A(n_2591),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_2481),
.Y(n_3203)
);

AND2x4_ASAP7_75t_L g3204 ( 
.A(n_2289),
.B(n_71),
.Y(n_3204)
);

AND2x2_ASAP7_75t_L g3205 ( 
.A(n_2591),
.B(n_72),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2226),
.Y(n_3206)
);

AND2x4_ASAP7_75t_L g3207 ( 
.A(n_2289),
.B(n_73),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2247),
.B(n_74),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2413),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_2228),
.B(n_74),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2247),
.B(n_75),
.Y(n_3211)
);

AND2x4_ASAP7_75t_L g3212 ( 
.A(n_2289),
.B(n_75),
.Y(n_3212)
);

CKINVDCx5p33_ASAP7_75t_R g3213 ( 
.A(n_2481),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2226),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2226),
.Y(n_3215)
);

AO22x2_ASAP7_75t_L g3216 ( 
.A1(n_2367),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_3216)
);

AND2x4_ASAP7_75t_L g3217 ( 
.A(n_2289),
.B(n_76),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2413),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2226),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2247),
.B(n_76),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2226),
.Y(n_3221)
);

INVxp67_ASAP7_75t_L g3222 ( 
.A(n_2591),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_2226),
.Y(n_3223)
);

AND2x4_ASAP7_75t_L g3224 ( 
.A(n_2289),
.B(n_77),
.Y(n_3224)
);

AO22x2_ASAP7_75t_L g3225 ( 
.A1(n_2367),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_3225)
);

AO22x2_ASAP7_75t_L g3226 ( 
.A1(n_2367),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_2413),
.Y(n_3227)
);

NAND2x1p5_ASAP7_75t_L g3228 ( 
.A(n_2223),
.B(n_78),
.Y(n_3228)
);

INVxp67_ASAP7_75t_L g3229 ( 
.A(n_2591),
.Y(n_3229)
);

OAI22xp33_ASAP7_75t_L g3230 ( 
.A1(n_2228),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3230)
);

OAI22xp5_ASAP7_75t_L g3231 ( 
.A1(n_2299),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_3231)
);

AND2x4_ASAP7_75t_L g3232 ( 
.A(n_2289),
.B(n_81),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2226),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2413),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2226),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2226),
.Y(n_3236)
);

AND2x4_ASAP7_75t_L g3237 ( 
.A(n_2289),
.B(n_82),
.Y(n_3237)
);

AOI21x1_ASAP7_75t_L g3238 ( 
.A1(n_2863),
.A2(n_3014),
.B(n_2701),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2697),
.Y(n_3239)
);

AOI21xp5_ASAP7_75t_L g3240 ( 
.A1(n_2842),
.A2(n_83),
.B(n_84),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_2865),
.B(n_83),
.Y(n_3241)
);

INVxp33_ASAP7_75t_SL g3242 ( 
.A(n_2832),
.Y(n_3242)
);

AOI22xp5_ASAP7_75t_L g3243 ( 
.A1(n_3106),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_3243)
);

INVxp67_ASAP7_75t_L g3244 ( 
.A(n_3175),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_3027),
.A2(n_85),
.B(n_86),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_2650),
.Y(n_3246)
);

AOI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_2922),
.A2(n_86),
.B(n_87),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3073),
.A2(n_87),
.B(n_88),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_2968),
.B(n_2696),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2772),
.B(n_87),
.Y(n_3250)
);

AOI21x1_ASAP7_75t_L g3251 ( 
.A1(n_2701),
.A2(n_88),
.B(n_89),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2653),
.Y(n_3252)
);

OR2x2_ASAP7_75t_L g3253 ( 
.A(n_2640),
.B(n_89),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2655),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2782),
.B(n_89),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_SL g3256 ( 
.A(n_2886),
.B(n_2933),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_3092),
.A2(n_3118),
.B(n_3094),
.Y(n_3257)
);

AND2x4_ASAP7_75t_L g3258 ( 
.A(n_2921),
.B(n_90),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_SL g3259 ( 
.A(n_3014),
.B(n_120),
.Y(n_3259)
);

CKINVDCx10_ASAP7_75t_R g3260 ( 
.A(n_2823),
.Y(n_3260)
);

AOI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_2750),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_3261)
);

AOI22x1_ASAP7_75t_L g3262 ( 
.A1(n_2860),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_2784),
.B(n_91),
.Y(n_3263)
);

OAI22xp5_ASAP7_75t_L g3264 ( 
.A1(n_3099),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_3264)
);

OAI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_2610),
.A2(n_94),
.B(n_95),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_3125),
.A2(n_3137),
.B(n_3127),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2786),
.B(n_94),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_2868),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_3182),
.A2(n_96),
.B(n_97),
.Y(n_3269)
);

AOI21xp33_ASAP7_75t_L g3270 ( 
.A1(n_3185),
.A2(n_98),
.B(n_99),
.Y(n_3270)
);

AOI21x1_ASAP7_75t_L g3271 ( 
.A1(n_3099),
.A2(n_98),
.B(n_99),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3208),
.A2(n_98),
.B(n_99),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3211),
.A2(n_100),
.B(n_101),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_2601),
.B(n_100),
.Y(n_3274)
);

O2A1O1Ixp33_ASAP7_75t_L g3275 ( 
.A1(n_3230),
.A2(n_2620),
.B(n_3220),
.C(n_3135),
.Y(n_3275)
);

AOI21xp5_ASAP7_75t_L g3276 ( 
.A1(n_3085),
.A2(n_101),
.B(n_102),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3011),
.B(n_101),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_3111),
.A2(n_102),
.B(n_103),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2602),
.B(n_102),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_3174),
.A2(n_2888),
.B(n_2670),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_2664),
.A2(n_103),
.B(n_104),
.Y(n_3281)
);

OAI21x1_ASAP7_75t_L g3282 ( 
.A1(n_2934),
.A2(n_103),
.B(n_104),
.Y(n_3282)
);

AOI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_2692),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_2693),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_2674),
.A2(n_105),
.B(n_106),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2607),
.B(n_106),
.Y(n_3286)
);

AOI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_2680),
.A2(n_107),
.B(n_108),
.Y(n_3287)
);

AOI21x1_ASAP7_75t_L g3288 ( 
.A1(n_2866),
.A2(n_107),
.B(n_108),
.Y(n_3288)
);

AOI22x1_ASAP7_75t_L g3289 ( 
.A1(n_2600),
.A2(n_3030),
.B1(n_2976),
.B2(n_2814),
.Y(n_3289)
);

AOI21xp5_ASAP7_75t_L g3290 ( 
.A1(n_2681),
.A2(n_107),
.B(n_108),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2613),
.B(n_109),
.Y(n_3291)
);

A2O1A1Ixp33_ASAP7_75t_L g3292 ( 
.A1(n_3146),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2614),
.B(n_109),
.Y(n_3293)
);

OAI22xp5_ASAP7_75t_L g3294 ( 
.A1(n_2678),
.A2(n_113),
.B1(n_110),
.B2(n_112),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_2785),
.A2(n_113),
.B(n_114),
.Y(n_3295)
);

AOI22x1_ASAP7_75t_SL g3296 ( 
.A1(n_2605),
.A2(n_3088),
.B1(n_3193),
.B2(n_3144),
.Y(n_3296)
);

A2O1A1Ixp33_ASAP7_75t_L g3297 ( 
.A1(n_2749),
.A2(n_116),
.B(n_113),
.C(n_115),
.Y(n_3297)
);

AOI21xp5_ASAP7_75t_L g3298 ( 
.A1(n_2898),
.A2(n_115),
.B(n_116),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_SL g3299 ( 
.A(n_2971),
.B(n_120),
.Y(n_3299)
);

INVx3_ASAP7_75t_L g3300 ( 
.A(n_2626),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_2690),
.A2(n_115),
.B(n_116),
.Y(n_3301)
);

OAI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2755),
.A2(n_117),
.B(n_118),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_L g3303 ( 
.A(n_2760),
.B(n_117),
.Y(n_3303)
);

NAND2x1_ASAP7_75t_L g3304 ( 
.A(n_2988),
.B(n_2626),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_2767),
.A2(n_117),
.B(n_118),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_2597),
.Y(n_3306)
);

BUFx6f_ASAP7_75t_L g3307 ( 
.A(n_2768),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_2854),
.B(n_2953),
.Y(n_3308)
);

OR2x2_ASAP7_75t_L g3309 ( 
.A(n_3032),
.B(n_118),
.Y(n_3309)
);

OR2x6_ASAP7_75t_L g3310 ( 
.A(n_3161),
.B(n_119),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_2615),
.Y(n_3311)
);

OAI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2641),
.A2(n_119),
.B(n_121),
.Y(n_3312)
);

INVx3_ASAP7_75t_L g3313 ( 
.A(n_3017),
.Y(n_3313)
);

AOI21x1_ASAP7_75t_L g3314 ( 
.A1(n_2867),
.A2(n_119),
.B(n_123),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_2997),
.Y(n_3315)
);

BUFx8_ASAP7_75t_L g3316 ( 
.A(n_3082),
.Y(n_3316)
);

AOI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_3234),
.A2(n_124),
.B(n_125),
.Y(n_3317)
);

A2O1A1Ixp33_ASAP7_75t_L g3318 ( 
.A1(n_3067),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_2998),
.A2(n_3018),
.B(n_3016),
.Y(n_3319)
);

AOI21xp5_ASAP7_75t_L g3320 ( 
.A1(n_3028),
.A2(n_126),
.B(n_127),
.Y(n_3320)
);

OAI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_2811),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_3321)
);

AOI21xp5_ASAP7_75t_L g3322 ( 
.A1(n_3031),
.A2(n_128),
.B(n_129),
.Y(n_3322)
);

BUFx3_ASAP7_75t_L g3323 ( 
.A(n_3161),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2625),
.B(n_130),
.Y(n_3324)
);

AO21x2_ASAP7_75t_L g3325 ( 
.A1(n_2990),
.A2(n_132),
.B(n_133),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_3227),
.A2(n_132),
.B(n_134),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3037),
.A2(n_134),
.B(n_135),
.Y(n_3327)
);

CKINVDCx10_ASAP7_75t_R g3328 ( 
.A(n_2908),
.Y(n_3328)
);

AOI21xp5_ASAP7_75t_L g3329 ( 
.A1(n_3047),
.A2(n_135),
.B(n_136),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_3148),
.B(n_136),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_3048),
.A2(n_3054),
.B(n_3051),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2628),
.B(n_137),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2629),
.B(n_137),
.Y(n_3333)
);

NOR2xp33_ASAP7_75t_L g3334 ( 
.A(n_2928),
.B(n_138),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2630),
.B(n_139),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3062),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_2633),
.Y(n_3337)
);

BUFx6f_ASAP7_75t_L g3338 ( 
.A(n_2768),
.Y(n_3338)
);

AOI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_3070),
.A2(n_140),
.B(n_141),
.Y(n_3339)
);

AOI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_3093),
.A2(n_3103),
.B(n_3097),
.Y(n_3340)
);

OAI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_2999),
.A2(n_3006),
.B(n_3002),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2634),
.B(n_140),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3115),
.A2(n_141),
.B(n_142),
.Y(n_3343)
);

OAI21xp5_ASAP7_75t_L g3344 ( 
.A1(n_3020),
.A2(n_142),
.B(n_143),
.Y(n_3344)
);

AOI21xp5_ASAP7_75t_L g3345 ( 
.A1(n_3119),
.A2(n_143),
.B(n_144),
.Y(n_3345)
);

INVx11_ASAP7_75t_L g3346 ( 
.A(n_2644),
.Y(n_3346)
);

NOR2xp33_ASAP7_75t_L g3347 ( 
.A(n_2935),
.B(n_145),
.Y(n_3347)
);

OAI22xp5_ASAP7_75t_L g3348 ( 
.A1(n_2811),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_3348)
);

AOI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_3130),
.A2(n_3136),
.B(n_3134),
.Y(n_3349)
);

AOI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_3139),
.A2(n_146),
.B(n_148),
.Y(n_3350)
);

AOI21xp5_ASAP7_75t_L g3351 ( 
.A1(n_3142),
.A2(n_149),
.B(n_151),
.Y(n_3351)
);

BUFx6f_ASAP7_75t_L g3352 ( 
.A(n_2768),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3143),
.A2(n_149),
.B(n_152),
.Y(n_3353)
);

BUFx3_ASAP7_75t_L g3354 ( 
.A(n_3183),
.Y(n_3354)
);

AOI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_3147),
.A2(n_152),
.B(n_153),
.Y(n_3355)
);

OAI321xp33_ASAP7_75t_L g3356 ( 
.A1(n_3033),
.A2(n_3040),
.A3(n_3109),
.B1(n_3231),
.B2(n_3043),
.C(n_3025),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_2598),
.B(n_154),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_2635),
.B(n_155),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_2991),
.B(n_155),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_L g3360 ( 
.A(n_2950),
.B(n_156),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2637),
.B(n_157),
.Y(n_3361)
);

BUFx6f_ASAP7_75t_L g3362 ( 
.A(n_3017),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3004),
.B(n_158),
.Y(n_3363)
);

NOR2xp33_ASAP7_75t_L g3364 ( 
.A(n_2735),
.B(n_159),
.Y(n_3364)
);

OAI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_2874),
.A2(n_163),
.B1(n_159),
.B2(n_160),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_SL g3366 ( 
.A(n_3189),
.B(n_163),
.Y(n_3366)
);

INVxp67_ASAP7_75t_L g3367 ( 
.A(n_2732),
.Y(n_3367)
);

AOI22xp5_ASAP7_75t_L g3368 ( 
.A1(n_2939),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_3368)
);

AOI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_3166),
.A2(n_165),
.B(n_166),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_2638),
.B(n_167),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_2812),
.B(n_168),
.Y(n_3371)
);

OAI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_2744),
.A2(n_169),
.B(n_170),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_2639),
.B(n_170),
.Y(n_3373)
);

OAI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_2777),
.A2(n_171),
.B(n_172),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_3172),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_3178),
.Y(n_3376)
);

AOI33xp33_ASAP7_75t_L g3377 ( 
.A1(n_2754),
.A2(n_175),
.A3(n_177),
.B1(n_173),
.B2(n_174),
.B3(n_176),
.Y(n_3377)
);

AOI21xp5_ASAP7_75t_L g3378 ( 
.A1(n_3186),
.A2(n_173),
.B(n_175),
.Y(n_3378)
);

OR2x6_ASAP7_75t_L g3379 ( 
.A(n_3109),
.B(n_176),
.Y(n_3379)
);

AOI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_3190),
.A2(n_177),
.B(n_178),
.Y(n_3380)
);

NOR2xp33_ASAP7_75t_L g3381 ( 
.A(n_2833),
.B(n_178),
.Y(n_3381)
);

NAND3xp33_ASAP7_75t_L g3382 ( 
.A(n_2984),
.B(n_179),
.C(n_180),
.Y(n_3382)
);

NOR3xp33_ASAP7_75t_L g3383 ( 
.A(n_2852),
.B(n_179),
.C(n_180),
.Y(n_3383)
);

INVx3_ASAP7_75t_L g3384 ( 
.A(n_3066),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_2642),
.B(n_181),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_3090),
.B(n_181),
.Y(n_3386)
);

NOR2x1_ASAP7_75t_L g3387 ( 
.A(n_2728),
.B(n_182),
.Y(n_3387)
);

A2O1A1Ixp33_ASAP7_75t_L g3388 ( 
.A1(n_2847),
.A2(n_186),
.B(n_183),
.C(n_185),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_2649),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_3192),
.Y(n_3390)
);

O2A1O1Ixp5_ASAP7_75t_L g3391 ( 
.A1(n_2869),
.A2(n_186),
.B(n_183),
.C(n_185),
.Y(n_3391)
);

INVx4_ASAP7_75t_L g3392 ( 
.A(n_2921),
.Y(n_3392)
);

AND2x2_ASAP7_75t_L g3393 ( 
.A(n_3095),
.B(n_187),
.Y(n_3393)
);

OAI21x1_ASAP7_75t_L g3394 ( 
.A1(n_2745),
.A2(n_188),
.B(n_189),
.Y(n_3394)
);

AOI21xp5_ASAP7_75t_L g3395 ( 
.A1(n_3194),
.A2(n_188),
.B(n_189),
.Y(n_3395)
);

CKINVDCx8_ASAP7_75t_R g3396 ( 
.A(n_3203),
.Y(n_3396)
);

OAI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_2788),
.A2(n_190),
.B(n_191),
.Y(n_3397)
);

A2O1A1Ixp33_ASAP7_75t_L g3398 ( 
.A1(n_2717),
.A2(n_192),
.B(n_190),
.C(n_191),
.Y(n_3398)
);

O2A1O1Ixp33_ASAP7_75t_L g3399 ( 
.A1(n_2710),
.A2(n_195),
.B(n_192),
.C(n_193),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3195),
.A2(n_193),
.B(n_195),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_3198),
.Y(n_3401)
);

OAI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_2794),
.A2(n_196),
.B(n_197),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3201),
.A2(n_196),
.B(n_197),
.Y(n_3403)
);

AOI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_3209),
.A2(n_198),
.B(n_199),
.Y(n_3404)
);

AOI21xp5_ASAP7_75t_L g3405 ( 
.A1(n_3218),
.A2(n_199),
.B(n_200),
.Y(n_3405)
);

NAND2x1p5_ASAP7_75t_L g3406 ( 
.A(n_2627),
.B(n_200),
.Y(n_3406)
);

AOI21xp5_ASAP7_75t_L g3407 ( 
.A1(n_2604),
.A2(n_201),
.B(n_202),
.Y(n_3407)
);

AO21x1_ASAP7_75t_L g3408 ( 
.A1(n_2874),
.A2(n_203),
.B(n_204),
.Y(n_3408)
);

INVx3_ASAP7_75t_L g3409 ( 
.A(n_3066),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_2623),
.A2(n_203),
.B(n_204),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_2654),
.B(n_205),
.Y(n_3411)
);

OAI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_2806),
.A2(n_206),
.B(n_207),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_2656),
.B(n_206),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_2624),
.A2(n_207),
.B(n_208),
.Y(n_3414)
);

AOI22xp33_ASAP7_75t_L g3415 ( 
.A1(n_2805),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_2658),
.B(n_210),
.Y(n_3416)
);

O2A1O1Ixp33_ASAP7_75t_SL g3417 ( 
.A1(n_2679),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_2659),
.B(n_2989),
.Y(n_3418)
);

AOI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_2645),
.A2(n_212),
.B(n_215),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_2699),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_SL g3421 ( 
.A(n_3151),
.B(n_215),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_2704),
.A2(n_216),
.B(n_217),
.Y(n_3422)
);

BUFx2_ASAP7_75t_L g3423 ( 
.A(n_2688),
.Y(n_3423)
);

INVx1_ASAP7_75t_SL g3424 ( 
.A(n_3063),
.Y(n_3424)
);

OAI21xp5_ASAP7_75t_L g3425 ( 
.A1(n_2838),
.A2(n_216),
.B(n_218),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_2995),
.B(n_218),
.Y(n_3426)
);

AND2x4_ASAP7_75t_L g3427 ( 
.A(n_2921),
.B(n_3044),
.Y(n_3427)
);

AOI21x1_ASAP7_75t_L g3428 ( 
.A1(n_2870),
.A2(n_219),
.B(n_220),
.Y(n_3428)
);

BUFx4f_ASAP7_75t_L g3429 ( 
.A(n_2883),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3008),
.Y(n_3430)
);

INVx3_ASAP7_75t_L g3431 ( 
.A(n_3154),
.Y(n_3431)
);

AOI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_2715),
.A2(n_219),
.B(n_221),
.Y(n_3432)
);

BUFx12f_ASAP7_75t_L g3433 ( 
.A(n_2644),
.Y(n_3433)
);

OAI21x1_ASAP7_75t_L g3434 ( 
.A1(n_2952),
.A2(n_221),
.B(n_222),
.Y(n_3434)
);

AOI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_2792),
.A2(n_222),
.B(n_223),
.Y(n_3435)
);

AOI21xp5_ASAP7_75t_L g3436 ( 
.A1(n_2793),
.A2(n_2817),
.B(n_2803),
.Y(n_3436)
);

BUFx6f_ASAP7_75t_L g3437 ( 
.A(n_2988),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_L g3438 ( 
.A(n_2897),
.B(n_223),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_2702),
.Y(n_3439)
);

BUFx6f_ASAP7_75t_L g3440 ( 
.A(n_2988),
.Y(n_3440)
);

AOI21xp5_ASAP7_75t_L g3441 ( 
.A1(n_2819),
.A2(n_2858),
.B(n_2849),
.Y(n_3441)
);

AO21x1_ASAP7_75t_L g3442 ( 
.A1(n_3074),
.A2(n_224),
.B(n_225),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3009),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_3168),
.B(n_3191),
.Y(n_3444)
);

AOI21xp5_ASAP7_75t_L g3445 ( 
.A1(n_2862),
.A2(n_2733),
.B(n_2711),
.Y(n_3445)
);

AOI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_2706),
.A2(n_224),
.B(n_225),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3013),
.B(n_226),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3019),
.Y(n_3448)
);

O2A1O1Ixp33_ASAP7_75t_SL g3449 ( 
.A1(n_3076),
.A2(n_3078),
.B(n_3173),
.C(n_2985),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3021),
.Y(n_3450)
);

INVx4_ASAP7_75t_L g3451 ( 
.A(n_3081),
.Y(n_3451)
);

HB1xp67_ASAP7_75t_L g3452 ( 
.A(n_3202),
.Y(n_3452)
);

BUFx2_ASAP7_75t_L g3453 ( 
.A(n_2683),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3022),
.B(n_226),
.Y(n_3454)
);

AOI21xp5_ASAP7_75t_L g3455 ( 
.A1(n_2712),
.A2(n_227),
.B(n_228),
.Y(n_3455)
);

O2A1O1Ixp33_ASAP7_75t_L g3456 ( 
.A1(n_3058),
.A2(n_231),
.B(n_228),
.C(n_230),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_3023),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3024),
.B(n_231),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3026),
.Y(n_3459)
);

OA22x2_ASAP7_75t_L g3460 ( 
.A1(n_2987),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3035),
.Y(n_3461)
);

AOI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_2721),
.A2(n_233),
.B(n_234),
.Y(n_3462)
);

OR2x6_ASAP7_75t_L g3463 ( 
.A(n_2883),
.B(n_235),
.Y(n_3463)
);

AOI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_2722),
.A2(n_235),
.B(n_236),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_2723),
.A2(n_237),
.B(n_238),
.Y(n_3465)
);

AOI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_2729),
.A2(n_237),
.B(n_239),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_2902),
.B(n_239),
.Y(n_3467)
);

OAI22xp5_ASAP7_75t_L g3468 ( 
.A1(n_2713),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_3468)
);

OAI22xp5_ASAP7_75t_L g3469 ( 
.A1(n_2713),
.A2(n_2660),
.B1(n_3229),
.B2(n_3222),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_2731),
.A2(n_2889),
.B(n_2882),
.Y(n_3470)
);

OAI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_2844),
.A2(n_240),
.B(n_242),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_2893),
.A2(n_245),
.B(n_246),
.Y(n_3472)
);

BUFx4f_ASAP7_75t_L g3473 ( 
.A(n_2661),
.Y(n_3473)
);

NOR2xp33_ASAP7_75t_L g3474 ( 
.A(n_2912),
.B(n_246),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_2734),
.B(n_247),
.Y(n_3475)
);

NOR2xp33_ASAP7_75t_L g3476 ( 
.A(n_3003),
.B(n_247),
.Y(n_3476)
);

AOI21x1_ASAP7_75t_L g3477 ( 
.A1(n_2871),
.A2(n_248),
.B(n_249),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3045),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3055),
.B(n_248),
.Y(n_3479)
);

OAI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_2853),
.A2(n_249),
.B(n_250),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3056),
.B(n_250),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_SL g3482 ( 
.A(n_2992),
.B(n_252),
.Y(n_3482)
);

BUFx4f_ASAP7_75t_L g3483 ( 
.A(n_2661),
.Y(n_3483)
);

OAI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_2875),
.A2(n_252),
.B(n_253),
.Y(n_3484)
);

AOI21xp5_ASAP7_75t_L g3485 ( 
.A1(n_2896),
.A2(n_253),
.B(n_254),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3057),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3069),
.B(n_254),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3083),
.Y(n_3488)
);

A2O1A1Ixp33_ASAP7_75t_L g3489 ( 
.A1(n_2816),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_3489)
);

A2O1A1Ixp33_ASAP7_75t_L g3490 ( 
.A1(n_3053),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3086),
.B(n_258),
.Y(n_3491)
);

O2A1O1Ixp33_ASAP7_75t_L g3492 ( 
.A1(n_3077),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_2900),
.A2(n_259),
.B(n_260),
.Y(n_3493)
);

AOI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_2901),
.A2(n_261),
.B(n_262),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3089),
.B(n_263),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_2736),
.A2(n_263),
.B(n_264),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_2740),
.A2(n_265),
.B(n_266),
.Y(n_3497)
);

OAI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_2707),
.A2(n_265),
.B(n_266),
.Y(n_3498)
);

AOI21x1_ASAP7_75t_L g3499 ( 
.A1(n_2876),
.A2(n_267),
.B(n_268),
.Y(n_3499)
);

CKINVDCx5p33_ASAP7_75t_R g3500 ( 
.A(n_3080),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_2734),
.B(n_267),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_2719),
.B(n_268),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3096),
.B(n_269),
.Y(n_3503)
);

O2A1O1Ixp33_ASAP7_75t_L g3504 ( 
.A1(n_3091),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_3504)
);

NAND3xp33_ASAP7_75t_L g3505 ( 
.A(n_2617),
.B(n_271),
.C(n_274),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3100),
.B(n_274),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_2741),
.A2(n_275),
.B(n_276),
.Y(n_3507)
);

AND2x2_ASAP7_75t_SL g3508 ( 
.A(n_2987),
.B(n_275),
.Y(n_3508)
);

AND2x4_ASAP7_75t_L g3509 ( 
.A(n_3169),
.B(n_276),
.Y(n_3509)
);

AOI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_2743),
.A2(n_277),
.B(n_278),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3101),
.B(n_277),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3104),
.Y(n_3512)
);

AO21x1_ASAP7_75t_L g3513 ( 
.A1(n_2894),
.A2(n_278),
.B(n_279),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3108),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3116),
.B(n_279),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_SL g3516 ( 
.A(n_2992),
.B(n_280),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_2665),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3517)
);

INVxp67_ASAP7_75t_L g3518 ( 
.A(n_3007),
.Y(n_3518)
);

O2A1O1Ixp33_ASAP7_75t_L g3519 ( 
.A1(n_3112),
.A2(n_284),
.B(n_281),
.C(n_283),
.Y(n_3519)
);

AND2x2_ASAP7_75t_SL g3520 ( 
.A(n_2748),
.B(n_283),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3117),
.Y(n_3521)
);

AOI22xp5_ASAP7_75t_L g3522 ( 
.A1(n_3001),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3522)
);

CKINVDCx20_ASAP7_75t_R g3523 ( 
.A(n_2831),
.Y(n_3523)
);

INVx1_ASAP7_75t_SL g3524 ( 
.A(n_2751),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_2800),
.A2(n_286),
.B(n_287),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_2804),
.A2(n_287),
.B(n_288),
.Y(n_3526)
);

BUFx6f_ASAP7_75t_L g3527 ( 
.A(n_2781),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_2807),
.A2(n_291),
.B(n_292),
.Y(n_3528)
);

BUFx2_ASAP7_75t_L g3529 ( 
.A(n_2683),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3121),
.Y(n_3530)
);

OAI21x1_ASAP7_75t_L g3531 ( 
.A1(n_2756),
.A2(n_291),
.B(n_292),
.Y(n_3531)
);

AO32x1_ASAP7_75t_L g3532 ( 
.A1(n_2878),
.A2(n_299),
.A3(n_295),
.B1(n_297),
.B2(n_300),
.Y(n_3532)
);

AOI33xp33_ASAP7_75t_L g3533 ( 
.A1(n_2666),
.A2(n_299),
.A3(n_302),
.B1(n_295),
.B2(n_297),
.B3(n_301),
.Y(n_3533)
);

BUFx12f_ASAP7_75t_L g3534 ( 
.A(n_3080),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3124),
.B(n_302),
.Y(n_3535)
);

O2A1O1Ixp33_ASAP7_75t_L g3536 ( 
.A1(n_3152),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3126),
.B(n_303),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_3129),
.B(n_304),
.Y(n_3538)
);

BUFx6f_ASAP7_75t_L g3539 ( 
.A(n_2827),
.Y(n_3539)
);

INVx2_ASAP7_75t_SL g3540 ( 
.A(n_2929),
.Y(n_3540)
);

INVx4_ASAP7_75t_L g3541 ( 
.A(n_2959),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3131),
.B(n_305),
.Y(n_3542)
);

A2O1A1Ixp33_ASAP7_75t_L g3543 ( 
.A1(n_3068),
.A2(n_309),
.B(n_307),
.C(n_308),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3132),
.B(n_3133),
.Y(n_3544)
);

AOI22xp5_ASAP7_75t_L g3545 ( 
.A1(n_3199),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3153),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_3007),
.B(n_310),
.Y(n_3547)
);

NOR2xp67_ASAP7_75t_L g3548 ( 
.A(n_2856),
.B(n_310),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_2818),
.A2(n_311),
.B(n_312),
.Y(n_3549)
);

AND2x4_ASAP7_75t_SL g3550 ( 
.A(n_2959),
.B(n_311),
.Y(n_3550)
);

AOI22xp5_ASAP7_75t_L g3551 ( 
.A1(n_3210),
.A2(n_315),
.B1(n_312),
.B2(n_313),
.Y(n_3551)
);

INVx4_ASAP7_75t_L g3552 ( 
.A(n_2727),
.Y(n_3552)
);

AOI21x1_ASAP7_75t_L g3553 ( 
.A1(n_2885),
.A2(n_313),
.B(n_316),
.Y(n_3553)
);

OA22x2_ASAP7_75t_L g3554 ( 
.A1(n_3084),
.A2(n_3176),
.B1(n_3171),
.B2(n_2894),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_2820),
.A2(n_316),
.B(n_317),
.Y(n_3555)
);

OAI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_2709),
.A2(n_317),
.B(n_319),
.Y(n_3556)
);

AOI22xp5_ASAP7_75t_L g3557 ( 
.A1(n_2774),
.A2(n_322),
.B1(n_319),
.B2(n_320),
.Y(n_3557)
);

AND2x2_ASAP7_75t_L g3558 ( 
.A(n_2775),
.B(n_320),
.Y(n_3558)
);

INVxp67_ASAP7_75t_L g3559 ( 
.A(n_3010),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3158),
.B(n_323),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3164),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_2821),
.A2(n_324),
.B(n_325),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3167),
.B(n_326),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3170),
.B(n_327),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_SL g3565 ( 
.A(n_3010),
.B(n_328),
.Y(n_3565)
);

BUFx8_ASAP7_75t_L g3566 ( 
.A(n_2879),
.Y(n_3566)
);

HB1xp67_ASAP7_75t_L g3567 ( 
.A(n_3071),
.Y(n_3567)
);

NOR3xp33_ASAP7_75t_L g3568 ( 
.A(n_2841),
.B(n_328),
.C(n_329),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3179),
.B(n_329),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_2822),
.A2(n_330),
.B(n_331),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_SL g3571 ( 
.A(n_3071),
.B(n_330),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3180),
.Y(n_3572)
);

AND2x4_ASAP7_75t_L g3573 ( 
.A(n_3206),
.B(n_331),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3214),
.B(n_332),
.Y(n_3574)
);

OAI22xp5_ASAP7_75t_L g3575 ( 
.A1(n_2665),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_3575)
);

INVx4_ASAP7_75t_L g3576 ( 
.A(n_3046),
.Y(n_3576)
);

AOI33xp33_ASAP7_75t_L g3577 ( 
.A1(n_2836),
.A2(n_336),
.A3(n_338),
.B1(n_333),
.B2(n_334),
.B3(n_337),
.Y(n_3577)
);

NAND2xp33_ASAP7_75t_L g3578 ( 
.A(n_2965),
.B(n_946),
.Y(n_3578)
);

OAI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_2691),
.A2(n_339),
.B(n_340),
.Y(n_3579)
);

AOI21xp5_ASAP7_75t_L g3580 ( 
.A1(n_2828),
.A2(n_339),
.B(n_341),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3215),
.B(n_342),
.Y(n_3581)
);

OAI21x1_ASAP7_75t_L g3582 ( 
.A1(n_2761),
.A2(n_343),
.B(n_344),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3219),
.B(n_344),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_L g3584 ( 
.A(n_2903),
.B(n_345),
.Y(n_3584)
);

NOR2xp67_ASAP7_75t_L g3585 ( 
.A(n_3184),
.B(n_345),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3221),
.B(n_346),
.Y(n_3586)
);

OAI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_2667),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_SL g3588 ( 
.A(n_3110),
.B(n_348),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3223),
.B(n_349),
.Y(n_3589)
);

AOI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_2632),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_3590)
);

A2O1A1Ixp33_ASAP7_75t_L g3591 ( 
.A1(n_3233),
.A2(n_353),
.B(n_351),
.C(n_352),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_2830),
.A2(n_353),
.B(n_354),
.Y(n_3592)
);

AO22x1_ASAP7_75t_L g3593 ( 
.A1(n_3213),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_2632),
.A2(n_361),
.B1(n_356),
.B2(n_360),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_2834),
.A2(n_361),
.B(n_362),
.Y(n_3595)
);

OAI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_2667),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_3596)
);

BUFx2_ASAP7_75t_L g3597 ( 
.A(n_2839),
.Y(n_3597)
);

AOI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_2837),
.A2(n_364),
.B(n_365),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3235),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_2775),
.B(n_366),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_SL g3601 ( 
.A(n_3110),
.B(n_367),
.Y(n_3601)
);

OAI22xp5_ASAP7_75t_L g3602 ( 
.A1(n_2825),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_2910),
.A2(n_2923),
.B(n_2873),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_2662),
.A2(n_368),
.B(n_369),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3236),
.B(n_370),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_2663),
.Y(n_3606)
);

O2A1O1Ixp33_ASAP7_75t_L g3607 ( 
.A1(n_2779),
.A2(n_373),
.B(n_371),
.C(n_372),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_2669),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_2671),
.A2(n_371),
.B(n_375),
.Y(n_3609)
);

AOI21xp5_ASAP7_75t_L g3610 ( 
.A1(n_2672),
.A2(n_377),
.B(n_378),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_2673),
.A2(n_379),
.B(n_380),
.Y(n_3611)
);

AND2x4_ASAP7_75t_L g3612 ( 
.A(n_2790),
.B(n_379),
.Y(n_3612)
);

OAI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_2972),
.A2(n_380),
.B(n_381),
.Y(n_3613)
);

AND2x2_ASAP7_75t_L g3614 ( 
.A(n_3034),
.B(n_381),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_SL g3615 ( 
.A(n_3128),
.B(n_383),
.Y(n_3615)
);

AOI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_2684),
.A2(n_384),
.B(n_385),
.Y(n_3616)
);

INVx2_ASAP7_75t_SL g3617 ( 
.A(n_2929),
.Y(n_3617)
);

NOR2xp33_ASAP7_75t_L g3618 ( 
.A(n_2726),
.B(n_2926),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_2694),
.Y(n_3619)
);

O2A1O1Ixp33_ASAP7_75t_L g3620 ( 
.A1(n_2695),
.A2(n_387),
.B(n_384),
.C(n_386),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_2705),
.A2(n_387),
.B(n_388),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_SL g3622 ( 
.A(n_3128),
.B(n_388),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2941),
.A2(n_389),
.B(n_390),
.Y(n_3623)
);

BUFx2_ASAP7_75t_L g3624 ( 
.A(n_2880),
.Y(n_3624)
);

AOI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_2936),
.A2(n_389),
.B(n_390),
.Y(n_3625)
);

O2A1O1Ixp5_ASAP7_75t_L g3626 ( 
.A1(n_2887),
.A2(n_393),
.B(n_391),
.C(n_392),
.Y(n_3626)
);

OAI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_2682),
.A2(n_391),
.B(n_392),
.Y(n_3627)
);

AOI22xp5_ASAP7_75t_L g3628 ( 
.A1(n_2753),
.A2(n_395),
.B1(n_393),
.B2(n_394),
.Y(n_3628)
);

AO22x1_ASAP7_75t_L g3629 ( 
.A1(n_2965),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_2937),
.B(n_396),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_2924),
.A2(n_397),
.B(n_398),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_SL g3632 ( 
.A(n_3138),
.B(n_398),
.Y(n_3632)
);

AOI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_2931),
.A2(n_399),
.B(n_401),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_2942),
.B(n_399),
.Y(n_3634)
);

AOI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_2899),
.A2(n_401),
.B(n_402),
.Y(n_3635)
);

INVxp67_ASAP7_75t_L g3636 ( 
.A(n_3138),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_2944),
.B(n_402),
.Y(n_3637)
);

BUFx6f_ASAP7_75t_L g3638 ( 
.A(n_2962),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_2907),
.A2(n_403),
.B(n_404),
.Y(n_3639)
);

A2O1A1Ixp33_ASAP7_75t_L g3640 ( 
.A1(n_2686),
.A2(n_409),
.B(n_406),
.C(n_408),
.Y(n_3640)
);

AOI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_2957),
.A2(n_408),
.B(n_409),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_2945),
.B(n_410),
.Y(n_3642)
);

O2A1O1Ixp33_ASAP7_75t_SL g3643 ( 
.A1(n_2890),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_2917),
.A2(n_412),
.B(n_413),
.Y(n_3644)
);

A2O1A1Ixp33_ASAP7_75t_L g3645 ( 
.A1(n_2675),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_3645)
);

OR2x6_ASAP7_75t_L g3646 ( 
.A(n_3038),
.B(n_415),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_2958),
.B(n_416),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_2967),
.B(n_2974),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_2864),
.Y(n_3649)
);

NAND2x1p5_ASAP7_75t_L g3650 ( 
.A(n_2606),
.B(n_417),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3052),
.B(n_417),
.Y(n_3651)
);

A2O1A1Ixp33_ASAP7_75t_L g3652 ( 
.A1(n_2675),
.A2(n_420),
.B(n_418),
.C(n_419),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_SL g3653 ( 
.A(n_3162),
.B(n_418),
.Y(n_3653)
);

INVxp67_ASAP7_75t_L g3654 ( 
.A(n_3162),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_2911),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3105),
.B(n_421),
.Y(n_3656)
);

NAND3xp33_ASAP7_75t_L g3657 ( 
.A(n_2918),
.B(n_422),
.C(n_423),
.Y(n_3657)
);

INVx3_ASAP7_75t_L g3658 ( 
.A(n_2904),
.Y(n_3658)
);

AOI22xp33_ASAP7_75t_L g3659 ( 
.A1(n_2791),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_3659)
);

AOI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_2780),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_SL g3661 ( 
.A(n_3187),
.B(n_425),
.Y(n_3661)
);

INVx3_ASAP7_75t_L g3662 ( 
.A(n_2616),
.Y(n_3662)
);

INVx2_ASAP7_75t_L g3663 ( 
.A(n_2746),
.Y(n_3663)
);

AND2x2_ASAP7_75t_L g3664 ( 
.A(n_3123),
.B(n_3157),
.Y(n_3664)
);

A2O1A1Ixp33_ASAP7_75t_L g3665 ( 
.A1(n_2676),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_3665)
);

OAI21xp33_ASAP7_75t_L g3666 ( 
.A1(n_2808),
.A2(n_2631),
.B(n_2703),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3181),
.B(n_428),
.Y(n_3667)
);

CKINVDCx5p33_ASAP7_75t_R g3668 ( 
.A(n_2764),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_2762),
.A2(n_429),
.B(n_430),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3205),
.B(n_429),
.Y(n_3670)
);

NOR2xp33_ASAP7_75t_L g3671 ( 
.A(n_2840),
.B(n_2845),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_2763),
.A2(n_431),
.B(n_432),
.Y(n_3672)
);

OAI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_2913),
.A2(n_432),
.B(n_433),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_2769),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_2966),
.B(n_434),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_2925),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_2846),
.B(n_2850),
.Y(n_3677)
);

AOI21xp5_ASAP7_75t_L g3678 ( 
.A1(n_2771),
.A2(n_434),
.B(n_436),
.Y(n_3678)
);

INVx4_ASAP7_75t_L g3679 ( 
.A(n_2799),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_2920),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_2857),
.B(n_436),
.Y(n_3681)
);

AOI22xp33_ASAP7_75t_L g3682 ( 
.A1(n_2791),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_3682)
);

AND2x2_ASAP7_75t_L g3683 ( 
.A(n_2927),
.B(n_437),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_2783),
.Y(n_3684)
);

OR2x2_ASAP7_75t_L g3685 ( 
.A(n_2813),
.B(n_438),
.Y(n_3685)
);

AOI21xp5_ASAP7_75t_L g3686 ( 
.A1(n_2789),
.A2(n_439),
.B(n_441),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_2798),
.B(n_441),
.Y(n_3687)
);

INVxp67_ASAP7_75t_L g3688 ( 
.A(n_3187),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_2905),
.A2(n_442),
.B(n_444),
.Y(n_3689)
);

OAI321xp33_ASAP7_75t_L g3690 ( 
.A1(n_3049),
.A2(n_445),
.A3(n_447),
.B1(n_442),
.B2(n_444),
.C(n_446),
.Y(n_3690)
);

O2A1O1Ixp33_ASAP7_75t_L g3691 ( 
.A1(n_2916),
.A2(n_447),
.B(n_445),
.C(n_446),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_2906),
.A2(n_448),
.B(n_449),
.Y(n_3692)
);

OAI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_3012),
.A2(n_451),
.B1(n_448),
.B2(n_450),
.Y(n_3693)
);

O2A1O1Ixp33_ASAP7_75t_L g3694 ( 
.A1(n_2714),
.A2(n_453),
.B(n_451),
.C(n_452),
.Y(n_3694)
);

NOR2xp67_ASAP7_75t_L g3695 ( 
.A(n_3041),
.B(n_452),
.Y(n_3695)
);

AOI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_2938),
.A2(n_454),
.B(n_455),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_2940),
.A2(n_454),
.B(n_455),
.Y(n_3697)
);

BUFx3_ASAP7_75t_L g3698 ( 
.A(n_2879),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_2801),
.B(n_2946),
.Y(n_3699)
);

BUFx2_ASAP7_75t_L g3700 ( 
.A(n_2872),
.Y(n_3700)
);

INVx3_ASAP7_75t_L g3701 ( 
.A(n_2687),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_2920),
.Y(n_3702)
);

AOI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_2982),
.A2(n_456),
.B(n_457),
.Y(n_3703)
);

NOR2xp33_ASAP7_75t_L g3704 ( 
.A(n_2738),
.B(n_2720),
.Y(n_3704)
);

OAI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_2855),
.A2(n_456),
.B(n_458),
.Y(n_3705)
);

AOI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_2747),
.A2(n_458),
.B(n_459),
.Y(n_3706)
);

AOI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_2773),
.A2(n_460),
.B(n_461),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_2776),
.A2(n_460),
.B(n_461),
.Y(n_3708)
);

CKINVDCx10_ASAP7_75t_R g3709 ( 
.A(n_2619),
.Y(n_3709)
);

AND2x2_ASAP7_75t_SL g3710 ( 
.A(n_3204),
.B(n_462),
.Y(n_3710)
);

HB1xp67_ASAP7_75t_L g3711 ( 
.A(n_3204),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_2969),
.A2(n_463),
.B(n_464),
.Y(n_3712)
);

AOI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_2983),
.A2(n_464),
.B(n_465),
.Y(n_3713)
);

O2A1O1Ixp33_ASAP7_75t_L g3714 ( 
.A1(n_2757),
.A2(n_2657),
.B(n_3061),
.C(n_3039),
.Y(n_3714)
);

OAI22xp5_ASAP7_75t_L g3715 ( 
.A1(n_3114),
.A2(n_3122),
.B1(n_3149),
.B2(n_3120),
.Y(n_3715)
);

AOI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_2909),
.A2(n_465),
.B(n_466),
.Y(n_3716)
);

OAI321xp33_ASAP7_75t_L g3717 ( 
.A1(n_3050),
.A2(n_469),
.A3(n_471),
.B1(n_467),
.B2(n_468),
.C(n_470),
.Y(n_3717)
);

AOI21xp33_ASAP7_75t_L g3718 ( 
.A1(n_2724),
.A2(n_470),
.B(n_471),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_2725),
.B(n_2752),
.Y(n_3719)
);

BUFx6f_ASAP7_75t_L g3720 ( 
.A(n_2796),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_2892),
.A2(n_472),
.B(n_473),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_2725),
.B(n_472),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_2802),
.B(n_473),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3207),
.Y(n_3724)
);

NOR2xp67_ASAP7_75t_L g3725 ( 
.A(n_3059),
.B(n_474),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_2752),
.B(n_476),
.Y(n_3726)
);

AOI21xp5_ASAP7_75t_L g3727 ( 
.A1(n_2895),
.A2(n_476),
.B(n_477),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_2927),
.B(n_477),
.Y(n_3728)
);

OAI321xp33_ASAP7_75t_L g3729 ( 
.A1(n_3098),
.A2(n_480),
.A3(n_482),
.B1(n_478),
.B2(n_479),
.C(n_481),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3207),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_2676),
.B(n_2770),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_2770),
.B(n_478),
.Y(n_3732)
);

NOR2xp33_ASAP7_75t_R g3733 ( 
.A(n_2835),
.B(n_947),
.Y(n_3733)
);

INVx3_ASAP7_75t_L g3734 ( 
.A(n_2700),
.Y(n_3734)
);

NOR2xp33_ASAP7_75t_L g3735 ( 
.A(n_2802),
.B(n_482),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_2961),
.B(n_483),
.Y(n_3736)
);

INVx3_ASAP7_75t_L g3737 ( 
.A(n_2716),
.Y(n_3737)
);

AOI21x1_ASAP7_75t_L g3738 ( 
.A1(n_2932),
.A2(n_483),
.B(n_484),
.Y(n_3738)
);

OAI21xp5_ASAP7_75t_L g3739 ( 
.A1(n_2973),
.A2(n_485),
.B(n_487),
.Y(n_3739)
);

AOI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_2978),
.A2(n_487),
.B(n_488),
.Y(n_3740)
);

OAI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_2708),
.A2(n_489),
.B(n_490),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_2730),
.A2(n_489),
.B(n_494),
.Y(n_3742)
);

OR2x6_ASAP7_75t_L g3743 ( 
.A(n_3107),
.B(n_495),
.Y(n_3743)
);

INVx3_ASAP7_75t_L g3744 ( 
.A(n_3212),
.Y(n_3744)
);

O2A1O1Ixp33_ASAP7_75t_L g3745 ( 
.A1(n_2648),
.A2(n_497),
.B(n_495),
.C(n_496),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_2765),
.A2(n_496),
.B(n_497),
.Y(n_3746)
);

NOR2x1p5_ASAP7_75t_L g3747 ( 
.A(n_2956),
.B(n_498),
.Y(n_3747)
);

OAI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_2612),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_2981),
.A2(n_499),
.B(n_501),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_SL g3750 ( 
.A(n_3212),
.B(n_501),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3217),
.Y(n_3751)
);

OAI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_2977),
.A2(n_502),
.B(n_503),
.Y(n_3752)
);

OAI22xp5_ASAP7_75t_L g3753 ( 
.A1(n_2797),
.A2(n_2851),
.B1(n_2877),
.B2(n_2698),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_2621),
.A2(n_503),
.B(n_504),
.Y(n_3754)
);

OAI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_2980),
.A2(n_2599),
.B(n_2809),
.Y(n_3755)
);

AOI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_2932),
.A2(n_504),
.B(n_505),
.Y(n_3756)
);

O2A1O1Ixp5_ASAP7_75t_L g3757 ( 
.A1(n_2778),
.A2(n_507),
.B(n_505),
.C(n_506),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_2947),
.B(n_506),
.Y(n_3758)
);

O2A1O1Ixp33_ASAP7_75t_L g3759 ( 
.A1(n_2668),
.A2(n_3000),
.B(n_2608),
.C(n_2848),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_2943),
.A2(n_509),
.B(n_510),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3217),
.B(n_510),
.Y(n_3761)
);

BUFx2_ASAP7_75t_L g3762 ( 
.A(n_2954),
.Y(n_3762)
);

AOI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_2618),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_3763)
);

AOI21xp5_ASAP7_75t_L g3764 ( 
.A1(n_2943),
.A2(n_513),
.B(n_514),
.Y(n_3764)
);

OAI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_2599),
.A2(n_515),
.B(n_516),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_2718),
.A2(n_515),
.B(n_516),
.Y(n_3766)
);

OAI21xp33_ASAP7_75t_L g3767 ( 
.A1(n_2795),
.A2(n_517),
.B(n_518),
.Y(n_3767)
);

NAND3xp33_ASAP7_75t_L g3768 ( 
.A(n_2824),
.B(n_518),
.C(n_519),
.Y(n_3768)
);

AOI21xp5_ASAP7_75t_L g3769 ( 
.A1(n_3072),
.A2(n_519),
.B(n_520),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3224),
.B(n_520),
.Y(n_3770)
);

AND2x4_ASAP7_75t_L g3771 ( 
.A(n_3160),
.B(n_521),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3224),
.Y(n_3772)
);

NOR2xp33_ASAP7_75t_L g3773 ( 
.A(n_2859),
.B(n_521),
.Y(n_3773)
);

AOI21xp5_ASAP7_75t_L g3774 ( 
.A1(n_3163),
.A2(n_523),
.B(n_524),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3232),
.B(n_523),
.Y(n_3775)
);

OAI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_2809),
.A2(n_2810),
.B(n_2758),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3232),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_SL g3778 ( 
.A(n_3237),
.B(n_524),
.Y(n_3778)
);

NOR3xp33_ASAP7_75t_L g3779 ( 
.A(n_2881),
.B(n_525),
.C(n_526),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3237),
.B(n_525),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_2851),
.Y(n_3781)
);

NAND3xp33_ASAP7_75t_L g3782 ( 
.A(n_2685),
.B(n_526),
.C(n_527),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3196),
.B(n_2797),
.Y(n_3783)
);

AOI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_2651),
.A2(n_527),
.B(n_528),
.Y(n_3784)
);

O2A1O1Ixp33_ASAP7_75t_L g3785 ( 
.A1(n_3753),
.A2(n_3228),
.B(n_3197),
.C(n_3155),
.Y(n_3785)
);

O2A1O1Ixp33_ASAP7_75t_L g3786 ( 
.A1(n_3341),
.A2(n_3140),
.B(n_2884),
.C(n_2787),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_3257),
.A2(n_2996),
.B(n_2994),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3246),
.Y(n_3788)
);

O2A1O1Ixp33_ASAP7_75t_L g3789 ( 
.A1(n_3666),
.A2(n_2815),
.B(n_2609),
.C(n_2611),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3284),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3655),
.Y(n_3791)
);

AOI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3266),
.A2(n_2996),
.B(n_2994),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3664),
.B(n_2795),
.Y(n_3793)
);

O2A1O1Ixp33_ASAP7_75t_L g3794 ( 
.A1(n_3699),
.A2(n_2951),
.B(n_2891),
.C(n_3005),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3508),
.B(n_2877),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3311),
.B(n_2698),
.Y(n_3796)
);

AND2x4_ASAP7_75t_L g3797 ( 
.A(n_3323),
.B(n_2742),
.Y(n_3797)
);

AOI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_3280),
.A2(n_3029),
.B(n_3015),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3475),
.B(n_2914),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_R g3800 ( 
.A(n_3523),
.B(n_3500),
.Y(n_3800)
);

A2O1A1Ixp33_ASAP7_75t_SL g3801 ( 
.A1(n_3584),
.A2(n_2915),
.B(n_2993),
.C(n_2970),
.Y(n_3801)
);

NOR2xp67_ASAP7_75t_SL g3802 ( 
.A(n_3249),
.B(n_3065),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3578),
.A2(n_3029),
.B(n_3015),
.Y(n_3803)
);

AOI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_3240),
.A2(n_3064),
.B(n_3036),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3239),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3648),
.Y(n_3806)
);

AND2x4_ASAP7_75t_L g3807 ( 
.A(n_3354),
.B(n_2759),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3649),
.Y(n_3808)
);

INVx8_ASAP7_75t_L g3809 ( 
.A(n_3433),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3337),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3389),
.B(n_3430),
.Y(n_3811)
);

NAND2xp33_ASAP7_75t_SL g3812 ( 
.A(n_3437),
.B(n_2766),
.Y(n_3812)
);

NOR3xp33_ASAP7_75t_SL g3813 ( 
.A(n_3668),
.B(n_2964),
.C(n_3042),
.Y(n_3813)
);

NAND2x1p5_ASAP7_75t_L g3814 ( 
.A(n_3473),
.B(n_2843),
.Y(n_3814)
);

BUFx2_ASAP7_75t_L g3815 ( 
.A(n_3700),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3275),
.A2(n_3064),
.B(n_3036),
.Y(n_3816)
);

INVx1_ASAP7_75t_SL g3817 ( 
.A(n_3427),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3436),
.A2(n_3079),
.B(n_3075),
.Y(n_3818)
);

AOI21x1_ASAP7_75t_L g3819 ( 
.A1(n_3238),
.A2(n_3079),
.B(n_3075),
.Y(n_3819)
);

BUFx6f_ASAP7_75t_L g3820 ( 
.A(n_3483),
.Y(n_3820)
);

A2O1A1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_3276),
.A2(n_2891),
.B(n_2618),
.C(n_2652),
.Y(n_3821)
);

OAI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_3710),
.A2(n_2914),
.B1(n_2646),
.B2(n_3113),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_SL g3823 ( 
.A(n_3437),
.B(n_2919),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3443),
.Y(n_3824)
);

AND2x4_ASAP7_75t_L g3825 ( 
.A(n_3658),
.B(n_3427),
.Y(n_3825)
);

AND2x4_ASAP7_75t_L g3826 ( 
.A(n_3658),
.B(n_3087),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3448),
.B(n_2737),
.Y(n_3827)
);

A2O1A1Ixp33_ASAP7_75t_L g3828 ( 
.A1(n_3278),
.A2(n_2651),
.B(n_2652),
.C(n_2643),
.Y(n_3828)
);

BUFx3_ASAP7_75t_L g3829 ( 
.A(n_3566),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3450),
.Y(n_3830)
);

O2A1O1Ixp33_ASAP7_75t_L g3831 ( 
.A1(n_3367),
.A2(n_2737),
.B(n_2739),
.C(n_2643),
.Y(n_3831)
);

NOR2xp33_ASAP7_75t_L g3832 ( 
.A(n_3242),
.B(n_2603),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3441),
.A2(n_3141),
.B(n_3113),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_R g3834 ( 
.A(n_3709),
.B(n_2919),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3319),
.A2(n_3145),
.B(n_3141),
.Y(n_3835)
);

NOR2xp33_ASAP7_75t_L g3836 ( 
.A(n_3618),
.B(n_2986),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3461),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3331),
.A2(n_3159),
.B(n_3145),
.Y(n_3838)
);

AOI22xp5_ASAP7_75t_L g3839 ( 
.A1(n_3554),
.A2(n_2647),
.B1(n_2739),
.B2(n_2636),
.Y(n_3839)
);

AO31x2_ASAP7_75t_L g3840 ( 
.A1(n_3680),
.A2(n_2948),
.A3(n_2955),
.B(n_2960),
.Y(n_3840)
);

BUFx8_ASAP7_75t_L g3841 ( 
.A(n_3534),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3437),
.B(n_3102),
.Y(n_3842)
);

AOI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3783),
.A2(n_2636),
.B1(n_2622),
.B2(n_3200),
.Y(n_3843)
);

NOR3xp33_ASAP7_75t_SL g3844 ( 
.A(n_3767),
.B(n_3177),
.C(n_3060),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3340),
.A2(n_3165),
.B(n_3159),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3420),
.Y(n_3846)
);

HB1xp67_ASAP7_75t_L g3847 ( 
.A(n_3452),
.Y(n_3847)
);

NOR2xp67_ASAP7_75t_L g3848 ( 
.A(n_3451),
.B(n_3150),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3349),
.A2(n_3200),
.B(n_3165),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3439),
.Y(n_3850)
);

AOI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3603),
.A2(n_3225),
.B(n_3216),
.Y(n_3851)
);

INVx1_ASAP7_75t_SL g3852 ( 
.A(n_3424),
.Y(n_3852)
);

INVx4_ASAP7_75t_L g3853 ( 
.A(n_3346),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3512),
.B(n_2810),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3501),
.B(n_3216),
.Y(n_3855)
);

HB1xp67_ASAP7_75t_L g3856 ( 
.A(n_3244),
.Y(n_3856)
);

NAND2x1p5_ASAP7_75t_L g3857 ( 
.A(n_3392),
.B(n_2930),
.Y(n_3857)
);

AOI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3364),
.A2(n_2622),
.B1(n_2979),
.B2(n_2689),
.Y(n_3858)
);

NOR2xp33_ASAP7_75t_R g3859 ( 
.A(n_3260),
.B(n_3156),
.Y(n_3859)
);

NOR2xp33_ASAP7_75t_L g3860 ( 
.A(n_3518),
.B(n_2829),
.Y(n_3860)
);

INVx2_ASAP7_75t_L g3861 ( 
.A(n_3457),
.Y(n_3861)
);

BUFx2_ASAP7_75t_L g3862 ( 
.A(n_3392),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3558),
.B(n_3225),
.Y(n_3863)
);

NOR2xp33_ASAP7_75t_L g3864 ( 
.A(n_3559),
.B(n_3636),
.Y(n_3864)
);

O2A1O1Ixp33_ASAP7_75t_L g3865 ( 
.A1(n_3292),
.A2(n_3188),
.B(n_2689),
.C(n_2677),
.Y(n_3865)
);

NOR2xp33_ASAP7_75t_L g3866 ( 
.A(n_3654),
.B(n_2677),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3440),
.B(n_3539),
.Y(n_3867)
);

AOI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3470),
.A2(n_3226),
.B(n_2963),
.Y(n_3868)
);

AOI21xp5_ASAP7_75t_L g3869 ( 
.A1(n_3445),
.A2(n_3256),
.B(n_3304),
.Y(n_3869)
);

A2O1A1Ixp33_ASAP7_75t_SL g3870 ( 
.A1(n_3476),
.A2(n_2975),
.B(n_2826),
.C(n_2861),
.Y(n_3870)
);

INVxp67_ASAP7_75t_L g3871 ( 
.A(n_3379),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3521),
.B(n_2949),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_SL g3873 ( 
.A(n_3440),
.B(n_3539),
.Y(n_3873)
);

O2A1O1Ixp33_ASAP7_75t_L g3874 ( 
.A1(n_3714),
.A2(n_3226),
.B(n_2965),
.C(n_533),
.Y(n_3874)
);

AOI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3449),
.A2(n_530),
.B(n_531),
.Y(n_3875)
);

O2A1O1Ixp33_ASAP7_75t_L g3876 ( 
.A1(n_3759),
.A2(n_534),
.B(n_531),
.C(n_533),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3546),
.Y(n_3877)
);

AOI21xp5_ASAP7_75t_L g3878 ( 
.A1(n_3434),
.A2(n_535),
.B(n_536),
.Y(n_3878)
);

INVx11_ASAP7_75t_L g3879 ( 
.A(n_3316),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3561),
.B(n_535),
.Y(n_3880)
);

CKINVDCx16_ASAP7_75t_R g3881 ( 
.A(n_3379),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3572),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3599),
.B(n_537),
.Y(n_3883)
);

NOR2xp33_ASAP7_75t_SL g3884 ( 
.A(n_3396),
.B(n_537),
.Y(n_3884)
);

O2A1O1Ixp33_ASAP7_75t_SL g3885 ( 
.A1(n_3645),
.A2(n_540),
.B(n_538),
.C(n_539),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3600),
.B(n_538),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_3619),
.B(n_539),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_L g3888 ( 
.A(n_3688),
.B(n_540),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3715),
.A2(n_541),
.B(n_542),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3676),
.Y(n_3890)
);

BUFx2_ASAP7_75t_L g3891 ( 
.A(n_3451),
.Y(n_3891)
);

CKINVDCx16_ASAP7_75t_R g3892 ( 
.A(n_3310),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3418),
.B(n_541),
.Y(n_3893)
);

BUFx3_ASAP7_75t_L g3894 ( 
.A(n_3566),
.Y(n_3894)
);

BUFx6f_ASAP7_75t_L g3895 ( 
.A(n_3362),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3544),
.B(n_542),
.Y(n_3896)
);

AOI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3308),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_3897)
);

AOI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_3469),
.A2(n_543),
.B(n_544),
.Y(n_3898)
);

NAND2x1p5_ASAP7_75t_L g3899 ( 
.A(n_3679),
.B(n_545),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3781),
.B(n_546),
.Y(n_3900)
);

INVx2_ASAP7_75t_L g3901 ( 
.A(n_3459),
.Y(n_3901)
);

BUFx6f_ASAP7_75t_L g3902 ( 
.A(n_3362),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3731),
.B(n_3719),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_SL g3904 ( 
.A(n_3440),
.B(n_546),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3478),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3486),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3282),
.A2(n_547),
.B(n_548),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3488),
.B(n_547),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_SL g3909 ( 
.A(n_3539),
.B(n_548),
.Y(n_3909)
);

NOR3xp33_ASAP7_75t_SL g3910 ( 
.A(n_3468),
.B(n_549),
.C(n_550),
.Y(n_3910)
);

NOR2xp33_ASAP7_75t_L g3911 ( 
.A(n_3755),
.B(n_549),
.Y(n_3911)
);

AOI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3243),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_SL g3913 ( 
.A(n_3638),
.B(n_554),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3514),
.Y(n_3914)
);

HB1xp67_ASAP7_75t_L g3915 ( 
.A(n_3567),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3530),
.Y(n_3916)
);

OAI22xp5_ASAP7_75t_L g3917 ( 
.A1(n_3573),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3606),
.Y(n_3918)
);

AOI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_3394),
.A2(n_555),
.B(n_556),
.Y(n_3919)
);

OAI22xp5_ASAP7_75t_SL g3920 ( 
.A1(n_3520),
.A2(n_561),
.B1(n_559),
.B2(n_560),
.Y(n_3920)
);

OAI22xp5_ASAP7_75t_L g3921 ( 
.A1(n_3573),
.A2(n_562),
.B1(n_559),
.B2(n_560),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3608),
.B(n_563),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3245),
.A2(n_563),
.B(n_564),
.Y(n_3923)
);

INVx3_ASAP7_75t_L g3924 ( 
.A(n_3552),
.Y(n_3924)
);

NOR2xp33_ASAP7_75t_L g3925 ( 
.A(n_3711),
.B(n_565),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3252),
.Y(n_3926)
);

NOR2xp67_ASAP7_75t_SL g3927 ( 
.A(n_3762),
.B(n_566),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3247),
.A2(n_567),
.B(n_568),
.Y(n_3928)
);

CKINVDCx5p33_ASAP7_75t_R g3929 ( 
.A(n_3316),
.Y(n_3929)
);

AOI211xp5_ASAP7_75t_L g3930 ( 
.A1(n_3693),
.A2(n_570),
.B(n_567),
.C(n_569),
.Y(n_3930)
);

AND2x4_ASAP7_75t_L g3931 ( 
.A(n_3310),
.B(n_570),
.Y(n_3931)
);

AOI22xp5_ASAP7_75t_L g3932 ( 
.A1(n_3334),
.A2(n_3347),
.B1(n_3568),
.B2(n_3303),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3254),
.B(n_571),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3277),
.B(n_571),
.Y(n_3934)
);

AOI21xp5_ASAP7_75t_L g3935 ( 
.A1(n_3356),
.A2(n_3643),
.B(n_3255),
.Y(n_3935)
);

O2A1O1Ixp33_ASAP7_75t_L g3936 ( 
.A1(n_3482),
.A2(n_575),
.B(n_572),
.C(n_574),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3306),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_3250),
.A2(n_572),
.B(n_574),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3315),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3336),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3663),
.Y(n_3941)
);

CKINVDCx8_ASAP7_75t_R g3942 ( 
.A(n_3328),
.Y(n_3942)
);

AOI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_3302),
.A2(n_575),
.B(n_576),
.Y(n_3943)
);

AOI21xp5_ASAP7_75t_L g3944 ( 
.A1(n_3375),
.A2(n_576),
.B(n_577),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_SL g3945 ( 
.A(n_3638),
.B(n_578),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3677),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3638),
.B(n_578),
.Y(n_3947)
);

BUFx12f_ASAP7_75t_L g3948 ( 
.A(n_3453),
.Y(n_3948)
);

BUFx6f_ASAP7_75t_L g3949 ( 
.A(n_3362),
.Y(n_3949)
);

O2A1O1Ixp33_ASAP7_75t_L g3950 ( 
.A1(n_3516),
.A2(n_3547),
.B(n_3588),
.C(n_3565),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3376),
.Y(n_3951)
);

NOR2xp33_ASAP7_75t_L g3952 ( 
.A(n_3597),
.B(n_579),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3263),
.Y(n_3953)
);

AOI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3390),
.A2(n_579),
.B(n_580),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3401),
.Y(n_3955)
);

AOI22xp5_ASAP7_75t_L g3956 ( 
.A1(n_3360),
.A2(n_584),
.B1(n_580),
.B2(n_583),
.Y(n_3956)
);

BUFx12f_ASAP7_75t_L g3957 ( 
.A(n_3529),
.Y(n_3957)
);

O2A1O1Ixp33_ASAP7_75t_L g3958 ( 
.A1(n_3571),
.A2(n_587),
.B(n_584),
.C(n_585),
.Y(n_3958)
);

OAI22xp5_ASAP7_75t_L g3959 ( 
.A1(n_3463),
.A2(n_589),
.B1(n_585),
.B2(n_588),
.Y(n_3959)
);

AOI21xp5_ASAP7_75t_L g3960 ( 
.A1(n_3744),
.A2(n_3417),
.B(n_3312),
.Y(n_3960)
);

NOR2xp33_ASAP7_75t_L g3961 ( 
.A(n_3624),
.B(n_590),
.Y(n_3961)
);

BUFx6f_ASAP7_75t_L g3962 ( 
.A(n_3698),
.Y(n_3962)
);

INVxp67_ASAP7_75t_L g3963 ( 
.A(n_3704),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3744),
.A2(n_590),
.B(n_591),
.Y(n_3964)
);

O2A1O1Ixp33_ASAP7_75t_L g3965 ( 
.A1(n_3601),
.A2(n_595),
.B(n_591),
.C(n_594),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3671),
.B(n_595),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3267),
.Y(n_3967)
);

AOI221xp5_ASAP7_75t_L g3968 ( 
.A1(n_3294),
.A2(n_598),
.B1(n_596),
.B2(n_597),
.C(n_599),
.Y(n_3968)
);

BUFx3_ASAP7_75t_L g3969 ( 
.A(n_3541),
.Y(n_3969)
);

AOI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_3723),
.A2(n_3735),
.B1(n_3502),
.B2(n_3371),
.Y(n_3970)
);

OAI22x1_ASAP7_75t_L g3971 ( 
.A1(n_3747),
.A2(n_3406),
.B1(n_3509),
.B2(n_3650),
.Y(n_3971)
);

BUFx6f_ASAP7_75t_L g3972 ( 
.A(n_3720),
.Y(n_3972)
);

BUFx5_ASAP7_75t_L g3973 ( 
.A(n_3258),
.Y(n_3973)
);

BUFx2_ASAP7_75t_L g3974 ( 
.A(n_3576),
.Y(n_3974)
);

NOR2xp33_ASAP7_75t_L g3975 ( 
.A(n_3524),
.B(n_3423),
.Y(n_3975)
);

O2A1O1Ixp33_ASAP7_75t_L g3976 ( 
.A1(n_3615),
.A2(n_602),
.B(n_600),
.C(n_601),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3241),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3531),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_SL g3979 ( 
.A(n_3429),
.B(n_604),
.Y(n_3979)
);

NAND2x1_ASAP7_75t_L g3980 ( 
.A(n_3307),
.B(n_604),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_3582),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_3776),
.B(n_951),
.Y(n_3982)
);

A2O1A1Ixp33_ASAP7_75t_L g3983 ( 
.A1(n_3301),
.A2(n_608),
.B(n_606),
.C(n_607),
.Y(n_3983)
);

BUFx3_ASAP7_75t_L g3984 ( 
.A(n_3541),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3259),
.A2(n_606),
.B(n_607),
.Y(n_3985)
);

HB1xp67_ASAP7_75t_L g3986 ( 
.A(n_3724),
.Y(n_3986)
);

OR2x6_ASAP7_75t_SL g3987 ( 
.A(n_3309),
.B(n_608),
.Y(n_3987)
);

INVx2_ASAP7_75t_SL g3988 ( 
.A(n_3720),
.Y(n_3988)
);

HB1xp67_ASAP7_75t_L g3989 ( 
.A(n_3730),
.Y(n_3989)
);

AND2x6_ASAP7_75t_L g3990 ( 
.A(n_3702),
.B(n_609),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_3756),
.A2(n_609),
.B(n_610),
.Y(n_3991)
);

O2A1O1Ixp33_ASAP7_75t_L g3992 ( 
.A1(n_3622),
.A2(n_612),
.B(n_610),
.C(n_611),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3274),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3279),
.Y(n_3994)
);

AOI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3760),
.A2(n_611),
.B(n_613),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3286),
.Y(n_3996)
);

BUFx3_ASAP7_75t_L g3997 ( 
.A(n_3720),
.Y(n_3997)
);

NOR2xp33_ASAP7_75t_L g3998 ( 
.A(n_3772),
.B(n_613),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3751),
.B(n_951),
.Y(n_3999)
);

INVx1_ASAP7_75t_SL g4000 ( 
.A(n_3431),
.Y(n_4000)
);

AND2x4_ASAP7_75t_L g4001 ( 
.A(n_3463),
.B(n_614),
.Y(n_4001)
);

INVx3_ASAP7_75t_L g4002 ( 
.A(n_3552),
.Y(n_4002)
);

A2O1A1Ixp33_ASAP7_75t_L g4003 ( 
.A1(n_3305),
.A2(n_616),
.B(n_614),
.C(n_615),
.Y(n_4003)
);

BUFx2_ASAP7_75t_L g4004 ( 
.A(n_3576),
.Y(n_4004)
);

INVx2_ASAP7_75t_SL g4005 ( 
.A(n_3540),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3764),
.A2(n_615),
.B(n_617),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3291),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_L g4008 ( 
.A(n_3679),
.B(n_617),
.Y(n_4008)
);

CKINVDCx20_ASAP7_75t_R g4009 ( 
.A(n_3296),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3253),
.B(n_618),
.Y(n_4010)
);

OAI22xp5_ASAP7_75t_L g4011 ( 
.A1(n_3646),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_4011)
);

AOI22xp5_ASAP7_75t_SL g4012 ( 
.A1(n_3617),
.A2(n_621),
.B1(n_619),
.B2(n_620),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3777),
.B(n_622),
.Y(n_4013)
);

AOI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_3344),
.A2(n_623),
.B(n_624),
.Y(n_4014)
);

OAI21x1_ASAP7_75t_L g4015 ( 
.A1(n_3289),
.A2(n_623),
.B(n_624),
.Y(n_4015)
);

INVxp67_ASAP7_75t_SL g4016 ( 
.A(n_3307),
.Y(n_4016)
);

HB1xp67_ASAP7_75t_L g4017 ( 
.A(n_3444),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3438),
.B(n_949),
.Y(n_4018)
);

O2A1O1Ixp33_ASAP7_75t_L g4019 ( 
.A1(n_3632),
.A2(n_627),
.B(n_625),
.C(n_626),
.Y(n_4019)
);

NOR2xp33_ASAP7_75t_L g4020 ( 
.A(n_3685),
.B(n_626),
.Y(n_4020)
);

BUFx2_ASAP7_75t_L g4021 ( 
.A(n_3431),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3674),
.Y(n_4022)
);

NOR2xp33_ASAP7_75t_L g4023 ( 
.A(n_3736),
.B(n_627),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_SL g4024 ( 
.A(n_3602),
.B(n_629),
.Y(n_4024)
);

OAI22xp5_ASAP7_75t_L g4025 ( 
.A1(n_3646),
.A2(n_632),
.B1(n_630),
.B2(n_631),
.Y(n_4025)
);

O2A1O1Ixp33_ASAP7_75t_L g4026 ( 
.A1(n_3653),
.A2(n_632),
.B(n_630),
.C(n_631),
.Y(n_4026)
);

OAI22xp5_ASAP7_75t_L g4027 ( 
.A1(n_3743),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.Y(n_4027)
);

INVx4_ASAP7_75t_L g4028 ( 
.A(n_3743),
.Y(n_4028)
);

INVxp67_ASAP7_75t_L g4029 ( 
.A(n_3612),
.Y(n_4029)
);

AND2x2_ASAP7_75t_L g4030 ( 
.A(n_3683),
.B(n_633),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_SL g4031 ( 
.A(n_3765),
.B(n_634),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3293),
.Y(n_4032)
);

NOR2xp33_ASAP7_75t_L g4033 ( 
.A(n_3661),
.B(n_635),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3659),
.A2(n_642),
.B1(n_636),
.B2(n_638),
.Y(n_4034)
);

AOI21xp5_ASAP7_75t_L g4035 ( 
.A1(n_3374),
.A2(n_636),
.B(n_638),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3728),
.B(n_643),
.Y(n_4036)
);

A2O1A1Ixp33_ASAP7_75t_SL g4037 ( 
.A1(n_3627),
.A2(n_645),
.B(n_643),
.C(n_644),
.Y(n_4037)
);

O2A1O1Ixp33_ASAP7_75t_L g4038 ( 
.A1(n_3750),
.A2(n_646),
.B(n_644),
.C(n_645),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3705),
.B(n_646),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3732),
.B(n_647),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3662),
.B(n_647),
.Y(n_4041)
);

AOI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_3397),
.A2(n_648),
.B(n_649),
.Y(n_4042)
);

OR2x6_ASAP7_75t_SL g4043 ( 
.A(n_3748),
.B(n_3517),
.Y(n_4043)
);

NOR2xp33_ASAP7_75t_L g4044 ( 
.A(n_3778),
.B(n_649),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3630),
.Y(n_4045)
);

AOI21xp5_ASAP7_75t_L g4046 ( 
.A1(n_3402),
.A2(n_651),
.B(n_652),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3634),
.Y(n_4047)
);

NAND2x1p5_ASAP7_75t_L g4048 ( 
.A(n_3662),
.B(n_652),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3637),
.Y(n_4049)
);

INVx4_ASAP7_75t_L g4050 ( 
.A(n_3258),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3642),
.Y(n_4051)
);

AND2x4_ASAP7_75t_L g4052 ( 
.A(n_3612),
.B(n_949),
.Y(n_4052)
);

OR2x6_ASAP7_75t_L g4053 ( 
.A(n_3509),
.B(n_3629),
.Y(n_4053)
);

CKINVDCx5p33_ASAP7_75t_R g4054 ( 
.A(n_3733),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3467),
.B(n_653),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3474),
.B(n_653),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_SL g4057 ( 
.A(n_3701),
.B(n_654),
.Y(n_4057)
);

BUFx6f_ASAP7_75t_L g4058 ( 
.A(n_3307),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3684),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3614),
.B(n_948),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3647),
.Y(n_4061)
);

OAI21x1_ASAP7_75t_L g4062 ( 
.A1(n_3288),
.A2(n_654),
.B(n_655),
.Y(n_4062)
);

A2O1A1Ixp33_ASAP7_75t_L g4063 ( 
.A1(n_3295),
.A2(n_658),
.B(n_655),
.C(n_657),
.Y(n_4063)
);

NOR2xp33_ASAP7_75t_L g4064 ( 
.A(n_3758),
.B(n_658),
.Y(n_4064)
);

O2A1O1Ixp33_ASAP7_75t_L g4065 ( 
.A1(n_3299),
.A2(n_661),
.B(n_659),
.C(n_660),
.Y(n_4065)
);

NAND2x2_ASAP7_75t_L g4066 ( 
.A(n_3738),
.B(n_3251),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_SL g4067 ( 
.A(n_3701),
.B(n_660),
.Y(n_4067)
);

AOI21xp5_ASAP7_75t_L g4068 ( 
.A1(n_3412),
.A2(n_661),
.B(n_662),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3261),
.B(n_662),
.Y(n_4069)
);

OAI21xp5_ASAP7_75t_L g4070 ( 
.A1(n_3757),
.A2(n_3298),
.B(n_3607),
.Y(n_4070)
);

INVx4_ASAP7_75t_L g4071 ( 
.A(n_3734),
.Y(n_4071)
);

AOI21x1_ASAP7_75t_L g4072 ( 
.A1(n_3271),
.A2(n_3477),
.B(n_3428),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3675),
.Y(n_4073)
);

AOI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_3425),
.A2(n_663),
.B(n_664),
.Y(n_4074)
);

OR2x6_ASAP7_75t_SL g4075 ( 
.A(n_3575),
.B(n_664),
.Y(n_4075)
);

OAI22xp5_ASAP7_75t_L g4076 ( 
.A1(n_3682),
.A2(n_668),
.B1(n_666),
.B2(n_667),
.Y(n_4076)
);

AOI21xp5_ASAP7_75t_L g4077 ( 
.A1(n_3471),
.A2(n_667),
.B(n_668),
.Y(n_4077)
);

OR2x6_ASAP7_75t_L g4078 ( 
.A(n_3771),
.B(n_669),
.Y(n_4078)
);

O2A1O1Ixp33_ASAP7_75t_L g4079 ( 
.A1(n_3456),
.A2(n_672),
.B(n_669),
.C(n_670),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3324),
.Y(n_4080)
);

INVx6_ASAP7_75t_L g4081 ( 
.A(n_3338),
.Y(n_4081)
);

CKINVDCx14_ASAP7_75t_R g4082 ( 
.A(n_3771),
.Y(n_4082)
);

INVx1_ASAP7_75t_SL g4083 ( 
.A(n_3550),
.Y(n_4083)
);

INVxp33_ASAP7_75t_L g4084 ( 
.A(n_3387),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_3332),
.Y(n_4085)
);

HB1xp67_ASAP7_75t_L g4086 ( 
.A(n_3357),
.Y(n_4086)
);

CKINVDCx20_ASAP7_75t_R g4087 ( 
.A(n_3300),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3333),
.Y(n_4088)
);

INVx3_ASAP7_75t_L g4089 ( 
.A(n_3734),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3262),
.Y(n_4090)
);

NOR2x1_ASAP7_75t_R g4091 ( 
.A(n_3737),
.B(n_673),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3533),
.B(n_948),
.Y(n_4092)
);

NOR3xp33_ASAP7_75t_L g4093 ( 
.A(n_3593),
.B(n_673),
.C(n_674),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3359),
.B(n_674),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3268),
.B(n_676),
.Y(n_4095)
);

AO32x1_ASAP7_75t_L g4096 ( 
.A1(n_3587),
.A2(n_678),
.A3(n_676),
.B1(n_677),
.B2(n_679),
.Y(n_4096)
);

NOR2xp33_ASAP7_75t_L g4097 ( 
.A(n_3726),
.B(n_3722),
.Y(n_4097)
);

AOI21xp5_ASAP7_75t_L g4098 ( 
.A1(n_3480),
.A2(n_3484),
.B(n_3498),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3335),
.Y(n_4099)
);

AOI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_3556),
.A2(n_3352),
.B(n_3338),
.Y(n_4100)
);

NOR2xp33_ASAP7_75t_L g4101 ( 
.A(n_3381),
.B(n_678),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3338),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3363),
.B(n_3393),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3651),
.B(n_947),
.Y(n_4104)
);

AOI21xp5_ASAP7_75t_L g4105 ( 
.A1(n_3352),
.A2(n_679),
.B(n_680),
.Y(n_4105)
);

AOI21xp5_ASAP7_75t_L g4106 ( 
.A1(n_3352),
.A2(n_681),
.B(n_682),
.Y(n_4106)
);

BUFx12f_ASAP7_75t_L g4107 ( 
.A(n_3527),
.Y(n_4107)
);

NOR2xp33_ASAP7_75t_L g4108 ( 
.A(n_3656),
.B(n_681),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_SL g4109 ( 
.A(n_3737),
.B(n_682),
.Y(n_4109)
);

NOR2xp33_ASAP7_75t_R g4110 ( 
.A(n_3300),
.B(n_684),
.Y(n_4110)
);

OAI22xp5_ASAP7_75t_L g4111 ( 
.A1(n_3741),
.A2(n_686),
.B1(n_684),
.B2(n_685),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3667),
.B(n_946),
.Y(n_4112)
);

INVx5_ASAP7_75t_L g4113 ( 
.A(n_3527),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_3579),
.A2(n_687),
.B(n_688),
.Y(n_4114)
);

OAI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3283),
.A2(n_689),
.B1(n_687),
.B2(n_688),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3325),
.Y(n_4116)
);

NOR2xp33_ASAP7_75t_SL g4117 ( 
.A(n_3548),
.B(n_3768),
.Y(n_4117)
);

A2O1A1Ixp33_ASAP7_75t_L g4118 ( 
.A1(n_3265),
.A2(n_692),
.B(n_690),
.C(n_691),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_3460),
.B(n_690),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3342),
.Y(n_4120)
);

AOI21xp5_ASAP7_75t_L g4121 ( 
.A1(n_3613),
.A2(n_691),
.B(n_692),
.Y(n_4121)
);

NOR2xp33_ASAP7_75t_L g4122 ( 
.A(n_3670),
.B(n_694),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_SL g4123 ( 
.A(n_3408),
.B(n_694),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3358),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_3361),
.Y(n_4125)
);

NOR2xp33_ASAP7_75t_L g4126 ( 
.A(n_3761),
.B(n_695),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3545),
.B(n_695),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3370),
.Y(n_4128)
);

A2O1A1Ixp33_ASAP7_75t_L g4129 ( 
.A1(n_3752),
.A2(n_698),
.B(n_696),
.C(n_697),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_3373),
.Y(n_4130)
);

O2A1O1Ixp33_ASAP7_75t_L g4131 ( 
.A1(n_3492),
.A2(n_698),
.B(n_696),
.C(n_697),
.Y(n_4131)
);

BUFx12f_ASAP7_75t_L g4132 ( 
.A(n_3527),
.Y(n_4132)
);

CKINVDCx8_ASAP7_75t_R g4133 ( 
.A(n_3773),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3385),
.Y(n_4134)
);

INVx3_ASAP7_75t_L g4135 ( 
.A(n_3313),
.Y(n_4135)
);

AOI22xp33_ASAP7_75t_L g4136 ( 
.A1(n_3383),
.A2(n_702),
.B1(n_699),
.B2(n_700),
.Y(n_4136)
);

AOI22xp5_ASAP7_75t_L g4137 ( 
.A1(n_3779),
.A2(n_704),
.B1(n_700),
.B2(n_702),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3372),
.A2(n_704),
.B(n_706),
.Y(n_4138)
);

NOR2xp33_ASAP7_75t_L g4139 ( 
.A(n_3770),
.B(n_706),
.Y(n_4139)
);

AOI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_3382),
.A2(n_707),
.B(n_708),
.Y(n_4140)
);

INVx5_ASAP7_75t_L g4141 ( 
.A(n_3313),
.Y(n_4141)
);

AOI21xp5_ASAP7_75t_L g4142 ( 
.A1(n_3318),
.A2(n_707),
.B(n_708),
.Y(n_4142)
);

BUFx6f_ASAP7_75t_L g4143 ( 
.A(n_4107),
.Y(n_4143)
);

INVx4_ASAP7_75t_L g4144 ( 
.A(n_3879),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3791),
.Y(n_4145)
);

NAND2x1p5_ASAP7_75t_L g4146 ( 
.A(n_3853),
.B(n_3384),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3805),
.Y(n_4147)
);

INVx4_ASAP7_75t_L g4148 ( 
.A(n_3809),
.Y(n_4148)
);

INVx3_ASAP7_75t_SL g4149 ( 
.A(n_3809),
.Y(n_4149)
);

BUFx6f_ASAP7_75t_L g4150 ( 
.A(n_4132),
.Y(n_4150)
);

INVx6_ASAP7_75t_L g4151 ( 
.A(n_3841),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3806),
.B(n_3377),
.Y(n_4152)
);

BUFx6f_ASAP7_75t_L g4153 ( 
.A(n_3820),
.Y(n_4153)
);

INVx5_ASAP7_75t_L g4154 ( 
.A(n_3820),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_3788),
.Y(n_4155)
);

CKINVDCx5p33_ASAP7_75t_R g4156 ( 
.A(n_3929),
.Y(n_4156)
);

BUFx2_ASAP7_75t_L g4157 ( 
.A(n_3891),
.Y(n_4157)
);

BUFx6f_ASAP7_75t_L g4158 ( 
.A(n_3829),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_3886),
.B(n_3590),
.Y(n_4159)
);

BUFx2_ASAP7_75t_L g4160 ( 
.A(n_3974),
.Y(n_4160)
);

INVx2_ASAP7_75t_SL g4161 ( 
.A(n_3894),
.Y(n_4161)
);

BUFx6f_ASAP7_75t_L g4162 ( 
.A(n_3962),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_3790),
.Y(n_4163)
);

AOI22xp33_ASAP7_75t_L g4164 ( 
.A1(n_3795),
.A2(n_3513),
.B1(n_3782),
.B2(n_3596),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_3846),
.Y(n_4165)
);

INVx1_ASAP7_75t_SL g4166 ( 
.A(n_4004),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_3850),
.Y(n_4167)
);

INVx2_ASAP7_75t_L g4168 ( 
.A(n_3937),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_3946),
.B(n_3577),
.Y(n_4169)
);

INVx1_ASAP7_75t_SL g4170 ( 
.A(n_4087),
.Y(n_4170)
);

INVx1_ASAP7_75t_SL g4171 ( 
.A(n_3797),
.Y(n_4171)
);

BUFx3_ASAP7_75t_L g4172 ( 
.A(n_3948),
.Y(n_4172)
);

INVx5_ASAP7_75t_L g4173 ( 
.A(n_3957),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_4030),
.B(n_3594),
.Y(n_4174)
);

AOI22xp33_ASAP7_75t_SL g4175 ( 
.A1(n_3822),
.A2(n_3739),
.B1(n_3365),
.B2(n_3348),
.Y(n_4175)
);

BUFx3_ASAP7_75t_L g4176 ( 
.A(n_3962),
.Y(n_4176)
);

INVx6_ASAP7_75t_L g4177 ( 
.A(n_3892),
.Y(n_4177)
);

INVx3_ASAP7_75t_SL g4178 ( 
.A(n_3881),
.Y(n_4178)
);

BUFx6f_ASAP7_75t_L g4179 ( 
.A(n_3969),
.Y(n_4179)
);

NAND2x1_ASAP7_75t_L g4180 ( 
.A(n_4053),
.B(n_3384),
.Y(n_4180)
);

INVx3_ASAP7_75t_L g4181 ( 
.A(n_3924),
.Y(n_4181)
);

CKINVDCx11_ASAP7_75t_R g4182 ( 
.A(n_3942),
.Y(n_4182)
);

BUFx6f_ASAP7_75t_L g4183 ( 
.A(n_3984),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_3939),
.Y(n_4184)
);

INVxp67_ASAP7_75t_SL g4185 ( 
.A(n_3815),
.Y(n_4185)
);

INVx4_ASAP7_75t_L g4186 ( 
.A(n_4002),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3808),
.Y(n_4187)
);

INVx5_ASAP7_75t_L g4188 ( 
.A(n_4028),
.Y(n_4188)
);

BUFx6f_ASAP7_75t_L g4189 ( 
.A(n_3972),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3810),
.Y(n_4190)
);

BUFx2_ASAP7_75t_L g4191 ( 
.A(n_3862),
.Y(n_4191)
);

INVx4_ASAP7_75t_L g4192 ( 
.A(n_3825),
.Y(n_4192)
);

BUFx12f_ASAP7_75t_L g4193 ( 
.A(n_4054),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3824),
.Y(n_4194)
);

BUFx4_ASAP7_75t_SL g4195 ( 
.A(n_4009),
.Y(n_4195)
);

CKINVDCx5p33_ASAP7_75t_R g4196 ( 
.A(n_3800),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_3855),
.A2(n_3321),
.B1(n_3442),
.B2(n_3264),
.Y(n_4197)
);

INVx3_ASAP7_75t_SL g4198 ( 
.A(n_3826),
.Y(n_4198)
);

INVx4_ASAP7_75t_L g4199 ( 
.A(n_3814),
.Y(n_4199)
);

BUFx3_ASAP7_75t_L g4200 ( 
.A(n_3807),
.Y(n_4200)
);

BUFx12f_ASAP7_75t_L g4201 ( 
.A(n_3931),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_3830),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_3940),
.Y(n_4203)
);

INVx3_ASAP7_75t_L g4204 ( 
.A(n_4071),
.Y(n_4204)
);

BUFx6f_ASAP7_75t_L g4205 ( 
.A(n_3972),
.Y(n_4205)
);

BUFx3_ASAP7_75t_L g4206 ( 
.A(n_3997),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_3951),
.Y(n_4207)
);

AOI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_3920),
.A2(n_3551),
.B1(n_3368),
.B2(n_3763),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3837),
.Y(n_4209)
);

INVxp67_ASAP7_75t_SL g4210 ( 
.A(n_3847),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_4036),
.B(n_3775),
.Y(n_4211)
);

BUFx8_ASAP7_75t_SL g4212 ( 
.A(n_4001),
.Y(n_4212)
);

BUFx4_ASAP7_75t_SL g4213 ( 
.A(n_4078),
.Y(n_4213)
);

BUFx2_ASAP7_75t_L g4214 ( 
.A(n_4021),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4040),
.B(n_3780),
.Y(n_4215)
);

BUFx3_ASAP7_75t_L g4216 ( 
.A(n_3857),
.Y(n_4216)
);

INVx3_ASAP7_75t_L g4217 ( 
.A(n_4050),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3877),
.Y(n_4218)
);

AND2x2_ASAP7_75t_L g4219 ( 
.A(n_3799),
.B(n_3695),
.Y(n_4219)
);

BUFx3_ASAP7_75t_L g4220 ( 
.A(n_4005),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3955),
.Y(n_4221)
);

INVx2_ASAP7_75t_SL g4222 ( 
.A(n_3859),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3882),
.Y(n_4223)
);

HB1xp67_ASAP7_75t_L g4224 ( 
.A(n_3856),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3890),
.Y(n_4225)
);

BUFx2_ASAP7_75t_R g4226 ( 
.A(n_3987),
.Y(n_4226)
);

INVx3_ASAP7_75t_L g4227 ( 
.A(n_3817),
.Y(n_4227)
);

BUFx6f_ASAP7_75t_L g4228 ( 
.A(n_3895),
.Y(n_4228)
);

INVx3_ASAP7_75t_L g4229 ( 
.A(n_4000),
.Y(n_4229)
);

INVx8_ASAP7_75t_L g4230 ( 
.A(n_4078),
.Y(n_4230)
);

AND2x4_ASAP7_75t_L g4231 ( 
.A(n_3848),
.B(n_3409),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_3811),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4103),
.B(n_3725),
.Y(n_4233)
);

INVx1_ASAP7_75t_SL g4234 ( 
.A(n_3852),
.Y(n_4234)
);

BUFx3_ASAP7_75t_L g4235 ( 
.A(n_3988),
.Y(n_4235)
);

INVxp67_ASAP7_75t_SL g4236 ( 
.A(n_3973),
.Y(n_4236)
);

INVx8_ASAP7_75t_L g4237 ( 
.A(n_4053),
.Y(n_4237)
);

BUFx24_ASAP7_75t_SL g4238 ( 
.A(n_3839),
.Y(n_4238)
);

INVx3_ASAP7_75t_L g4239 ( 
.A(n_4089),
.Y(n_4239)
);

INVx3_ASAP7_75t_L g4240 ( 
.A(n_4048),
.Y(n_4240)
);

INVx3_ASAP7_75t_SL g4241 ( 
.A(n_4052),
.Y(n_4241)
);

INVx5_ASAP7_75t_L g4242 ( 
.A(n_3895),
.Y(n_4242)
);

BUFx2_ASAP7_75t_R g4243 ( 
.A(n_4075),
.Y(n_4243)
);

BUFx10_ASAP7_75t_L g4244 ( 
.A(n_3975),
.Y(n_4244)
);

INVx4_ASAP7_75t_L g4245 ( 
.A(n_4113),
.Y(n_4245)
);

BUFx3_ASAP7_75t_L g4246 ( 
.A(n_4113),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3905),
.Y(n_4247)
);

BUFx6f_ASAP7_75t_L g4248 ( 
.A(n_3902),
.Y(n_4248)
);

INVx1_ASAP7_75t_SL g4249 ( 
.A(n_4083),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_3906),
.Y(n_4250)
);

NOR2xp33_ASAP7_75t_L g4251 ( 
.A(n_3832),
.B(n_3687),
.Y(n_4251)
);

BUFx3_ASAP7_75t_L g4252 ( 
.A(n_4113),
.Y(n_4252)
);

CKINVDCx11_ASAP7_75t_R g4253 ( 
.A(n_4133),
.Y(n_4253)
);

INVxp33_ASAP7_75t_L g4254 ( 
.A(n_4091),
.Y(n_4254)
);

INVx3_ASAP7_75t_SL g4255 ( 
.A(n_3973),
.Y(n_4255)
);

INVx1_ASAP7_75t_SL g4256 ( 
.A(n_3812),
.Y(n_4256)
);

BUFx3_ASAP7_75t_L g4257 ( 
.A(n_3902),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_3793),
.B(n_3411),
.Y(n_4258)
);

BUFx3_ASAP7_75t_L g4259 ( 
.A(n_3949),
.Y(n_4259)
);

INVx3_ASAP7_75t_L g4260 ( 
.A(n_4141),
.Y(n_4260)
);

BUFx12f_ASAP7_75t_L g4261 ( 
.A(n_3899),
.Y(n_4261)
);

BUFx4_ASAP7_75t_SL g4262 ( 
.A(n_3834),
.Y(n_4262)
);

INVx2_ASAP7_75t_R g4263 ( 
.A(n_4141),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_4082),
.B(n_709),
.Y(n_4264)
);

BUFx12f_ASAP7_75t_L g4265 ( 
.A(n_3949),
.Y(n_4265)
);

INVx6_ASAP7_75t_SL g4266 ( 
.A(n_3813),
.Y(n_4266)
);

BUFx8_ASAP7_75t_L g4267 ( 
.A(n_4119),
.Y(n_4267)
);

INVx8_ASAP7_75t_L g4268 ( 
.A(n_4141),
.Y(n_4268)
);

INVx4_ASAP7_75t_L g4269 ( 
.A(n_3973),
.Y(n_4269)
);

INVx1_ASAP7_75t_SL g4270 ( 
.A(n_4110),
.Y(n_4270)
);

INVx6_ASAP7_75t_L g4271 ( 
.A(n_3973),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_3903),
.B(n_709),
.Y(n_4272)
);

BUFx24_ASAP7_75t_L g4273 ( 
.A(n_3884),
.Y(n_4273)
);

INVx2_ASAP7_75t_SL g4274 ( 
.A(n_3971),
.Y(n_4274)
);

INVx2_ASAP7_75t_L g4275 ( 
.A(n_3861),
.Y(n_4275)
);

INVx1_ASAP7_75t_SL g4276 ( 
.A(n_3872),
.Y(n_4276)
);

INVx1_ASAP7_75t_SL g4277 ( 
.A(n_4081),
.Y(n_4277)
);

INVx3_ASAP7_75t_L g4278 ( 
.A(n_4135),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3953),
.B(n_3413),
.Y(n_4279)
);

BUFx2_ASAP7_75t_SL g4280 ( 
.A(n_3823),
.Y(n_4280)
);

BUFx3_ASAP7_75t_L g4281 ( 
.A(n_4081),
.Y(n_4281)
);

INVx4_ASAP7_75t_L g4282 ( 
.A(n_4058),
.Y(n_4282)
);

INVx3_ASAP7_75t_SL g4283 ( 
.A(n_4012),
.Y(n_4283)
);

NAND2x1p5_ASAP7_75t_L g4284 ( 
.A(n_3927),
.B(n_3409),
.Y(n_4284)
);

BUFx3_ASAP7_75t_L g4285 ( 
.A(n_3926),
.Y(n_4285)
);

CKINVDCx5p33_ASAP7_75t_R g4286 ( 
.A(n_3871),
.Y(n_4286)
);

CKINVDCx20_ASAP7_75t_R g4287 ( 
.A(n_3952),
.Y(n_4287)
);

BUFx3_ASAP7_75t_L g4288 ( 
.A(n_3941),
.Y(n_4288)
);

BUFx6f_ASAP7_75t_L g4289 ( 
.A(n_4058),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_3916),
.Y(n_4290)
);

INVx2_ASAP7_75t_L g4291 ( 
.A(n_3901),
.Y(n_4291)
);

NAND2x1p5_ASAP7_75t_L g4292 ( 
.A(n_3802),
.B(n_3585),
.Y(n_4292)
);

INVxp67_ASAP7_75t_L g4293 ( 
.A(n_3860),
.Y(n_4293)
);

CKINVDCx14_ASAP7_75t_R g4294 ( 
.A(n_3836),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_3967),
.B(n_3977),
.Y(n_4295)
);

BUFx6f_ASAP7_75t_L g4296 ( 
.A(n_4102),
.Y(n_4296)
);

CKINVDCx6p67_ASAP7_75t_R g4297 ( 
.A(n_3979),
.Y(n_4297)
);

AND2x2_ASAP7_75t_L g4298 ( 
.A(n_3863),
.B(n_710),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_3918),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_3914),
.Y(n_4300)
);

INVx1_ASAP7_75t_SL g4301 ( 
.A(n_3827),
.Y(n_4301)
);

BUFx6f_ASAP7_75t_L g4302 ( 
.A(n_3842),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_3867),
.Y(n_4303)
);

AND2x2_ASAP7_75t_L g4304 ( 
.A(n_4094),
.B(n_710),
.Y(n_4304)
);

BUFx6f_ASAP7_75t_L g4305 ( 
.A(n_3873),
.Y(n_4305)
);

INVx6_ASAP7_75t_L g4306 ( 
.A(n_3990),
.Y(n_4306)
);

INVx3_ASAP7_75t_L g4307 ( 
.A(n_4022),
.Y(n_4307)
);

OAI22xp5_ASAP7_75t_L g4308 ( 
.A1(n_3843),
.A2(n_3660),
.B1(n_3557),
.B2(n_3628),
.Y(n_4308)
);

BUFx4_ASAP7_75t_SL g4309 ( 
.A(n_3993),
.Y(n_4309)
);

BUFx6f_ASAP7_75t_L g4310 ( 
.A(n_4059),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_L g4311 ( 
.A(n_3963),
.B(n_3330),
.Y(n_4311)
);

BUFx2_ASAP7_75t_SL g4312 ( 
.A(n_3915),
.Y(n_4312)
);

INVx5_ASAP7_75t_L g4313 ( 
.A(n_3990),
.Y(n_4313)
);

CKINVDCx14_ASAP7_75t_R g4314 ( 
.A(n_3961),
.Y(n_4314)
);

INVx8_ASAP7_75t_L g4315 ( 
.A(n_3990),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3900),
.Y(n_4316)
);

INVx5_ASAP7_75t_SL g4317 ( 
.A(n_3844),
.Y(n_4317)
);

HB1xp67_ASAP7_75t_L g4318 ( 
.A(n_3986),
.Y(n_4318)
);

NAND2x1p5_ASAP7_75t_L g4319 ( 
.A(n_4041),
.B(n_3522),
.Y(n_4319)
);

INVx2_ASAP7_75t_SL g4320 ( 
.A(n_3989),
.Y(n_4320)
);

INVx5_ASAP7_75t_L g4321 ( 
.A(n_4127),
.Y(n_4321)
);

BUFx2_ASAP7_75t_L g4322 ( 
.A(n_4029),
.Y(n_4322)
);

INVx6_ASAP7_75t_SL g4323 ( 
.A(n_3785),
.Y(n_4323)
);

CKINVDCx5p33_ASAP7_75t_R g4324 ( 
.A(n_4008),
.Y(n_4324)
);

BUFx6f_ASAP7_75t_L g4325 ( 
.A(n_3980),
.Y(n_4325)
);

INVx3_ASAP7_75t_SL g4326 ( 
.A(n_4057),
.Y(n_4326)
);

NAND2x1p5_ASAP7_75t_L g4327 ( 
.A(n_4067),
.B(n_3386),
.Y(n_4327)
);

BUFx8_ASAP7_75t_SL g4328 ( 
.A(n_3854),
.Y(n_4328)
);

BUFx2_ASAP7_75t_L g4329 ( 
.A(n_4016),
.Y(n_4329)
);

BUFx3_ASAP7_75t_L g4330 ( 
.A(n_3866),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_3796),
.Y(n_4331)
);

AND2x4_ASAP7_75t_L g4332 ( 
.A(n_3821),
.B(n_3652),
.Y(n_4332)
);

BUFx6f_ASAP7_75t_L g4333 ( 
.A(n_3864),
.Y(n_4333)
);

BUFx5_ASAP7_75t_L g4334 ( 
.A(n_3994),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_3840),
.Y(n_4335)
);

INVx3_ASAP7_75t_SL g4336 ( 
.A(n_4109),
.Y(n_4336)
);

OR2x6_ASAP7_75t_L g4337 ( 
.A(n_3831),
.B(n_3784),
.Y(n_4337)
);

BUFx4_ASAP7_75t_SL g4338 ( 
.A(n_3996),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_3840),
.Y(n_4339)
);

AOI22xp33_ASAP7_75t_L g4340 ( 
.A1(n_4093),
.A2(n_3270),
.B1(n_3718),
.B2(n_3366),
.Y(n_4340)
);

INVx8_ASAP7_75t_L g4341 ( 
.A(n_4084),
.Y(n_4341)
);

INVx3_ASAP7_75t_L g4342 ( 
.A(n_3819),
.Y(n_4342)
);

NAND2x1p5_ASAP7_75t_L g4343 ( 
.A(n_3913),
.B(n_3421),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4086),
.B(n_711),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_4007),
.B(n_3416),
.Y(n_4345)
);

INVx1_ASAP7_75t_SL g4346 ( 
.A(n_4017),
.Y(n_4346)
);

INVx5_ASAP7_75t_L g4347 ( 
.A(n_4125),
.Y(n_4347)
);

BUFx3_ASAP7_75t_L g4348 ( 
.A(n_3934),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_L g4349 ( 
.A(n_4032),
.B(n_3426),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4010),
.B(n_713),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_3880),
.Y(n_4351)
);

INVx3_ASAP7_75t_L g4352 ( 
.A(n_4015),
.Y(n_4352)
);

CKINVDCx5p33_ASAP7_75t_R g4353 ( 
.A(n_3959),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3883),
.Y(n_4354)
);

INVx5_ASAP7_75t_L g4355 ( 
.A(n_4128),
.Y(n_4355)
);

INVx2_ASAP7_75t_SL g4356 ( 
.A(n_4060),
.Y(n_4356)
);

HB1xp67_ASAP7_75t_L g4357 ( 
.A(n_3982),
.Y(n_4357)
);

CKINVDCx11_ASAP7_75t_R g4358 ( 
.A(n_4043),
.Y(n_4358)
);

INVx2_ASAP7_75t_SL g4359 ( 
.A(n_4011),
.Y(n_4359)
);

BUFx10_ASAP7_75t_L g4360 ( 
.A(n_4020),
.Y(n_4360)
);

INVx3_ASAP7_75t_L g4361 ( 
.A(n_4130),
.Y(n_4361)
);

INVx1_ASAP7_75t_SL g4362 ( 
.A(n_3908),
.Y(n_4362)
);

BUFx3_ASAP7_75t_L g4363 ( 
.A(n_3925),
.Y(n_4363)
);

INVx1_ASAP7_75t_SL g4364 ( 
.A(n_3922),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_3887),
.Y(n_4365)
);

AOI22xp33_ASAP7_75t_L g4366 ( 
.A1(n_3911),
.A2(n_3673),
.B1(n_3415),
.B2(n_3269),
.Y(n_4366)
);

INVx3_ASAP7_75t_L g4367 ( 
.A(n_3933),
.Y(n_4367)
);

BUFx3_ASAP7_75t_L g4368 ( 
.A(n_3858),
.Y(n_4368)
);

BUFx6f_ASAP7_75t_L g4369 ( 
.A(n_3999),
.Y(n_4369)
);

BUFx6f_ASAP7_75t_L g4370 ( 
.A(n_4013),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4062),
.Y(n_4371)
);

INVx2_ASAP7_75t_SL g4372 ( 
.A(n_4025),
.Y(n_4372)
);

BUFx4_ASAP7_75t_SL g4373 ( 
.A(n_4045),
.Y(n_4373)
);

INVxp67_ASAP7_75t_SL g4374 ( 
.A(n_3787),
.Y(n_4374)
);

BUFx6f_ASAP7_75t_L g4375 ( 
.A(n_4092),
.Y(n_4375)
);

BUFx12f_ASAP7_75t_L g4376 ( 
.A(n_4027),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4047),
.Y(n_4377)
);

NOR2xp33_ASAP7_75t_L g4378 ( 
.A(n_3970),
.B(n_3681),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_4049),
.Y(n_4379)
);

INVxp67_ASAP7_75t_SL g4380 ( 
.A(n_3792),
.Y(n_4380)
);

INVx3_ASAP7_75t_L g4381 ( 
.A(n_3893),
.Y(n_4381)
);

INVx3_ASAP7_75t_L g4382 ( 
.A(n_3896),
.Y(n_4382)
);

NAND2x1p5_ASAP7_75t_L g4383 ( 
.A(n_3945),
.B(n_3769),
.Y(n_4383)
);

INVx3_ASAP7_75t_L g4384 ( 
.A(n_4148),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4155),
.Y(n_4385)
);

OAI21x1_ASAP7_75t_SL g4386 ( 
.A1(n_4274),
.A2(n_3803),
.B(n_3816),
.Y(n_4386)
);

OAI21x1_ASAP7_75t_L g4387 ( 
.A1(n_4352),
.A2(n_4072),
.B(n_4100),
.Y(n_4387)
);

OAI21x1_ASAP7_75t_L g4388 ( 
.A1(n_4342),
.A2(n_4116),
.B(n_3981),
.Y(n_4388)
);

NOR2xp33_ASAP7_75t_L g4389 ( 
.A(n_4254),
.B(n_3932),
.Y(n_4389)
);

AND2x4_ASAP7_75t_L g4390 ( 
.A(n_4157),
.B(n_3828),
.Y(n_4390)
);

OA21x2_ASAP7_75t_L g4391 ( 
.A1(n_4374),
.A2(n_3798),
.B(n_3818),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_4163),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4232),
.B(n_4051),
.Y(n_4393)
);

INVx3_ASAP7_75t_L g4394 ( 
.A(n_4179),
.Y(n_4394)
);

OAI21xp5_ASAP7_75t_L g4395 ( 
.A1(n_4378),
.A2(n_3935),
.B(n_3804),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4145),
.Y(n_4396)
);

OAI22xp5_ASAP7_75t_L g4397 ( 
.A1(n_4243),
.A2(n_3930),
.B1(n_3910),
.B2(n_3912),
.Y(n_4397)
);

AND2x4_ASAP7_75t_L g4398 ( 
.A(n_4160),
.B(n_4191),
.Y(n_4398)
);

OAI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_4175),
.A2(n_3868),
.B(n_3874),
.Y(n_4399)
);

A2O1A1Ixp33_ASAP7_75t_L g4400 ( 
.A1(n_4315),
.A2(n_3865),
.B(n_3950),
.C(n_3876),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4147),
.Y(n_4401)
);

OAI21x1_ASAP7_75t_SL g4402 ( 
.A1(n_4269),
.A2(n_3851),
.B(n_3845),
.Y(n_4402)
);

AOI22xp33_ASAP7_75t_L g4403 ( 
.A1(n_4376),
.A2(n_4039),
.B1(n_4031),
.B2(n_4024),
.Y(n_4403)
);

INVx2_ASAP7_75t_L g4404 ( 
.A(n_4165),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4187),
.Y(n_4405)
);

HB1xp67_ASAP7_75t_L g4406 ( 
.A(n_4288),
.Y(n_4406)
);

INVx2_ASAP7_75t_SL g4407 ( 
.A(n_4179),
.Y(n_4407)
);

NOR2xp67_ASAP7_75t_L g4408 ( 
.A(n_4188),
.B(n_3833),
.Y(n_4408)
);

BUFx2_ASAP7_75t_SL g4409 ( 
.A(n_4144),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_4285),
.B(n_4061),
.Y(n_4410)
);

NOR3xp33_ASAP7_75t_L g4411 ( 
.A(n_4251),
.B(n_3801),
.C(n_3789),
.Y(n_4411)
);

OAI21x1_ASAP7_75t_L g4412 ( 
.A1(n_4371),
.A2(n_3978),
.B(n_3869),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4190),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_4301),
.B(n_4073),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4194),
.Y(n_4415)
);

OR2x2_ASAP7_75t_L g4416 ( 
.A(n_4210),
.B(n_4080),
.Y(n_4416)
);

HB1xp67_ASAP7_75t_L g4417 ( 
.A(n_4318),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_L g4418 ( 
.A(n_4377),
.B(n_4085),
.Y(n_4418)
);

AOI22xp33_ASAP7_75t_L g4419 ( 
.A1(n_4368),
.A2(n_4332),
.B1(n_4321),
.B2(n_4317),
.Y(n_4419)
);

O2A1O1Ixp33_ASAP7_75t_L g4420 ( 
.A1(n_4381),
.A2(n_3870),
.B(n_3794),
.C(n_4018),
.Y(n_4420)
);

NAND2x1p5_ASAP7_75t_L g4421 ( 
.A(n_4173),
.B(n_3947),
.Y(n_4421)
);

INVx2_ASAP7_75t_L g4422 ( 
.A(n_4167),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4202),
.Y(n_4423)
);

OAI21x1_ASAP7_75t_L g4424 ( 
.A1(n_4180),
.A2(n_3838),
.B(n_3835),
.Y(n_4424)
);

AND2x4_ASAP7_75t_L g4425 ( 
.A(n_4166),
.B(n_4088),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_4209),
.Y(n_4426)
);

OAI21x1_ASAP7_75t_L g4427 ( 
.A1(n_4339),
.A2(n_3849),
.B(n_3960),
.Y(n_4427)
);

OAI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_4340),
.A2(n_3729),
.B(n_3717),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_4218),
.Y(n_4429)
);

AOI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_4236),
.A2(n_4098),
.B(n_4123),
.Y(n_4430)
);

NOR2xp33_ASAP7_75t_L g4431 ( 
.A(n_4328),
.B(n_4097),
.Y(n_4431)
);

OR2x2_ASAP7_75t_L g4432 ( 
.A(n_4185),
.B(n_4224),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4223),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4379),
.B(n_4099),
.Y(n_4434)
);

A2O1A1Ixp33_ASAP7_75t_L g4435 ( 
.A1(n_4237),
.A2(n_3786),
.B(n_3958),
.C(n_3936),
.Y(n_4435)
);

OAI22xp5_ASAP7_75t_L g4436 ( 
.A1(n_4283),
.A2(n_4118),
.B1(n_4129),
.B2(n_3897),
.Y(n_4436)
);

BUFx3_ASAP7_75t_L g4437 ( 
.A(n_4149),
.Y(n_4437)
);

AOI21xp5_ASAP7_75t_L g4438 ( 
.A1(n_4380),
.A2(n_4090),
.B(n_4037),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4225),
.Y(n_4439)
);

OAI21xp5_ASAP7_75t_L g4440 ( 
.A1(n_4208),
.A2(n_3898),
.B(n_3875),
.Y(n_4440)
);

CKINVDCx5p33_ASAP7_75t_R g4441 ( 
.A(n_4262),
.Y(n_4441)
);

OAI21x1_ASAP7_75t_L g4442 ( 
.A1(n_4335),
.A2(n_3878),
.B(n_3907),
.Y(n_4442)
);

A2O1A1Ixp33_ASAP7_75t_L g4443 ( 
.A1(n_4230),
.A2(n_3976),
.B(n_3992),
.C(n_3965),
.Y(n_4443)
);

OAI21x1_ASAP7_75t_L g4444 ( 
.A1(n_4383),
.A2(n_3919),
.B(n_4070),
.Y(n_4444)
);

INVx3_ASAP7_75t_SL g4445 ( 
.A(n_4151),
.Y(n_4445)
);

OAI21x1_ASAP7_75t_L g4446 ( 
.A1(n_4292),
.A2(n_3553),
.B(n_3499),
.Y(n_4446)
);

OAI21x1_ASAP7_75t_L g4447 ( 
.A1(n_4260),
.A2(n_3314),
.B(n_4140),
.Y(n_4447)
);

OAI21x1_ASAP7_75t_L g4448 ( 
.A1(n_4343),
.A2(n_3626),
.B(n_3391),
.Y(n_4448)
);

OAI21xp5_ASAP7_75t_L g4449 ( 
.A1(n_4164),
.A2(n_3889),
.B(n_4014),
.Y(n_4449)
);

AO21x2_ASAP7_75t_L g4450 ( 
.A1(n_4169),
.A2(n_3904),
.B(n_4035),
.Y(n_4450)
);

NAND3xp33_ASAP7_75t_SL g4451 ( 
.A(n_4270),
.B(n_4117),
.C(n_3968),
.Y(n_4451)
);

O2A1O1Ixp33_ASAP7_75t_SL g4452 ( 
.A1(n_4222),
.A2(n_3665),
.B(n_3921),
.C(n_3917),
.Y(n_4452)
);

NOR2xp33_ASAP7_75t_L g4453 ( 
.A(n_4294),
.B(n_4101),
.Y(n_4453)
);

AND2x4_ASAP7_75t_L g4454 ( 
.A(n_4214),
.B(n_4120),
.Y(n_4454)
);

AND2x4_ASAP7_75t_L g4455 ( 
.A(n_4183),
.B(n_4124),
.Y(n_4455)
);

OAI21x1_ASAP7_75t_L g4456 ( 
.A1(n_4204),
.A2(n_3995),
.B(n_3991),
.Y(n_4456)
);

OAI21x1_ASAP7_75t_L g4457 ( 
.A1(n_4361),
.A2(n_4006),
.B(n_4138),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4276),
.B(n_4134),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4320),
.B(n_3888),
.Y(n_4459)
);

OAI22xp33_ASAP7_75t_L g4460 ( 
.A1(n_4321),
.A2(n_4111),
.B1(n_4137),
.B2(n_4066),
.Y(n_4460)
);

OAI21xp5_ASAP7_75t_L g4461 ( 
.A1(n_4152),
.A2(n_4046),
.B(n_4042),
.Y(n_4461)
);

OAI21x1_ASAP7_75t_L g4462 ( 
.A1(n_4319),
.A2(n_3943),
.B(n_4114),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4247),
.Y(n_4463)
);

AOI221xp5_ASAP7_75t_L g4464 ( 
.A1(n_4357),
.A2(n_4064),
.B1(n_4108),
.B2(n_4122),
.C(n_4126),
.Y(n_4464)
);

OAI21x1_ASAP7_75t_L g4465 ( 
.A1(n_4275),
.A2(n_4074),
.B(n_4068),
.Y(n_4465)
);

NOR2xp33_ASAP7_75t_L g4466 ( 
.A(n_4170),
.B(n_3966),
.Y(n_4466)
);

OAI21x1_ASAP7_75t_L g4467 ( 
.A1(n_4291),
.A2(n_4121),
.B(n_4077),
.Y(n_4467)
);

CKINVDCx5p33_ASAP7_75t_R g4468 ( 
.A(n_4182),
.Y(n_4468)
);

HB1xp67_ASAP7_75t_L g4469 ( 
.A(n_4329),
.Y(n_4469)
);

CKINVDCx5p33_ASAP7_75t_R g4470 ( 
.A(n_4156),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4316),
.B(n_3998),
.Y(n_4471)
);

BUFx2_ASAP7_75t_L g4472 ( 
.A(n_4323),
.Y(n_4472)
);

BUFx4f_ASAP7_75t_SL g4473 ( 
.A(n_4193),
.Y(n_4473)
);

BUFx2_ASAP7_75t_SL g4474 ( 
.A(n_4173),
.Y(n_4474)
);

NOR2x1_ASAP7_75t_SL g4475 ( 
.A(n_4313),
.B(n_3909),
.Y(n_4475)
);

AOI22xp33_ASAP7_75t_L g4476 ( 
.A1(n_4359),
.A2(n_4372),
.B1(n_4358),
.B2(n_4308),
.Y(n_4476)
);

NOR3xp33_ASAP7_75t_L g4477 ( 
.A(n_4382),
.B(n_4311),
.C(n_4240),
.Y(n_4477)
);

AOI21xp5_ASAP7_75t_L g4478 ( 
.A1(n_4337),
.A2(n_3885),
.B(n_4079),
.Y(n_4478)
);

OA21x2_ASAP7_75t_L g4479 ( 
.A1(n_4258),
.A2(n_3640),
.B(n_3983),
.Y(n_4479)
);

OAI21x1_ASAP7_75t_L g4480 ( 
.A1(n_4168),
.A2(n_4142),
.B(n_4106),
.Y(n_4480)
);

OAI21x1_ASAP7_75t_L g4481 ( 
.A1(n_4184),
.A2(n_4207),
.B(n_4203),
.Y(n_4481)
);

OR2x2_ASAP7_75t_L g4482 ( 
.A(n_4312),
.B(n_4346),
.Y(n_4482)
);

INVx2_ASAP7_75t_L g4483 ( 
.A(n_4221),
.Y(n_4483)
);

HB1xp67_ASAP7_75t_L g4484 ( 
.A(n_4310),
.Y(n_4484)
);

BUFx2_ASAP7_75t_L g4485 ( 
.A(n_4334),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_4307),
.Y(n_4486)
);

OAI21x1_ASAP7_75t_L g4487 ( 
.A1(n_4229),
.A2(n_4105),
.B(n_3954),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_4310),
.Y(n_4488)
);

AOI221xp5_ASAP7_75t_L g4489 ( 
.A1(n_4351),
.A2(n_4139),
.B1(n_4023),
.B2(n_3519),
.C(n_3536),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4250),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_4300),
.Y(n_4491)
);

AND2x4_ASAP7_75t_L g4492 ( 
.A(n_4183),
.B(n_3956),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4290),
.Y(n_4493)
);

OAI21x1_ASAP7_75t_L g4494 ( 
.A1(n_4327),
.A2(n_3944),
.B(n_3672),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4299),
.Y(n_4495)
);

OAI21x1_ASAP7_75t_L g4496 ( 
.A1(n_4284),
.A2(n_4217),
.B(n_4181),
.Y(n_4496)
);

OAI21x1_ASAP7_75t_L g4497 ( 
.A1(n_4278),
.A2(n_4197),
.B(n_4295),
.Y(n_4497)
);

INVx2_ASAP7_75t_SL g4498 ( 
.A(n_4309),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4322),
.Y(n_4499)
);

CKINVDCx5p33_ASAP7_75t_R g4500 ( 
.A(n_4195),
.Y(n_4500)
);

OAI21x1_ASAP7_75t_L g4501 ( 
.A1(n_4227),
.A2(n_4367),
.B(n_3678),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4331),
.Y(n_4502)
);

AOI221xp5_ASAP7_75t_L g4503 ( 
.A1(n_4354),
.A2(n_3504),
.B1(n_4115),
.B2(n_4033),
.C(n_4044),
.Y(n_4503)
);

BUFx3_ASAP7_75t_L g4504 ( 
.A(n_4143),
.Y(n_4504)
);

HB1xp67_ASAP7_75t_L g4505 ( 
.A(n_4347),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4334),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4334),
.Y(n_4507)
);

HB1xp67_ASAP7_75t_L g4508 ( 
.A(n_4347),
.Y(n_4508)
);

OAI21x1_ASAP7_75t_L g4509 ( 
.A1(n_4279),
.A2(n_3686),
.B(n_3669),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4355),
.Y(n_4510)
);

OAI22xp5_ASAP7_75t_L g4511 ( 
.A1(n_4306),
.A2(n_4136),
.B1(n_4069),
.B2(n_3490),
.Y(n_4511)
);

OAI21x1_ASAP7_75t_L g4512 ( 
.A1(n_4345),
.A2(n_3435),
.B(n_4131),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_4234),
.B(n_4104),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4355),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4365),
.Y(n_4515)
);

AO31x2_ASAP7_75t_L g4516 ( 
.A1(n_4238),
.A2(n_4003),
.A3(n_4063),
.B(n_3591),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4219),
.B(n_4112),
.Y(n_4517)
);

AND2x4_ASAP7_75t_L g4518 ( 
.A(n_4186),
.B(n_3964),
.Y(n_4518)
);

OAI21x1_ASAP7_75t_L g4519 ( 
.A1(n_4349),
.A2(n_3320),
.B(n_3317),
.Y(n_4519)
);

AND2x6_ASAP7_75t_L g4520 ( 
.A(n_4256),
.B(n_4095),
.Y(n_4520)
);

INVxp67_ASAP7_75t_SL g4521 ( 
.A(n_4296),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4233),
.B(n_713),
.Y(n_4522)
);

AOI22xp33_ASAP7_75t_L g4523 ( 
.A1(n_4375),
.A2(n_4076),
.B1(n_4034),
.B2(n_3928),
.Y(n_4523)
);

OAI21x1_ASAP7_75t_L g4524 ( 
.A1(n_4366),
.A2(n_3326),
.B(n_3322),
.Y(n_4524)
);

OAI21x1_ASAP7_75t_L g4525 ( 
.A1(n_4239),
.A2(n_3329),
.B(n_3327),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_4159),
.B(n_4055),
.Y(n_4526)
);

OR2x6_ASAP7_75t_L g4527 ( 
.A(n_4268),
.B(n_4261),
.Y(n_4527)
);

CKINVDCx6p67_ASAP7_75t_R g4528 ( 
.A(n_4273),
.Y(n_4528)
);

INVx2_ASAP7_75t_L g4529 ( 
.A(n_4296),
.Y(n_4529)
);

INVxp67_ASAP7_75t_L g4530 ( 
.A(n_4220),
.Y(n_4530)
);

AOI22xp5_ASAP7_75t_L g4531 ( 
.A1(n_4353),
.A2(n_4056),
.B1(n_3543),
.B2(n_3938),
.Y(n_4531)
);

OAI21x1_ASAP7_75t_L g4532 ( 
.A1(n_4146),
.A2(n_3343),
.B(n_3339),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4189),
.Y(n_4533)
);

OAI21x1_ASAP7_75t_L g4534 ( 
.A1(n_4263),
.A2(n_3350),
.B(n_3345),
.Y(n_4534)
);

BUFx6f_ASAP7_75t_L g4535 ( 
.A(n_4143),
.Y(n_4535)
);

OAI21x1_ASAP7_75t_L g4536 ( 
.A1(n_4298),
.A2(n_3353),
.B(n_3351),
.Y(n_4536)
);

INVx1_ASAP7_75t_SL g4537 ( 
.A(n_4338),
.Y(n_4537)
);

OR2x2_ASAP7_75t_L g4538 ( 
.A(n_4330),
.B(n_3447),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4189),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4344),
.Y(n_4540)
);

OAI21xp5_ASAP7_75t_L g4541 ( 
.A1(n_4350),
.A2(n_3774),
.B(n_4065),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4375),
.Y(n_4542)
);

AO21x2_ASAP7_75t_L g4543 ( 
.A1(n_4272),
.A2(n_3985),
.B(n_3690),
.Y(n_4543)
);

AO21x2_ASAP7_75t_L g4544 ( 
.A1(n_4231),
.A2(n_3497),
.B(n_3496),
.Y(n_4544)
);

INVxp67_ASAP7_75t_L g4545 ( 
.A(n_4348),
.Y(n_4545)
);

AND2x4_ASAP7_75t_L g4546 ( 
.A(n_4313),
.B(n_3454),
.Y(n_4546)
);

OR2x2_ASAP7_75t_L g4547 ( 
.A(n_4198),
.B(n_3458),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4385),
.Y(n_4548)
);

INVx3_ASAP7_75t_L g4549 ( 
.A(n_4398),
.Y(n_4549)
);

INVx3_ASAP7_75t_L g4550 ( 
.A(n_4485),
.Y(n_4550)
);

BUFx6f_ASAP7_75t_L g4551 ( 
.A(n_4496),
.Y(n_4551)
);

INVx2_ASAP7_75t_L g4552 ( 
.A(n_4392),
.Y(n_4552)
);

BUFx2_ASAP7_75t_L g4553 ( 
.A(n_4528),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4404),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4422),
.Y(n_4555)
);

INVx2_ASAP7_75t_SL g4556 ( 
.A(n_4437),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_4483),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4491),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_4481),
.Y(n_4559)
);

AOI22xp33_ASAP7_75t_L g4560 ( 
.A1(n_4411),
.A2(n_4174),
.B1(n_4363),
.B2(n_4314),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_4417),
.Y(n_4561)
);

AO21x2_ASAP7_75t_L g4562 ( 
.A1(n_4386),
.A2(n_4264),
.B(n_4304),
.Y(n_4562)
);

HB1xp67_ASAP7_75t_L g4563 ( 
.A(n_4469),
.Y(n_4563)
);

BUFx3_ASAP7_75t_L g4564 ( 
.A(n_4384),
.Y(n_4564)
);

AOI22xp33_ASAP7_75t_SL g4565 ( 
.A1(n_4406),
.A2(n_4280),
.B1(n_4201),
.B2(n_4267),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4396),
.Y(n_4566)
);

INVx3_ASAP7_75t_L g4567 ( 
.A(n_4485),
.Y(n_4567)
);

AOI22xp33_ASAP7_75t_SL g4568 ( 
.A1(n_4390),
.A2(n_4188),
.B1(n_4216),
.B2(n_4177),
.Y(n_4568)
);

OAI22xp5_ASAP7_75t_L g4569 ( 
.A1(n_4476),
.A2(n_4226),
.B1(n_4336),
.B2(n_4326),
.Y(n_4569)
);

INVx2_ASAP7_75t_SL g4570 ( 
.A(n_4535),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4401),
.Y(n_4571)
);

CKINVDCx11_ASAP7_75t_R g4572 ( 
.A(n_4445),
.Y(n_4572)
);

INVx2_ASAP7_75t_L g4573 ( 
.A(n_4495),
.Y(n_4573)
);

OAI21x1_ASAP7_75t_L g4574 ( 
.A1(n_4387),
.A2(n_3712),
.B(n_3410),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4405),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4413),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_4415),
.Y(n_4577)
);

AND2x2_ASAP7_75t_L g4578 ( 
.A(n_4499),
.B(n_4333),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_4515),
.B(n_4502),
.Y(n_4579)
);

INVx2_ASAP7_75t_L g4580 ( 
.A(n_4423),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4458),
.B(n_4333),
.Y(n_4581)
);

AOI22xp33_ASAP7_75t_L g4582 ( 
.A1(n_4397),
.A2(n_4356),
.B1(n_4370),
.B2(n_4369),
.Y(n_4582)
);

HB1xp67_ASAP7_75t_L g4583 ( 
.A(n_4432),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4426),
.Y(n_4584)
);

NAND2x1_ASAP7_75t_L g4585 ( 
.A(n_4498),
.B(n_4158),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4429),
.Y(n_4586)
);

OAI22xp5_ASAP7_75t_L g4587 ( 
.A1(n_4403),
.A2(n_4178),
.B1(n_4324),
.B2(n_4241),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4433),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4439),
.Y(n_4589)
);

INVx2_ASAP7_75t_L g4590 ( 
.A(n_4463),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4490),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4493),
.Y(n_4592)
);

INVx3_ASAP7_75t_L g4593 ( 
.A(n_4482),
.Y(n_4593)
);

AO21x2_ASAP7_75t_L g4594 ( 
.A1(n_4438),
.A2(n_3510),
.B(n_3507),
.Y(n_4594)
);

OAI21x1_ASAP7_75t_L g4595 ( 
.A1(n_4388),
.A2(n_3414),
.B(n_3407),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4542),
.Y(n_4596)
);

AOI22xp5_ASAP7_75t_L g4597 ( 
.A1(n_4436),
.A2(n_4297),
.B1(n_4287),
.B2(n_4362),
.Y(n_4597)
);

BUFx3_ASAP7_75t_L g4598 ( 
.A(n_4535),
.Y(n_4598)
);

OAI21x1_ASAP7_75t_L g4599 ( 
.A1(n_4424),
.A2(n_3419),
.B(n_3631),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4410),
.B(n_4244),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4486),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4454),
.B(n_4249),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4416),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4418),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4434),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_4484),
.Y(n_4606)
);

INVx2_ASAP7_75t_L g4607 ( 
.A(n_4488),
.Y(n_4607)
);

HB1xp67_ASAP7_75t_L g4608 ( 
.A(n_4505),
.Y(n_4608)
);

OR2x2_ASAP7_75t_L g4609 ( 
.A(n_4414),
.B(n_4171),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4393),
.Y(n_4610)
);

AOI21x1_ASAP7_75t_L g4611 ( 
.A1(n_4472),
.A2(n_4213),
.B(n_4161),
.Y(n_4611)
);

INVx3_ASAP7_75t_L g4612 ( 
.A(n_4506),
.Y(n_4612)
);

BUFx3_ASAP7_75t_L g4613 ( 
.A(n_4504),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4425),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4508),
.Y(n_4615)
);

CKINVDCx5p33_ASAP7_75t_R g4616 ( 
.A(n_4441),
.Y(n_4616)
);

NAND2x1p5_ASAP7_75t_L g4617 ( 
.A(n_4537),
.B(n_4150),
.Y(n_4617)
);

AO21x1_ASAP7_75t_L g4618 ( 
.A1(n_4460),
.A2(n_4395),
.B(n_4510),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4529),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4540),
.B(n_4364),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4545),
.B(n_4293),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4514),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4507),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4533),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4497),
.Y(n_4625)
);

HB1xp67_ASAP7_75t_L g4626 ( 
.A(n_4455),
.Y(n_4626)
);

INVx2_ASAP7_75t_L g4627 ( 
.A(n_4539),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4513),
.Y(n_4628)
);

HB1xp67_ASAP7_75t_L g4629 ( 
.A(n_4521),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4517),
.Y(n_4630)
);

INVx2_ASAP7_75t_L g4631 ( 
.A(n_4391),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4391),
.Y(n_4632)
);

OAI21xp5_ASAP7_75t_L g4633 ( 
.A1(n_4420),
.A2(n_3297),
.B(n_4019),
.Y(n_4633)
);

OAI21x1_ASAP7_75t_L g4634 ( 
.A1(n_4427),
.A2(n_3633),
.B(n_3369),
.Y(n_4634)
);

INVx2_ASAP7_75t_L g4635 ( 
.A(n_4412),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4459),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4394),
.Y(n_4637)
);

INVx1_ASAP7_75t_SL g4638 ( 
.A(n_4474),
.Y(n_4638)
);

HB1xp67_ASAP7_75t_L g4639 ( 
.A(n_4530),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4407),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4402),
.Y(n_4641)
);

BUFx8_ASAP7_75t_L g4642 ( 
.A(n_4472),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4522),
.B(n_4176),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4402),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4408),
.Y(n_4645)
);

HB1xp67_ASAP7_75t_L g4646 ( 
.A(n_4538),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4430),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4501),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4492),
.Y(n_4649)
);

CKINVDCx16_ASAP7_75t_R g4650 ( 
.A(n_4613),
.Y(n_4650)
);

OA21x2_ASAP7_75t_L g4651 ( 
.A1(n_4645),
.A2(n_4399),
.B(n_4444),
.Y(n_4651)
);

BUFx2_ASAP7_75t_L g4652 ( 
.A(n_4629),
.Y(n_4652)
);

CKINVDCx5p33_ASAP7_75t_R g4653 ( 
.A(n_4572),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4566),
.Y(n_4654)
);

INVxp67_ASAP7_75t_L g4655 ( 
.A(n_4608),
.Y(n_4655)
);

NOR2xp33_ASAP7_75t_L g4656 ( 
.A(n_4553),
.B(n_4389),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4571),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4593),
.B(n_4419),
.Y(n_4658)
);

NOR2x1p5_ASAP7_75t_L g4659 ( 
.A(n_4611),
.B(n_4500),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4577),
.Y(n_4660)
);

AOI22xp33_ASAP7_75t_L g4661 ( 
.A1(n_4618),
.A2(n_4451),
.B1(n_4440),
.B2(n_4449),
.Y(n_4661)
);

OAI22xp5_ASAP7_75t_L g4662 ( 
.A1(n_4597),
.A2(n_4400),
.B1(n_4527),
.B2(n_4547),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_4563),
.Y(n_4663)
);

BUFx10_ASAP7_75t_L g4664 ( 
.A(n_4556),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4584),
.Y(n_4665)
);

AND2x2_ASAP7_75t_L g4666 ( 
.A(n_4593),
.B(n_4477),
.Y(n_4666)
);

HB1xp67_ASAP7_75t_L g4667 ( 
.A(n_4583),
.Y(n_4667)
);

AND2x2_ASAP7_75t_L g4668 ( 
.A(n_4549),
.B(n_4466),
.Y(n_4668)
);

HB1xp67_ASAP7_75t_L g4669 ( 
.A(n_4646),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4552),
.Y(n_4670)
);

INVx3_ASAP7_75t_L g4671 ( 
.A(n_4564),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4549),
.B(n_4286),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4586),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4581),
.B(n_4453),
.Y(n_4674)
);

INVx3_ASAP7_75t_L g4675 ( 
.A(n_4585),
.Y(n_4675)
);

CKINVDCx5p33_ASAP7_75t_R g4676 ( 
.A(n_4616),
.Y(n_4676)
);

NAND2xp33_ASAP7_75t_R g4677 ( 
.A(n_4600),
.B(n_4527),
.Y(n_4677)
);

CKINVDCx5p33_ASAP7_75t_R g4678 ( 
.A(n_4642),
.Y(n_4678)
);

NAND2xp5_ASAP7_75t_L g4679 ( 
.A(n_4628),
.B(n_4526),
.Y(n_4679)
);

HB1xp67_ASAP7_75t_L g4680 ( 
.A(n_4626),
.Y(n_4680)
);

AOI22xp33_ASAP7_75t_SL g4681 ( 
.A1(n_4562),
.A2(n_4520),
.B1(n_4409),
.B2(n_4475),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4614),
.B(n_4431),
.Y(n_4682)
);

CKINVDCx5p33_ASAP7_75t_R g4683 ( 
.A(n_4642),
.Y(n_4683)
);

HB1xp67_ASAP7_75t_L g4684 ( 
.A(n_4558),
.Y(n_4684)
);

OR2x6_ASAP7_75t_L g4685 ( 
.A(n_4617),
.B(n_4341),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4557),
.Y(n_4686)
);

NOR2xp33_ASAP7_75t_L g4687 ( 
.A(n_4638),
.B(n_4212),
.Y(n_4687)
);

AND2x2_ASAP7_75t_L g4688 ( 
.A(n_4578),
.B(n_4518),
.Y(n_4688)
);

INVx2_ASAP7_75t_L g4689 ( 
.A(n_4548),
.Y(n_4689)
);

OR2x2_ASAP7_75t_L g4690 ( 
.A(n_4603),
.B(n_4561),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4548),
.Y(n_4691)
);

NOR2xp33_ASAP7_75t_L g4692 ( 
.A(n_4598),
.B(n_4158),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4588),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4589),
.Y(n_4694)
);

AND2x4_ASAP7_75t_L g4695 ( 
.A(n_4649),
.B(n_4206),
.Y(n_4695)
);

AND2x2_ASAP7_75t_L g4696 ( 
.A(n_4602),
.B(n_4520),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4636),
.B(n_4520),
.Y(n_4697)
);

O2A1O1Ixp33_ASAP7_75t_L g4698 ( 
.A1(n_4569),
.A2(n_4443),
.B(n_4452),
.C(n_4435),
.Y(n_4698)
);

NAND3xp33_ASAP7_75t_L g4699 ( 
.A(n_4625),
.B(n_4464),
.C(n_4428),
.Y(n_4699)
);

INVx2_ASAP7_75t_L g4700 ( 
.A(n_4554),
.Y(n_4700)
);

INVx2_ASAP7_75t_L g4701 ( 
.A(n_4554),
.Y(n_4701)
);

CKINVDCx16_ASAP7_75t_R g4702 ( 
.A(n_4643),
.Y(n_4702)
);

AND2x4_ASAP7_75t_L g4703 ( 
.A(n_4606),
.B(n_4235),
.Y(n_4703)
);

NAND2xp33_ASAP7_75t_R g4704 ( 
.A(n_4550),
.B(n_4196),
.Y(n_4704)
);

OR2x2_ASAP7_75t_L g4705 ( 
.A(n_4604),
.B(n_4471),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4575),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4630),
.B(n_4546),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4610),
.B(n_4604),
.Y(n_4708)
);

INVx2_ASAP7_75t_SL g4709 ( 
.A(n_4570),
.Y(n_4709)
);

AND2x2_ASAP7_75t_L g4710 ( 
.A(n_4615),
.B(n_4302),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4576),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4639),
.B(n_4605),
.Y(n_4712)
);

HB1xp67_ASAP7_75t_L g4713 ( 
.A(n_4573),
.Y(n_4713)
);

OR2x6_ASAP7_75t_L g4714 ( 
.A(n_4587),
.B(n_4150),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4580),
.Y(n_4715)
);

AOI22xp33_ASAP7_75t_SL g4716 ( 
.A1(n_4641),
.A2(n_4421),
.B1(n_4360),
.B2(n_4302),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4605),
.B(n_4479),
.Y(n_4717)
);

INVx1_ASAP7_75t_L g4718 ( 
.A(n_4590),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4591),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4601),
.B(n_4172),
.Y(n_4720)
);

INVx2_ASAP7_75t_L g4721 ( 
.A(n_4555),
.Y(n_4721)
);

BUFx6f_ASAP7_75t_L g4722 ( 
.A(n_4637),
.Y(n_4722)
);

AO32x2_ASAP7_75t_L g4723 ( 
.A1(n_4622),
.A2(n_4511),
.A3(n_4282),
.B1(n_4245),
.B2(n_4199),
.Y(n_4723)
);

CKINVDCx5p33_ASAP7_75t_R g4724 ( 
.A(n_4565),
.Y(n_4724)
);

INVx4_ASAP7_75t_L g4725 ( 
.A(n_4640),
.Y(n_4725)
);

OR2x6_ASAP7_75t_L g4726 ( 
.A(n_4551),
.B(n_4373),
.Y(n_4726)
);

OAI21xp5_ASAP7_75t_L g4727 ( 
.A1(n_4560),
.A2(n_4478),
.B(n_4462),
.Y(n_4727)
);

BUFx2_ASAP7_75t_L g4728 ( 
.A(n_4550),
.Y(n_4728)
);

CKINVDCx5p33_ASAP7_75t_R g4729 ( 
.A(n_4621),
.Y(n_4729)
);

AND2x2_ASAP7_75t_L g4730 ( 
.A(n_4609),
.B(n_4162),
.Y(n_4730)
);

OR2x2_ASAP7_75t_L g4731 ( 
.A(n_4592),
.B(n_4479),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4579),
.Y(n_4732)
);

INVx2_ASAP7_75t_SL g4733 ( 
.A(n_4650),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4688),
.B(n_4652),
.Y(n_4734)
);

INVx2_ASAP7_75t_L g4735 ( 
.A(n_4652),
.Y(n_4735)
);

BUFx6f_ASAP7_75t_L g4736 ( 
.A(n_4653),
.Y(n_4736)
);

NOR4xp25_ASAP7_75t_SL g4737 ( 
.A(n_4677),
.B(n_4468),
.C(n_4645),
.D(n_4470),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_4669),
.Y(n_4738)
);

AOI221xp5_ASAP7_75t_L g4739 ( 
.A1(n_4698),
.A2(n_4582),
.B1(n_4620),
.B2(n_4633),
.C(n_4596),
.Y(n_4739)
);

AND2x2_ASAP7_75t_L g4740 ( 
.A(n_4696),
.B(n_4567),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4717),
.B(n_4732),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4658),
.B(n_4666),
.Y(n_4742)
);

HB1xp67_ASAP7_75t_L g4743 ( 
.A(n_4667),
.Y(n_4743)
);

NOR2xp67_ASAP7_75t_SL g4744 ( 
.A(n_4671),
.B(n_4675),
.Y(n_4744)
);

INVx2_ASAP7_75t_L g4745 ( 
.A(n_4684),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4706),
.Y(n_4746)
);

CKINVDCx20_ASAP7_75t_R g4747 ( 
.A(n_4678),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4711),
.Y(n_4748)
);

INVxp67_ASAP7_75t_L g4749 ( 
.A(n_4656),
.Y(n_4749)
);

OR2x2_ASAP7_75t_L g4750 ( 
.A(n_4705),
.B(n_4555),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4713),
.Y(n_4751)
);

AND2x2_ASAP7_75t_L g4752 ( 
.A(n_4680),
.B(n_4567),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4725),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4715),
.Y(n_4754)
);

AND2x4_ASAP7_75t_L g4755 ( 
.A(n_4726),
.B(n_4641),
.Y(n_4755)
);

INVx3_ASAP7_75t_L g4756 ( 
.A(n_4726),
.Y(n_4756)
);

BUFx3_ASAP7_75t_L g4757 ( 
.A(n_4664),
.Y(n_4757)
);

OR2x2_ASAP7_75t_L g4758 ( 
.A(n_4690),
.B(n_4596),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4718),
.Y(n_4759)
);

OR2x2_ASAP7_75t_L g4760 ( 
.A(n_4663),
.B(n_4607),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4731),
.Y(n_4761)
);

NAND2x1p5_ASAP7_75t_L g4762 ( 
.A(n_4659),
.B(n_4154),
.Y(n_4762)
);

OR2x2_ASAP7_75t_L g4763 ( 
.A(n_4708),
.B(n_4619),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4719),
.Y(n_4764)
);

INVx2_ASAP7_75t_L g4765 ( 
.A(n_4689),
.Y(n_4765)
);

OR2x2_ASAP7_75t_L g4766 ( 
.A(n_4679),
.B(n_4647),
.Y(n_4766)
);

AND2x2_ASAP7_75t_L g4767 ( 
.A(n_4668),
.B(n_4612),
.Y(n_4767)
);

AND2x4_ASAP7_75t_L g4768 ( 
.A(n_4697),
.B(n_4644),
.Y(n_4768)
);

INVx2_ASAP7_75t_L g4769 ( 
.A(n_4691),
.Y(n_4769)
);

INVx2_ASAP7_75t_L g4770 ( 
.A(n_4700),
.Y(n_4770)
);

INVx4_ASAP7_75t_L g4771 ( 
.A(n_4685),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4701),
.Y(n_4772)
);

BUFx2_ASAP7_75t_L g4773 ( 
.A(n_4702),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4654),
.Y(n_4774)
);

INVx2_ASAP7_75t_L g4775 ( 
.A(n_4721),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4657),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4660),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4712),
.B(n_4647),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4730),
.B(n_4707),
.Y(n_4779)
);

AND2x2_ASAP7_75t_L g4780 ( 
.A(n_4710),
.B(n_4612),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4665),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4673),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_4728),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4728),
.Y(n_4784)
);

INVx2_ASAP7_75t_L g4785 ( 
.A(n_4670),
.Y(n_4785)
);

INVx1_ASAP7_75t_L g4786 ( 
.A(n_4686),
.Y(n_4786)
);

AND2x4_ASAP7_75t_L g4787 ( 
.A(n_4722),
.B(n_4644),
.Y(n_4787)
);

AND2x2_ASAP7_75t_L g4788 ( 
.A(n_4655),
.B(n_4624),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4699),
.B(n_4623),
.Y(n_4789)
);

INVx1_ASAP7_75t_SL g4790 ( 
.A(n_4683),
.Y(n_4790)
);

OR2x2_ASAP7_75t_L g4791 ( 
.A(n_4693),
.B(n_4627),
.Y(n_4791)
);

AND2x2_ASAP7_75t_L g4792 ( 
.A(n_4709),
.B(n_4551),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4694),
.B(n_4631),
.Y(n_4793)
);

AND2x4_ASAP7_75t_SL g4794 ( 
.A(n_4685),
.B(n_4162),
.Y(n_4794)
);

AND2x2_ASAP7_75t_L g4795 ( 
.A(n_4722),
.B(n_4551),
.Y(n_4795)
);

AND2x2_ASAP7_75t_L g4796 ( 
.A(n_4674),
.B(n_4632),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4651),
.Y(n_4797)
);

INVx3_ASAP7_75t_L g4798 ( 
.A(n_4714),
.Y(n_4798)
);

AOI221xp5_ASAP7_75t_L g4799 ( 
.A1(n_4661),
.A2(n_4662),
.B1(n_4727),
.B2(n_4724),
.C(n_4681),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4720),
.B(n_4568),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4651),
.B(n_4559),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4703),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4695),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4723),
.Y(n_4804)
);

INVx1_ASAP7_75t_SL g4805 ( 
.A(n_4773),
.Y(n_4805)
);

NAND2x1_ASAP7_75t_L g4806 ( 
.A(n_4744),
.B(n_4714),
.Y(n_4806)
);

INVx2_ASAP7_75t_L g4807 ( 
.A(n_4745),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4793),
.Y(n_4808)
);

OAI22xp5_ASAP7_75t_L g4809 ( 
.A1(n_4771),
.A2(n_4799),
.B1(n_4756),
.B2(n_4753),
.Y(n_4809)
);

BUFx2_ASAP7_75t_L g4810 ( 
.A(n_4771),
.Y(n_4810)
);

INVx2_ASAP7_75t_L g4811 ( 
.A(n_4751),
.Y(n_4811)
);

NAND4xp25_ASAP7_75t_L g4812 ( 
.A(n_4739),
.B(n_4716),
.C(n_4704),
.D(n_4687),
.Y(n_4812)
);

AOI22xp33_ASAP7_75t_L g4813 ( 
.A1(n_4742),
.A2(n_4682),
.B1(n_4729),
.B2(n_4266),
.Y(n_4813)
);

HB1xp67_ASAP7_75t_L g4814 ( 
.A(n_4738),
.Y(n_4814)
);

BUFx3_ASAP7_75t_L g4815 ( 
.A(n_4747),
.Y(n_4815)
);

OAI22xp33_ASAP7_75t_L g4816 ( 
.A1(n_4756),
.A2(n_4723),
.B1(n_4255),
.B2(n_4672),
.Y(n_4816)
);

AO31x2_ASAP7_75t_L g4817 ( 
.A1(n_4804),
.A2(n_4797),
.A3(n_4789),
.B(n_4801),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4766),
.Y(n_4818)
);

AND2x2_ASAP7_75t_L g4819 ( 
.A(n_4734),
.B(n_4792),
.Y(n_4819)
);

CKINVDCx5p33_ASAP7_75t_R g4820 ( 
.A(n_4736),
.Y(n_4820)
);

A2O1A1Ixp33_ASAP7_75t_L g4821 ( 
.A1(n_4794),
.A2(n_4692),
.B(n_4200),
.C(n_4723),
.Y(n_4821)
);

OAI21xp5_ASAP7_75t_L g4822 ( 
.A1(n_4744),
.A2(n_4461),
.B(n_4531),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4743),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4741),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4763),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4750),
.Y(n_4826)
);

BUFx3_ASAP7_75t_L g4827 ( 
.A(n_4736),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4746),
.Y(n_4828)
);

AND2x2_ASAP7_75t_L g4829 ( 
.A(n_4768),
.B(n_4648),
.Y(n_4829)
);

AOI22xp33_ASAP7_75t_SL g4830 ( 
.A1(n_4798),
.A2(n_4473),
.B1(n_4369),
.B2(n_4370),
.Y(n_4830)
);

AND2x2_ASAP7_75t_L g4831 ( 
.A(n_4768),
.B(n_4648),
.Y(n_4831)
);

INVxp67_ASAP7_75t_L g4832 ( 
.A(n_4733),
.Y(n_4832)
);

AOI22xp33_ASAP7_75t_L g4833 ( 
.A1(n_4798),
.A2(n_4749),
.B1(n_4803),
.B2(n_4800),
.Y(n_4833)
);

AO31x2_ASAP7_75t_L g4834 ( 
.A1(n_4797),
.A2(n_4635),
.A3(n_4192),
.B(n_3489),
.Y(n_4834)
);

INVxp67_ASAP7_75t_L g4835 ( 
.A(n_4757),
.Y(n_4835)
);

INVx2_ASAP7_75t_L g4836 ( 
.A(n_4761),
.Y(n_4836)
);

AOI22xp33_ASAP7_75t_L g4837 ( 
.A1(n_4803),
.A2(n_4489),
.B1(n_4594),
.B2(n_4543),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4748),
.Y(n_4838)
);

AOI21xp5_ASAP7_75t_L g4839 ( 
.A1(n_4737),
.A2(n_4676),
.B(n_4277),
.Y(n_4839)
);

OA21x2_ASAP7_75t_L g4840 ( 
.A1(n_4783),
.A2(n_4446),
.B(n_4599),
.Y(n_4840)
);

AOI211xp5_ASAP7_75t_L g4841 ( 
.A1(n_4755),
.A2(n_4541),
.B(n_4503),
.C(n_4153),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4754),
.Y(n_4842)
);

AND4x1_ASAP7_75t_L g4843 ( 
.A(n_4762),
.B(n_4253),
.C(n_4523),
.D(n_4026),
.Y(n_4843)
);

OAI21x1_ASAP7_75t_L g4844 ( 
.A1(n_4735),
.A2(n_4784),
.B(n_4795),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4814),
.Y(n_4845)
);

BUFx2_ASAP7_75t_L g4846 ( 
.A(n_4810),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4808),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4805),
.B(n_4755),
.Y(n_4848)
);

OAI22xp5_ASAP7_75t_L g4849 ( 
.A1(n_4833),
.A2(n_4802),
.B1(n_4778),
.B2(n_4779),
.Y(n_4849)
);

NAND2xp33_ASAP7_75t_R g4850 ( 
.A(n_4820),
.B(n_4787),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4824),
.B(n_4759),
.Y(n_4851)
);

AOI211x1_ASAP7_75t_L g4852 ( 
.A1(n_4809),
.A2(n_4752),
.B(n_4767),
.C(n_4740),
.Y(n_4852)
);

AOI221xp5_ASAP7_75t_L g4853 ( 
.A1(n_4812),
.A2(n_4774),
.B1(n_4781),
.B2(n_4777),
.C(n_4776),
.Y(n_4853)
);

INVx1_ASAP7_75t_L g4854 ( 
.A(n_4818),
.Y(n_4854)
);

INVx4_ASAP7_75t_L g4855 ( 
.A(n_4827),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4823),
.B(n_4764),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4837),
.B(n_4782),
.Y(n_4857)
);

BUFx3_ASAP7_75t_L g4858 ( 
.A(n_4815),
.Y(n_4858)
);

AND2x2_ASAP7_75t_L g4859 ( 
.A(n_4819),
.B(n_4787),
.Y(n_4859)
);

OR2x2_ASAP7_75t_L g4860 ( 
.A(n_4825),
.B(n_4758),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4832),
.B(n_4796),
.Y(n_4861)
);

BUFx2_ASAP7_75t_L g4862 ( 
.A(n_4806),
.Y(n_4862)
);

AND2x2_ASAP7_75t_L g4863 ( 
.A(n_4829),
.B(n_4780),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4826),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4828),
.Y(n_4865)
);

AND2x2_ASAP7_75t_L g4866 ( 
.A(n_4831),
.B(n_4788),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4841),
.B(n_4822),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4836),
.Y(n_4868)
);

INVx2_ASAP7_75t_SL g4869 ( 
.A(n_4807),
.Y(n_4869)
);

HB1xp67_ASAP7_75t_L g4870 ( 
.A(n_4817),
.Y(n_4870)
);

AO21x2_ASAP7_75t_L g4871 ( 
.A1(n_4816),
.A2(n_4772),
.B(n_4447),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4838),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4842),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4811),
.Y(n_4874)
);

CKINVDCx5p33_ASAP7_75t_R g4875 ( 
.A(n_4835),
.Y(n_4875)
);

AND2x2_ASAP7_75t_L g4876 ( 
.A(n_4813),
.B(n_4790),
.Y(n_4876)
);

INVx2_ASAP7_75t_L g4877 ( 
.A(n_4817),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4817),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4844),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4840),
.Y(n_4880)
);

INVx3_ASAP7_75t_L g4881 ( 
.A(n_4840),
.Y(n_4881)
);

HB1xp67_ASAP7_75t_L g4882 ( 
.A(n_4821),
.Y(n_4882)
);

NOR2x1_ASAP7_75t_L g4883 ( 
.A(n_4839),
.B(n_4736),
.Y(n_4883)
);

NAND3xp33_ASAP7_75t_L g4884 ( 
.A(n_4843),
.B(n_4786),
.C(n_4772),
.Y(n_4884)
);

HB1xp67_ASAP7_75t_L g4885 ( 
.A(n_4834),
.Y(n_4885)
);

AND2x2_ASAP7_75t_L g4886 ( 
.A(n_4830),
.B(n_4760),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4834),
.B(n_4785),
.Y(n_4887)
);

AOI22xp5_ASAP7_75t_L g4888 ( 
.A1(n_4834),
.A2(n_4786),
.B1(n_4769),
.B2(n_4770),
.Y(n_4888)
);

AOI221xp5_ASAP7_75t_L g4889 ( 
.A1(n_4809),
.A2(n_4775),
.B1(n_4765),
.B2(n_4791),
.C(n_3399),
.Y(n_4889)
);

INVx4_ASAP7_75t_L g4890 ( 
.A(n_4820),
.Y(n_4890)
);

NAND3xp33_ASAP7_75t_L g4891 ( 
.A(n_4809),
.B(n_3620),
.C(n_3694),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4814),
.Y(n_4892)
);

BUFx6f_ASAP7_75t_L g4893 ( 
.A(n_4827),
.Y(n_4893)
);

INVx3_ASAP7_75t_L g4894 ( 
.A(n_4806),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4810),
.B(n_4465),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4814),
.Y(n_4896)
);

INVx3_ASAP7_75t_L g4897 ( 
.A(n_4855),
.Y(n_4897)
);

AND2x2_ASAP7_75t_L g4898 ( 
.A(n_4876),
.B(n_4257),
.Y(n_4898)
);

AND2x2_ASAP7_75t_L g4899 ( 
.A(n_4848),
.B(n_4259),
.Y(n_4899)
);

OAI21xp5_ASAP7_75t_L g4900 ( 
.A1(n_4867),
.A2(n_4456),
.B(n_4512),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4846),
.B(n_4450),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4855),
.B(n_4153),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4870),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4886),
.B(n_4211),
.Y(n_4904)
);

AND2x2_ASAP7_75t_L g4905 ( 
.A(n_4862),
.B(n_4215),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4845),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4892),
.Y(n_4907)
);

INVxp67_ASAP7_75t_SL g4908 ( 
.A(n_4858),
.Y(n_4908)
);

AND2x2_ASAP7_75t_L g4909 ( 
.A(n_4893),
.B(n_4205),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_SL g4910 ( 
.A(n_4883),
.B(n_4242),
.Y(n_4910)
);

AND2x4_ASAP7_75t_L g4911 ( 
.A(n_4893),
.B(n_4154),
.Y(n_4911)
);

AND2x2_ASAP7_75t_L g4912 ( 
.A(n_4893),
.B(n_4205),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4894),
.B(n_4281),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4896),
.Y(n_4914)
);

INVx2_ASAP7_75t_L g4915 ( 
.A(n_4869),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_L g4916 ( 
.A(n_4847),
.B(n_4544),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_4894),
.B(n_4242),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4859),
.B(n_4246),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4863),
.B(n_4252),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_4853),
.B(n_4516),
.Y(n_4920)
);

OR2x2_ASAP7_75t_L g4921 ( 
.A(n_4864),
.B(n_4516),
.Y(n_4921)
);

AND2x2_ASAP7_75t_L g4922 ( 
.A(n_4866),
.B(n_4228),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4878),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4851),
.Y(n_4924)
);

OR2x2_ASAP7_75t_L g4925 ( 
.A(n_4854),
.B(n_4467),
.Y(n_4925)
);

AND2x2_ASAP7_75t_L g4926 ( 
.A(n_4882),
.B(n_4228),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4877),
.Y(n_4927)
);

OR2x2_ASAP7_75t_L g4928 ( 
.A(n_4860),
.B(n_4857),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_4868),
.Y(n_4929)
);

AND2x2_ASAP7_75t_L g4930 ( 
.A(n_4861),
.B(n_4248),
.Y(n_4930)
);

OR2x2_ASAP7_75t_L g4931 ( 
.A(n_4856),
.B(n_4524),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4865),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4889),
.B(n_4457),
.Y(n_4933)
);

INVx1_ASAP7_75t_SL g4934 ( 
.A(n_4875),
.Y(n_4934)
);

OR2x2_ASAP7_75t_L g4935 ( 
.A(n_4872),
.B(n_4519),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4873),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4849),
.B(n_4509),
.Y(n_4937)
);

OR2x2_ASAP7_75t_L g4938 ( 
.A(n_4874),
.B(n_4442),
.Y(n_4938)
);

AND2x2_ASAP7_75t_L g4939 ( 
.A(n_4895),
.B(n_4248),
.Y(n_4939)
);

OR2x2_ASAP7_75t_L g4940 ( 
.A(n_4884),
.B(n_4480),
.Y(n_4940)
);

OR2x2_ASAP7_75t_L g4941 ( 
.A(n_4879),
.B(n_4487),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_L g4942 ( 
.A(n_4852),
.B(n_4448),
.Y(n_4942)
);

AND2x2_ASAP7_75t_L g4943 ( 
.A(n_4890),
.B(n_4289),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4885),
.B(n_4536),
.Y(n_4944)
);

HB1xp67_ASAP7_75t_L g4945 ( 
.A(n_4850),
.Y(n_4945)
);

OR2x2_ASAP7_75t_L g4946 ( 
.A(n_4871),
.B(n_4574),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4880),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4881),
.Y(n_4948)
);

AND2x2_ASAP7_75t_L g4949 ( 
.A(n_4890),
.B(n_4289),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4887),
.B(n_4265),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4908),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4927),
.Y(n_4952)
);

INVx1_ASAP7_75t_L g4953 ( 
.A(n_4927),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4903),
.Y(n_4954)
);

OR2x2_ASAP7_75t_L g4955 ( 
.A(n_4924),
.B(n_4891),
.Y(n_4955)
);

AND2x2_ASAP7_75t_L g4956 ( 
.A(n_4945),
.B(n_4881),
.Y(n_4956)
);

HB1xp67_ASAP7_75t_L g4957 ( 
.A(n_4947),
.Y(n_4957)
);

INVx1_ASAP7_75t_SL g4958 ( 
.A(n_4934),
.Y(n_4958)
);

OR2x2_ASAP7_75t_L g4959 ( 
.A(n_4924),
.B(n_4906),
.Y(n_4959)
);

AND2x2_ASAP7_75t_L g4960 ( 
.A(n_4897),
.B(n_4888),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4905),
.B(n_4904),
.Y(n_4961)
);

AND2x2_ASAP7_75t_L g4962 ( 
.A(n_4897),
.B(n_4494),
.Y(n_4962)
);

AND2x2_ASAP7_75t_L g4963 ( 
.A(n_4913),
.B(n_4325),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4947),
.Y(n_4964)
);

INVx2_ASAP7_75t_SL g4965 ( 
.A(n_4902),
.Y(n_4965)
);

NAND2x1p5_ASAP7_75t_L g4966 ( 
.A(n_4911),
.B(n_4325),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4907),
.Y(n_4967)
);

HB1xp67_ASAP7_75t_L g4968 ( 
.A(n_4914),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4933),
.B(n_3706),
.Y(n_4969)
);

NOR2x1p5_ASAP7_75t_SL g4970 ( 
.A(n_4948),
.B(n_3532),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4917),
.B(n_4303),
.Y(n_4971)
);

OR2x2_ASAP7_75t_L g4972 ( 
.A(n_4928),
.B(n_714),
.Y(n_4972)
);

NOR2xp33_ASAP7_75t_L g4973 ( 
.A(n_4898),
.B(n_715),
.Y(n_4973)
);

AND2x2_ASAP7_75t_L g4974 ( 
.A(n_4926),
.B(n_4303),
.Y(n_4974)
);

INVx2_ASAP7_75t_L g4975 ( 
.A(n_4948),
.Y(n_4975)
);

OR2x2_ASAP7_75t_L g4976 ( 
.A(n_4929),
.B(n_715),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4923),
.Y(n_4977)
);

AND2x4_ASAP7_75t_L g4978 ( 
.A(n_4943),
.B(n_4532),
.Y(n_4978)
);

AND2x2_ASAP7_75t_L g4979 ( 
.A(n_4950),
.B(n_4305),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4932),
.Y(n_4980)
);

OR2x2_ASAP7_75t_L g4981 ( 
.A(n_4921),
.B(n_716),
.Y(n_4981)
);

OR2x2_ASAP7_75t_L g4982 ( 
.A(n_4931),
.B(n_717),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4915),
.B(n_4305),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_4936),
.Y(n_4984)
);

AND2x4_ASAP7_75t_L g4985 ( 
.A(n_4949),
.B(n_4525),
.Y(n_4985)
);

OR2x2_ASAP7_75t_L g4986 ( 
.A(n_4937),
.B(n_718),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4944),
.Y(n_4987)
);

CKINVDCx16_ASAP7_75t_R g4988 ( 
.A(n_4958),
.Y(n_4988)
);

OR2x2_ASAP7_75t_L g4989 ( 
.A(n_4951),
.B(n_4916),
.Y(n_4989)
);

INVxp67_ASAP7_75t_SL g4990 ( 
.A(n_4951),
.Y(n_4990)
);

OR2x2_ASAP7_75t_L g4991 ( 
.A(n_4955),
.B(n_4901),
.Y(n_4991)
);

AND2x2_ASAP7_75t_L g4992 ( 
.A(n_4965),
.B(n_4899),
.Y(n_4992)
);

INVx2_ASAP7_75t_SL g4993 ( 
.A(n_4983),
.Y(n_4993)
);

AND2x4_ASAP7_75t_L g4994 ( 
.A(n_4956),
.B(n_4911),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4957),
.Y(n_4995)
);

AOI21xp5_ASAP7_75t_L g4996 ( 
.A1(n_4960),
.A2(n_4910),
.B(n_4942),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4974),
.B(n_4909),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_4961),
.B(n_4920),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4964),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4975),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4971),
.B(n_4912),
.Y(n_5001)
);

AND2x2_ASAP7_75t_L g5002 ( 
.A(n_4979),
.B(n_4919),
.Y(n_5002)
);

OR2x2_ASAP7_75t_L g5003 ( 
.A(n_4972),
.B(n_4941),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4963),
.B(n_4918),
.Y(n_5004)
);

AND2x2_ASAP7_75t_L g5005 ( 
.A(n_4973),
.B(n_4939),
.Y(n_5005)
);

AND2x2_ASAP7_75t_L g5006 ( 
.A(n_4982),
.B(n_4930),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4986),
.B(n_4969),
.Y(n_5007)
);

AND2x2_ASAP7_75t_L g5008 ( 
.A(n_4987),
.B(n_4922),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4968),
.Y(n_5009)
);

AO21x2_ASAP7_75t_L g5010 ( 
.A1(n_4954),
.A2(n_4946),
.B(n_4940),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4952),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4953),
.Y(n_5012)
);

AND2x2_ASAP7_75t_L g5013 ( 
.A(n_4976),
.B(n_4938),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4959),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4962),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4967),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4977),
.Y(n_5017)
);

XOR2xp5_ASAP7_75t_L g5018 ( 
.A(n_4981),
.B(n_4900),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4980),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_SL g5020 ( 
.A(n_4984),
.B(n_4935),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4978),
.Y(n_5021)
);

INVx3_ASAP7_75t_L g5022 ( 
.A(n_4966),
.Y(n_5022)
);

INVx2_ASAP7_75t_L g5023 ( 
.A(n_4985),
.Y(n_5023)
);

AND2x2_ASAP7_75t_L g5024 ( 
.A(n_4978),
.B(n_4985),
.Y(n_5024)
);

INVx1_ASAP7_75t_L g5025 ( 
.A(n_4970),
.Y(n_5025)
);

NOR2xp33_ASAP7_75t_L g5026 ( 
.A(n_4958),
.B(n_4925),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_4951),
.B(n_718),
.Y(n_5027)
);

HB1xp67_ASAP7_75t_L g5028 ( 
.A(n_4951),
.Y(n_5028)
);

AND2x2_ASAP7_75t_L g5029 ( 
.A(n_4958),
.B(n_719),
.Y(n_5029)
);

INVx2_ASAP7_75t_L g5030 ( 
.A(n_4951),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_L g5031 ( 
.A(n_4951),
.B(n_719),
.Y(n_5031)
);

INVx1_ASAP7_75t_SL g5032 ( 
.A(n_4958),
.Y(n_5032)
);

INVx1_ASAP7_75t_SL g5033 ( 
.A(n_4958),
.Y(n_5033)
);

INVx1_ASAP7_75t_L g5034 ( 
.A(n_4951),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_5028),
.Y(n_5035)
);

INVxp67_ASAP7_75t_L g5036 ( 
.A(n_4990),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_4988),
.B(n_720),
.Y(n_5037)
);

NAND2xp33_ASAP7_75t_SL g5038 ( 
.A(n_4991),
.B(n_3479),
.Y(n_5038)
);

AND2x2_ASAP7_75t_L g5039 ( 
.A(n_5032),
.B(n_721),
.Y(n_5039)
);

INVx2_ASAP7_75t_L g5040 ( 
.A(n_5033),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_5002),
.B(n_722),
.Y(n_5041)
);

INVxp67_ASAP7_75t_L g5042 ( 
.A(n_5029),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_5030),
.B(n_722),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_5025),
.B(n_724),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_5004),
.B(n_724),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_L g5046 ( 
.A(n_5025),
.B(n_725),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_5034),
.Y(n_5047)
);

AND2x2_ASAP7_75t_L g5048 ( 
.A(n_4992),
.B(n_4994),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4995),
.Y(n_5049)
);

OR2x2_ASAP7_75t_L g5050 ( 
.A(n_5027),
.B(n_725),
.Y(n_5050)
);

OR2x2_ASAP7_75t_L g5051 ( 
.A(n_5031),
.B(n_726),
.Y(n_5051)
);

AND2x2_ASAP7_75t_L g5052 ( 
.A(n_4994),
.B(n_727),
.Y(n_5052)
);

AOI33xp33_ASAP7_75t_L g5053 ( 
.A1(n_5014),
.A2(n_4038),
.A3(n_3691),
.B1(n_3745),
.B2(n_729),
.B3(n_731),
.Y(n_5053)
);

AND2x2_ASAP7_75t_L g5054 ( 
.A(n_5001),
.B(n_4997),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_5000),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_5009),
.Y(n_5056)
);

NOR2x1_ASAP7_75t_L g5057 ( 
.A(n_5011),
.B(n_3749),
.Y(n_5057)
);

OR2x2_ASAP7_75t_L g5058 ( 
.A(n_4989),
.B(n_727),
.Y(n_5058)
);

OR2x2_ASAP7_75t_L g5059 ( 
.A(n_5007),
.B(n_728),
.Y(n_5059)
);

AND2x4_ASAP7_75t_L g5060 ( 
.A(n_4993),
.B(n_728),
.Y(n_5060)
);

INVx1_ASAP7_75t_SL g5061 ( 
.A(n_5022),
.Y(n_5061)
);

AND2x2_ASAP7_75t_L g5062 ( 
.A(n_5006),
.B(n_729),
.Y(n_5062)
);

INVx1_ASAP7_75t_SL g5063 ( 
.A(n_5022),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_5011),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_5026),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_5008),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_5021),
.B(n_730),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_5021),
.B(n_730),
.Y(n_5068)
);

NOR3xp33_ASAP7_75t_SL g5069 ( 
.A(n_4996),
.B(n_3272),
.C(n_3248),
.Y(n_5069)
);

NAND2x1_ASAP7_75t_L g5070 ( 
.A(n_5023),
.B(n_4271),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_5013),
.B(n_732),
.Y(n_5071)
);

AND2x2_ASAP7_75t_L g5072 ( 
.A(n_5005),
.B(n_732),
.Y(n_5072)
);

OR2x2_ASAP7_75t_L g5073 ( 
.A(n_5003),
.B(n_733),
.Y(n_5073)
);

NOR2xp33_ASAP7_75t_L g5074 ( 
.A(n_5061),
.B(n_4998),
.Y(n_5074)
);

AOI32xp33_ASAP7_75t_L g5075 ( 
.A1(n_5063),
.A2(n_5048),
.A3(n_5040),
.B1(n_5065),
.B2(n_5066),
.Y(n_5075)
);

OR2x2_ASAP7_75t_L g5076 ( 
.A(n_5044),
.B(n_5015),
.Y(n_5076)
);

HB1xp67_ASAP7_75t_L g5077 ( 
.A(n_5039),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_5037),
.Y(n_5078)
);

INVx1_ASAP7_75t_SL g5079 ( 
.A(n_5052),
.Y(n_5079)
);

INVx2_ASAP7_75t_L g5080 ( 
.A(n_5054),
.Y(n_5080)
);

AOI21xp33_ASAP7_75t_L g5081 ( 
.A1(n_5036),
.A2(n_5017),
.B(n_5016),
.Y(n_5081)
);

OAI22xp33_ASAP7_75t_L g5082 ( 
.A1(n_5046),
.A2(n_5019),
.B1(n_4999),
.B2(n_5012),
.Y(n_5082)
);

OR2x2_ASAP7_75t_L g5083 ( 
.A(n_5071),
.B(n_5020),
.Y(n_5083)
);

AOI21xp33_ASAP7_75t_L g5084 ( 
.A1(n_5035),
.A2(n_5018),
.B(n_5010),
.Y(n_5084)
);

INVx1_ASAP7_75t_SL g5085 ( 
.A(n_5060),
.Y(n_5085)
);

O2A1O1Ixp33_ASAP7_75t_SL g5086 ( 
.A1(n_5067),
.A2(n_5024),
.B(n_3398),
.C(n_3388),
.Y(n_5086)
);

AND2x2_ASAP7_75t_L g5087 ( 
.A(n_5041),
.B(n_734),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_5060),
.B(n_735),
.Y(n_5088)
);

OR2x2_ASAP7_75t_L g5089 ( 
.A(n_5068),
.B(n_735),
.Y(n_5089)
);

AOI21xp33_ASAP7_75t_L g5090 ( 
.A1(n_5035),
.A2(n_737),
.B(n_738),
.Y(n_5090)
);

OR2x2_ASAP7_75t_L g5091 ( 
.A(n_5043),
.B(n_737),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_5045),
.B(n_738),
.Y(n_5092)
);

INVx2_ASAP7_75t_SL g5093 ( 
.A(n_5070),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_5072),
.B(n_739),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_L g5095 ( 
.A(n_5062),
.B(n_739),
.Y(n_5095)
);

AOI222xp33_ASAP7_75t_L g5096 ( 
.A1(n_5055),
.A2(n_3495),
.B1(n_3487),
.B2(n_3503),
.C1(n_3491),
.C2(n_3481),
.Y(n_5096)
);

INVx1_ASAP7_75t_SL g5097 ( 
.A(n_5050),
.Y(n_5097)
);

OAI22xp33_ASAP7_75t_SL g5098 ( 
.A1(n_5058),
.A2(n_3506),
.B1(n_3515),
.B2(n_3511),
.Y(n_5098)
);

AOI22xp33_ASAP7_75t_L g5099 ( 
.A1(n_5038),
.A2(n_3766),
.B1(n_3754),
.B2(n_3707),
.Y(n_5099)
);

OR2x2_ASAP7_75t_L g5100 ( 
.A(n_5073),
.B(n_740),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_5051),
.Y(n_5101)
);

OR2x2_ASAP7_75t_L g5102 ( 
.A(n_5059),
.B(n_741),
.Y(n_5102)
);

OR2x2_ASAP7_75t_L g5103 ( 
.A(n_5056),
.B(n_741),
.Y(n_5103)
);

OAI21xp33_ASAP7_75t_SL g5104 ( 
.A1(n_5049),
.A2(n_3537),
.B(n_3535),
.Y(n_5104)
);

OAI22xp5_ASAP7_75t_L g5105 ( 
.A1(n_5042),
.A2(n_3708),
.B1(n_3742),
.B2(n_3273),
.Y(n_5105)
);

AND2x4_ASAP7_75t_L g5106 ( 
.A(n_5047),
.B(n_742),
.Y(n_5106)
);

OAI21xp33_ASAP7_75t_SL g5107 ( 
.A1(n_5064),
.A2(n_3542),
.B(n_3538),
.Y(n_5107)
);

OR2x2_ASAP7_75t_L g5108 ( 
.A(n_5069),
.B(n_744),
.Y(n_5108)
);

OR2x2_ASAP7_75t_L g5109 ( 
.A(n_5057),
.B(n_744),
.Y(n_5109)
);

INVx2_ASAP7_75t_L g5110 ( 
.A(n_5053),
.Y(n_5110)
);

OAI221xp5_ASAP7_75t_SL g5111 ( 
.A1(n_5061),
.A2(n_3923),
.B1(n_3528),
.B2(n_3549),
.C(n_3526),
.Y(n_5111)
);

AOI22xp5_ASAP7_75t_L g5112 ( 
.A1(n_5061),
.A2(n_3555),
.B1(n_3562),
.B2(n_3525),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_5080),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_5075),
.B(n_745),
.Y(n_5114)
);

NOR2x1_ASAP7_75t_L g5115 ( 
.A(n_5103),
.B(n_3560),
.Y(n_5115)
);

NAND2xp5_ASAP7_75t_L g5116 ( 
.A(n_5085),
.B(n_745),
.Y(n_5116)
);

OA21x2_ASAP7_75t_SL g5117 ( 
.A1(n_5079),
.A2(n_3564),
.B(n_3563),
.Y(n_5117)
);

AND2x2_ASAP7_75t_L g5118 ( 
.A(n_5074),
.B(n_746),
.Y(n_5118)
);

HB1xp67_ASAP7_75t_L g5119 ( 
.A(n_5088),
.Y(n_5119)
);

OR2x2_ASAP7_75t_L g5120 ( 
.A(n_5100),
.B(n_746),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_L g5121 ( 
.A(n_5087),
.B(n_747),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_L g5122 ( 
.A(n_5110),
.B(n_747),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_5102),
.Y(n_5123)
);

XNOR2xp5_ASAP7_75t_L g5124 ( 
.A(n_5077),
.B(n_748),
.Y(n_5124)
);

NAND3xp33_ASAP7_75t_L g5125 ( 
.A(n_5090),
.B(n_3639),
.C(n_3635),
.Y(n_5125)
);

INVxp67_ASAP7_75t_L g5126 ( 
.A(n_5092),
.Y(n_5126)
);

AND2x2_ASAP7_75t_L g5127 ( 
.A(n_5093),
.B(n_748),
.Y(n_5127)
);

NAND2xp5_ASAP7_75t_SL g5128 ( 
.A(n_5084),
.B(n_3641),
.Y(n_5128)
);

AND2x4_ASAP7_75t_L g5129 ( 
.A(n_5106),
.B(n_3746),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_L g5130 ( 
.A(n_5097),
.B(n_749),
.Y(n_5130)
);

OR2x2_ASAP7_75t_L g5131 ( 
.A(n_5108),
.B(n_750),
.Y(n_5131)
);

AND2x2_ASAP7_75t_L g5132 ( 
.A(n_5101),
.B(n_5078),
.Y(n_5132)
);

NAND2xp5_ASAP7_75t_L g5133 ( 
.A(n_5094),
.B(n_750),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_5089),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_5095),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_L g5136 ( 
.A(n_5082),
.B(n_751),
.Y(n_5136)
);

AND2x2_ASAP7_75t_L g5137 ( 
.A(n_5076),
.B(n_751),
.Y(n_5137)
);

INVx2_ASAP7_75t_L g5138 ( 
.A(n_5091),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_5109),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_5098),
.B(n_752),
.Y(n_5140)
);

INVx1_ASAP7_75t_SL g5141 ( 
.A(n_5083),
.Y(n_5141)
);

INVx2_ASAP7_75t_SL g5142 ( 
.A(n_5105),
.Y(n_5142)
);

NOR3xp33_ASAP7_75t_L g5143 ( 
.A(n_5081),
.B(n_3574),
.C(n_3569),
.Y(n_5143)
);

AND2x2_ASAP7_75t_L g5144 ( 
.A(n_5104),
.B(n_752),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_5127),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_5113),
.Y(n_5146)
);

INVxp67_ASAP7_75t_SL g5147 ( 
.A(n_5116),
.Y(n_5147)
);

OR2x2_ASAP7_75t_L g5148 ( 
.A(n_5114),
.B(n_5111),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_5118),
.B(n_5107),
.Y(n_5149)
);

AND2x4_ASAP7_75t_SL g5150 ( 
.A(n_5138),
.B(n_5112),
.Y(n_5150)
);

AND2x2_ASAP7_75t_L g5151 ( 
.A(n_5137),
.B(n_5096),
.Y(n_5151)
);

NOR2xp33_ASAP7_75t_L g5152 ( 
.A(n_5141),
.B(n_5086),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_5121),
.Y(n_5153)
);

NOR2xp33_ASAP7_75t_L g5154 ( 
.A(n_5122),
.B(n_5099),
.Y(n_5154)
);

AND2x2_ASAP7_75t_L g5155 ( 
.A(n_5144),
.B(n_5132),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_5131),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_5136),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_5130),
.Y(n_5158)
);

AOI21xp5_ASAP7_75t_L g5159 ( 
.A1(n_5140),
.A2(n_3580),
.B(n_3570),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_5133),
.Y(n_5160)
);

HB1xp67_ASAP7_75t_L g5161 ( 
.A(n_5120),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_L g5162 ( 
.A(n_5124),
.B(n_753),
.Y(n_5162)
);

AOI221xp5_ASAP7_75t_L g5163 ( 
.A1(n_5123),
.A2(n_3598),
.B1(n_3604),
.B2(n_3595),
.C(n_3592),
.Y(n_5163)
);

INVxp67_ASAP7_75t_SL g5164 ( 
.A(n_5119),
.Y(n_5164)
);

INVx1_ASAP7_75t_SL g5165 ( 
.A(n_5134),
.Y(n_5165)
);

AND2x2_ASAP7_75t_L g5166 ( 
.A(n_5139),
.B(n_753),
.Y(n_5166)
);

NAND2xp5_ASAP7_75t_L g5167 ( 
.A(n_5142),
.B(n_754),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5135),
.B(n_5126),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_5115),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_5143),
.B(n_754),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_5129),
.B(n_755),
.Y(n_5171)
);

NOR2xp67_ASAP7_75t_L g5172 ( 
.A(n_5128),
.B(n_755),
.Y(n_5172)
);

INVxp67_ASAP7_75t_L g5173 ( 
.A(n_5129),
.Y(n_5173)
);

INVx2_ASAP7_75t_SL g5174 ( 
.A(n_5146),
.Y(n_5174)
);

NAND2xp5_ASAP7_75t_L g5175 ( 
.A(n_5155),
.B(n_5166),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_SL g5176 ( 
.A(n_5172),
.B(n_5162),
.Y(n_5176)
);

NAND3xp33_ASAP7_75t_L g5177 ( 
.A(n_5167),
.B(n_5125),
.C(n_5117),
.Y(n_5177)
);

AOI211xp5_ASAP7_75t_L g5178 ( 
.A1(n_5152),
.A2(n_3610),
.B(n_3611),
.C(n_3609),
.Y(n_5178)
);

NAND2xp5_ASAP7_75t_L g5179 ( 
.A(n_5165),
.B(n_756),
.Y(n_5179)
);

OAI21x1_ASAP7_75t_L g5180 ( 
.A1(n_5145),
.A2(n_3583),
.B(n_3581),
.Y(n_5180)
);

NAND4xp25_ASAP7_75t_L g5181 ( 
.A(n_5157),
.B(n_3621),
.C(n_3616),
.D(n_3625),
.Y(n_5181)
);

INVx2_ASAP7_75t_SL g5182 ( 
.A(n_5150),
.Y(n_5182)
);

NAND3xp33_ASAP7_75t_L g5183 ( 
.A(n_5164),
.B(n_3589),
.C(n_3586),
.Y(n_5183)
);

AND2x2_ASAP7_75t_L g5184 ( 
.A(n_5151),
.B(n_756),
.Y(n_5184)
);

INVx2_ASAP7_75t_SL g5185 ( 
.A(n_5171),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_5170),
.Y(n_5186)
);

NOR4xp25_ASAP7_75t_L g5187 ( 
.A(n_5168),
.B(n_3605),
.C(n_3505),
.D(n_3657),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_5161),
.Y(n_5188)
);

HB1xp67_ASAP7_75t_L g5189 ( 
.A(n_5172),
.Y(n_5189)
);

INVx2_ASAP7_75t_L g5190 ( 
.A(n_5173),
.Y(n_5190)
);

NAND3xp33_ASAP7_75t_L g5191 ( 
.A(n_5158),
.B(n_5156),
.C(n_5160),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_5147),
.Y(n_5192)
);

NAND3xp33_ASAP7_75t_L g5193 ( 
.A(n_5153),
.B(n_3716),
.C(n_3455),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_5148),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_5169),
.Y(n_5195)
);

INVxp67_ASAP7_75t_L g5196 ( 
.A(n_5182),
.Y(n_5196)
);

A2O1A1Ixp33_ASAP7_75t_L g5197 ( 
.A1(n_5190),
.A2(n_5154),
.B(n_5149),
.C(n_5159),
.Y(n_5197)
);

AOI222xp33_ASAP7_75t_L g5198 ( 
.A1(n_5194),
.A2(n_5163),
.B1(n_4534),
.B2(n_4096),
.C1(n_4595),
.C2(n_759),
.Y(n_5198)
);

NOR2xp33_ASAP7_75t_L g5199 ( 
.A(n_5195),
.B(n_757),
.Y(n_5199)
);

OAI22xp33_ASAP7_75t_L g5200 ( 
.A1(n_5174),
.A2(n_3703),
.B1(n_3713),
.B2(n_3644),
.Y(n_5200)
);

AOI211xp5_ASAP7_75t_L g5201 ( 
.A1(n_5188),
.A2(n_3462),
.B(n_3464),
.C(n_3446),
.Y(n_5201)
);

NAND3xp33_ASAP7_75t_L g5202 ( 
.A(n_5179),
.B(n_3466),
.C(n_3465),
.Y(n_5202)
);

AOI211x1_ASAP7_75t_SL g5203 ( 
.A1(n_5191),
.A2(n_3692),
.B(n_3689),
.C(n_3721),
.Y(n_5203)
);

NOR2xp33_ASAP7_75t_L g5204 ( 
.A(n_5175),
.B(n_757),
.Y(n_5204)
);

OAI211xp5_ASAP7_75t_L g5205 ( 
.A1(n_5192),
.A2(n_3740),
.B(n_3378),
.C(n_3380),
.Y(n_5205)
);

NOR4xp75_ASAP7_75t_L g5206 ( 
.A(n_5176),
.B(n_760),
.C(n_758),
.D(n_759),
.Y(n_5206)
);

OAI211xp5_ASAP7_75t_L g5207 ( 
.A1(n_5184),
.A2(n_3395),
.B(n_3400),
.C(n_3355),
.Y(n_5207)
);

CKINVDCx5p33_ASAP7_75t_R g5208 ( 
.A(n_5189),
.Y(n_5208)
);

OAI21xp5_ASAP7_75t_L g5209 ( 
.A1(n_5177),
.A2(n_3727),
.B(n_3285),
.Y(n_5209)
);

AOI221xp5_ASAP7_75t_L g5210 ( 
.A1(n_5186),
.A2(n_3290),
.B1(n_3287),
.B2(n_3281),
.C(n_3422),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_5185),
.Y(n_5211)
);

AOI211xp5_ASAP7_75t_L g5212 ( 
.A1(n_5183),
.A2(n_3404),
.B(n_3405),
.C(n_3403),
.Y(n_5212)
);

HB1xp67_ASAP7_75t_L g5213 ( 
.A(n_5196),
.Y(n_5213)
);

NOR3xp33_ASAP7_75t_L g5214 ( 
.A(n_5211),
.B(n_5193),
.C(n_5180),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_5204),
.Y(n_5215)
);

AO22x2_ASAP7_75t_L g5216 ( 
.A1(n_5206),
.A2(n_5187),
.B1(n_5178),
.B2(n_5181),
.Y(n_5216)
);

AND3x2_ASAP7_75t_L g5217 ( 
.A(n_5199),
.B(n_758),
.C(n_761),
.Y(n_5217)
);

NOR3xp33_ASAP7_75t_L g5218 ( 
.A(n_5197),
.B(n_762),
.C(n_763),
.Y(n_5218)
);

AOI221xp5_ASAP7_75t_L g5219 ( 
.A1(n_5208),
.A2(n_3623),
.B1(n_3432),
.B2(n_3485),
.C(n_3493),
.Y(n_5219)
);

AOI221x1_ASAP7_75t_L g5220 ( 
.A1(n_5209),
.A2(n_3494),
.B1(n_3472),
.B2(n_3697),
.C(n_3696),
.Y(n_5220)
);

INVx1_ASAP7_75t_SL g5221 ( 
.A(n_5202),
.Y(n_5221)
);

AOI222xp33_ASAP7_75t_L g5222 ( 
.A1(n_5207),
.A2(n_3532),
.B1(n_4096),
.B2(n_766),
.C1(n_768),
.C2(n_763),
.Y(n_5222)
);

AOI221xp5_ASAP7_75t_L g5223 ( 
.A1(n_5201),
.A2(n_768),
.B1(n_764),
.B2(n_767),
.C(n_771),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_5198),
.Y(n_5224)
);

AO21x1_ASAP7_75t_L g5225 ( 
.A1(n_5212),
.A2(n_767),
.B(n_771),
.Y(n_5225)
);

OAI211xp5_ASAP7_75t_L g5226 ( 
.A1(n_5213),
.A2(n_5205),
.B(n_5210),
.C(n_5203),
.Y(n_5226)
);

OAI221xp5_ASAP7_75t_L g5227 ( 
.A1(n_5223),
.A2(n_5200),
.B1(n_775),
.B2(n_772),
.C(n_774),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_5217),
.B(n_772),
.Y(n_5228)
);

AOI21xp5_ASAP7_75t_L g5229 ( 
.A1(n_5218),
.A2(n_774),
.B(n_775),
.Y(n_5229)
);

AOI322xp5_ASAP7_75t_L g5230 ( 
.A1(n_5224),
.A2(n_776),
.A3(n_777),
.B1(n_778),
.B2(n_779),
.C1(n_780),
.C2(n_781),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5216),
.B(n_778),
.Y(n_5231)
);

NOR3xp33_ASAP7_75t_L g5232 ( 
.A(n_5215),
.B(n_782),
.C(n_783),
.Y(n_5232)
);

NOR2xp33_ASAP7_75t_SL g5233 ( 
.A(n_5221),
.B(n_784),
.Y(n_5233)
);

BUFx2_ASAP7_75t_L g5234 ( 
.A(n_5231),
.Y(n_5234)
);

NOR3xp33_ASAP7_75t_L g5235 ( 
.A(n_5232),
.B(n_5214),
.C(n_5225),
.Y(n_5235)
);

OR2x2_ASAP7_75t_L g5236 ( 
.A(n_5228),
.B(n_5216),
.Y(n_5236)
);

NAND2xp5_ASAP7_75t_SL g5237 ( 
.A(n_5230),
.B(n_5222),
.Y(n_5237)
);

INVx5_ASAP7_75t_L g5238 ( 
.A(n_5233),
.Y(n_5238)
);

O2A1O1Ixp33_ASAP7_75t_L g5239 ( 
.A1(n_5227),
.A2(n_5219),
.B(n_5220),
.C(n_787),
.Y(n_5239)
);

NOR3xp33_ASAP7_75t_L g5240 ( 
.A(n_5229),
.B(n_785),
.C(n_786),
.Y(n_5240)
);

CKINVDCx5p33_ASAP7_75t_R g5241 ( 
.A(n_5226),
.Y(n_5241)
);

NAND2xp33_ASAP7_75t_R g5242 ( 
.A(n_5241),
.B(n_785),
.Y(n_5242)
);

CKINVDCx16_ASAP7_75t_R g5243 ( 
.A(n_5236),
.Y(n_5243)
);

CKINVDCx14_ASAP7_75t_R g5244 ( 
.A(n_5234),
.Y(n_5244)
);

OR2x2_ASAP7_75t_L g5245 ( 
.A(n_5237),
.B(n_786),
.Y(n_5245)
);

AO21x2_ASAP7_75t_L g5246 ( 
.A1(n_5245),
.A2(n_5235),
.B(n_5240),
.Y(n_5246)
);

OAI22xp5_ASAP7_75t_L g5247 ( 
.A1(n_5243),
.A2(n_5238),
.B1(n_5239),
.B2(n_789),
.Y(n_5247)
);

NAND2xp5_ASAP7_75t_L g5248 ( 
.A(n_5244),
.B(n_5238),
.Y(n_5248)
);

OAI221xp5_ASAP7_75t_L g5249 ( 
.A1(n_5242),
.A2(n_789),
.B1(n_787),
.B2(n_788),
.C(n_791),
.Y(n_5249)
);

NAND3xp33_ASAP7_75t_L g5250 ( 
.A(n_5242),
.B(n_791),
.C(n_792),
.Y(n_5250)
);

OAI22xp5_ASAP7_75t_L g5251 ( 
.A1(n_5243),
.A2(n_794),
.B1(n_792),
.B2(n_793),
.Y(n_5251)
);

O2A1O1Ixp5_ASAP7_75t_L g5252 ( 
.A1(n_5247),
.A2(n_5248),
.B(n_5251),
.C(n_5250),
.Y(n_5252)
);

BUFx8_ASAP7_75t_L g5253 ( 
.A(n_5246),
.Y(n_5253)
);

OAI321xp33_ASAP7_75t_L g5254 ( 
.A1(n_5249),
.A2(n_798),
.A3(n_800),
.B1(n_794),
.B2(n_795),
.C(n_799),
.Y(n_5254)
);

XNOR2xp5_ASAP7_75t_L g5255 ( 
.A(n_5247),
.B(n_795),
.Y(n_5255)
);

BUFx2_ASAP7_75t_L g5256 ( 
.A(n_5253),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5255),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5252),
.Y(n_5258)
);

INVx2_ASAP7_75t_L g5259 ( 
.A(n_5254),
.Y(n_5259)
);

INVx2_ASAP7_75t_L g5260 ( 
.A(n_5253),
.Y(n_5260)
);

HB1xp67_ASAP7_75t_L g5261 ( 
.A(n_5258),
.Y(n_5261)
);

AOI21xp5_ASAP7_75t_L g5262 ( 
.A1(n_5259),
.A2(n_4634),
.B(n_799),
.Y(n_5262)
);

AO22x2_ASAP7_75t_L g5263 ( 
.A1(n_5260),
.A2(n_804),
.B1(n_801),
.B2(n_802),
.Y(n_5263)
);

OAI22xp5_ASAP7_75t_L g5264 ( 
.A1(n_5257),
.A2(n_805),
.B1(n_801),
.B2(n_804),
.Y(n_5264)
);

OR2x2_ASAP7_75t_L g5265 ( 
.A(n_5261),
.B(n_5256),
.Y(n_5265)
);

NAND2xp5_ASAP7_75t_L g5266 ( 
.A(n_5263),
.B(n_805),
.Y(n_5266)
);

AOI221xp5_ASAP7_75t_L g5267 ( 
.A1(n_5266),
.A2(n_5262),
.B1(n_5264),
.B2(n_809),
.C(n_806),
.Y(n_5267)
);

AOI22xp33_ASAP7_75t_SL g5268 ( 
.A1(n_5267),
.A2(n_5265),
.B1(n_810),
.B2(n_806),
.Y(n_5268)
);

AOI22xp33_ASAP7_75t_SL g5269 ( 
.A1(n_5268),
.A2(n_812),
.B1(n_807),
.B2(n_811),
.Y(n_5269)
);

OR2x6_ASAP7_75t_L g5270 ( 
.A(n_5269),
.B(n_811),
.Y(n_5270)
);

AOI21xp5_ASAP7_75t_L g5271 ( 
.A1(n_5270),
.A2(n_812),
.B(n_813),
.Y(n_5271)
);

AOI211xp5_ASAP7_75t_L g5272 ( 
.A1(n_5271),
.A2(n_815),
.B(n_813),
.C(n_814),
.Y(n_5272)
);


endmodule