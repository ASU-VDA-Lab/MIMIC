module fake_jpeg_17462_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_8),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_39),
.Y(n_42)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_22),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_28),
.B1(n_21),
.B2(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_15),
.B1(n_28),
.B2(n_16),
.Y(n_62)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_80),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_68),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_48),
.B1(n_28),
.B2(n_36),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_74),
.B1(n_79),
.B2(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_39),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_21),
.B1(n_16),
.B2(n_69),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_66),
.B1(n_31),
.B2(n_18),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_98),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_105),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_35),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_57),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_71),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_32),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_46),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_32),
.C(n_26),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_34),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_37),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_21),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_26),
.B(n_31),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_70),
.B1(n_74),
.B2(n_28),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_133),
.B1(n_95),
.B2(n_85),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_45),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_114),
.A2(n_120),
.B(n_121),
.Y(n_162)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_90),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_138),
.B1(n_100),
.B2(n_103),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_66),
.B1(n_21),
.B2(n_40),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_86),
.B1(n_111),
.B2(n_85),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_64),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_140),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_83),
.B(n_61),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_26),
.B(n_31),
.C(n_25),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_126),
.B(n_132),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_26),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_131),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_22),
.Y(n_132)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_128),
.Y(n_171)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_78),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_141),
.A2(n_148),
.B1(n_115),
.B2(n_19),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_142),
.B(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_89),
.B1(n_98),
.B2(n_88),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_143),
.A2(n_144),
.B1(n_169),
.B2(n_126),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_111),
.B1(n_96),
.B2(n_88),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_130),
.C(n_134),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_145),
.B(n_150),
.C(n_158),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_109),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_112),
.B1(n_107),
.B2(n_91),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_100),
.B1(n_18),
.B2(n_17),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_172),
.B1(n_24),
.B2(n_29),
.Y(n_201)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_90),
.A3(n_104),
.B1(n_91),
.B2(n_30),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_164),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_104),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_104),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_123),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_123),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_22),
.Y(n_166)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_73),
.B1(n_25),
.B2(n_30),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_37),
.B(n_23),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_124),
.B(n_135),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_128),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_116),
.A2(n_17),
.B1(n_24),
.B2(n_23),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_121),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_174),
.A2(n_182),
.B(n_141),
.Y(n_213)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_179),
.B(n_184),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_197),
.B(n_19),
.Y(n_220)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_132),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_199),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_124),
.B(n_117),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_149),
.B1(n_144),
.B2(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_202),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_127),
.B(n_29),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_133),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_188),
.B1(n_29),
.B2(n_180),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_157),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_162),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_192),
.B(n_176),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_225),
.B(n_227),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_149),
.B1(n_145),
.B2(n_147),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_212),
.A2(n_218),
.B1(n_189),
.B2(n_173),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_183),
.B(n_182),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_150),
.C(n_158),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_184),
.C(n_182),
.Y(n_233)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_143),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_115),
.B1(n_170),
.B2(n_2),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_19),
.B1(n_27),
.B2(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_201),
.B1(n_197),
.B2(n_175),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_189),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_178),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_183),
.A2(n_0),
.B(n_1),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_229),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_234),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_232),
.B(n_235),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_220),
.C(n_207),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_187),
.B1(n_185),
.B2(n_191),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_218),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_185),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_203),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_217),
.A2(n_1),
.B1(n_61),
.B2(n_4),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_27),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_27),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_247),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_10),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_213),
.B(n_203),
.C(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_260),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_210),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_261),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_257),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_262),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_243),
.A2(n_208),
.B1(n_225),
.B2(n_224),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_256),
.A2(n_232),
.B1(n_223),
.B2(n_224),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_263),
.C(n_236),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_208),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_227),
.B(n_211),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_215),
.C(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_276),
.C(n_277),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_215),
.B(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_249),
.A2(n_234),
.B1(n_247),
.B2(n_207),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_242),
.C(n_235),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_274),
.C(n_259),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_275),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_241),
.C(n_216),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_10),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_10),
.B1(n_3),
.B2(n_5),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_7),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_284),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_285),
.C(n_11),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_248),
.B1(n_253),
.B2(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_253),
.B(n_7),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_1),
.C(n_7),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_9),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_9),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_272),
.B(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_277),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_296),
.B(n_298),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_265),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_284),
.C(n_12),
.Y(n_300)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_278),
.B1(n_287),
.B2(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_11),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_304),
.B(n_290),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_293),
.A3(n_292),
.B1(n_13),
.B2(n_14),
.C1(n_12),
.C2(n_11),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_307),
.C(n_301),
.Y(n_309)
);

NAND2xp33_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_302),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_301),
.C(n_13),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_14),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_313),
.Y(n_314)
);


endmodule