module fake_jpeg_570_n_536 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_536);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_17),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_53),
.B(n_56),
.Y(n_130)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g133 ( 
.A(n_55),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_57),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g123 ( 
.A(n_64),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_65),
.B(n_74),
.Y(n_144)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_75),
.Y(n_114)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_17),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_38),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_83),
.B(n_101),
.Y(n_162)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_93),
.Y(n_127)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_92),
.B(n_94),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_15),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_37),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_47),
.Y(n_134)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_33),
.B1(n_21),
.B2(n_25),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_105),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_25),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_112),
.B(n_119),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_59),
.A2(n_39),
.B1(n_47),
.B2(n_33),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_126),
.A2(n_163),
.B1(n_36),
.B2(n_39),
.Y(n_194)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_128),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_134),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_21),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_135),
.B(n_139),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_24),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_143),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_64),
.A2(n_26),
.B1(n_29),
.B2(n_40),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_148),
.B1(n_91),
.B2(n_50),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_61),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_156),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_64),
.A2(n_26),
.B1(n_29),
.B2(n_40),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_68),
.B(n_24),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_155),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_67),
.B(n_24),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_82),
.B(n_47),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_82),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_69),
.A2(n_39),
.B1(n_29),
.B2(n_26),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_149),
.C(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_183),
.Y(n_234)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

CKINVDCx12_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_168),
.Y(n_228)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_171),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_172),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_173),
.A2(n_194),
.B1(n_136),
.B2(n_104),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_114),
.A2(n_102),
.B1(n_76),
.B2(n_95),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_174),
.A2(n_191),
.B1(n_204),
.B2(n_208),
.Y(n_239)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_101),
.B1(n_44),
.B2(n_43),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_176),
.B(n_203),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_103),
.B(n_47),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_181),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_178),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_127),
.B(n_42),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_182),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_42),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_116),
.B(n_47),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_184),
.Y(n_261)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_186),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_187),
.B(n_195),
.Y(n_248)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_117),
.A2(n_89),
.B1(n_87),
.B2(n_81),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_132),
.B(n_23),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_192),
.B(n_200),
.Y(n_238)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_115),
.A2(n_23),
.B(n_44),
.Y(n_195)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_126),
.A2(n_73),
.B1(n_66),
.B2(n_54),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_198),
.A2(n_220),
.B1(n_167),
.B2(n_172),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_150),
.B(n_41),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_199),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_108),
.B(n_43),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_146),
.B(n_41),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_142),
.A2(n_77),
.B1(n_80),
.B2(n_30),
.Y(n_204)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_148),
.A2(n_35),
.B1(n_32),
.B2(n_39),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_15),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_215),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_111),
.A2(n_36),
.B1(n_50),
.B2(n_10),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_213),
.B1(n_219),
.B2(n_104),
.Y(n_250)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_161),
.A2(n_36),
.B1(n_48),
.B2(n_93),
.Y(n_213)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_133),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_133),
.B(n_15),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_107),
.Y(n_218)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_111),
.A2(n_14),
.B1(n_11),
.B2(n_10),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_113),
.A2(n_48),
.B1(n_93),
.B2(n_2),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_113),
.B(n_0),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_0),
.C(n_1),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_159),
.B(n_10),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_0),
.Y(n_272)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_118),
.Y(n_225)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_171),
.A2(n_161),
.B1(n_157),
.B2(n_137),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_226),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_166),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_235),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_170),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_240),
.B(n_250),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_185),
.A2(n_160),
.B1(n_129),
.B2(n_147),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_256),
.B1(n_260),
.B2(n_221),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_176),
.A2(n_160),
.B1(n_136),
.B2(n_124),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_207),
.A2(n_124),
.B1(n_131),
.B2(n_140),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_202),
.B(n_122),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_180),
.B(n_157),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_140),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_186),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_274),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_2),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_199),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_184),
.B(n_152),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_275),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_109),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_188),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_183),
.B(n_203),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_278),
.A2(n_292),
.B(n_297),
.Y(n_354)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_279),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_220),
.B(n_213),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_280),
.A2(n_301),
.B(n_236),
.Y(n_338)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_231),
.Y(n_281)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

XOR2x2_ASAP7_75t_SL g332 ( 
.A(n_282),
.B(n_273),
.Y(n_332)
);

CKINVDCx11_ASAP7_75t_R g284 ( 
.A(n_253),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_284),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

BUFx24_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_288),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_291),
.Y(n_362)
);

OR2x4_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_214),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_275),
.Y(n_293)
);

BUFx24_ASAP7_75t_L g361 ( 
.A(n_293),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_258),
.Y(n_294)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_228),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_295),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_221),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_305),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_258),
.A2(n_198),
.B(n_205),
.Y(n_297)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_298),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_3),
.Y(n_363)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_300),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_212),
.B(n_225),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_231),
.Y(n_302)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_302),
.Y(n_342)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_230),
.Y(n_303)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_303),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_190),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_233),
.B(n_238),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_314),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_209),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_308),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_234),
.B(n_206),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_313),
.Y(n_343)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_241),
.Y(n_310)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

INVx3_ASAP7_75t_SL g312 ( 
.A(n_227),
.Y(n_312)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_312),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g313 ( 
.A(n_255),
.B(n_261),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_240),
.A2(n_191),
.B1(n_216),
.B2(n_169),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_315),
.A2(n_227),
.B1(n_264),
.B2(n_232),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_317),
.Y(n_345)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_319),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_265),
.B(n_197),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_321),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_277),
.B(n_196),
.Y(n_321)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_236),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_322),
.A2(n_267),
.B1(n_242),
.B2(n_247),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_239),
.A2(n_178),
.B1(n_218),
.B2(n_189),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_323),
.A2(n_249),
.B(n_245),
.Y(n_356)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_237),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_246),
.B1(n_243),
.B2(n_182),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_275),
.C(n_262),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_329),
.C(n_353),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_251),
.C(n_254),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_332),
.B(n_278),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_333),
.A2(n_339),
.B1(n_344),
.B2(n_350),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_334),
.A2(n_356),
.B1(n_311),
.B2(n_312),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_304),
.A2(n_315),
.B1(n_282),
.B2(n_296),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_335),
.A2(n_360),
.B1(n_341),
.B2(n_336),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_355),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_304),
.A2(n_323),
.B1(n_316),
.B2(n_285),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_304),
.A2(n_246),
.B1(n_179),
.B2(n_243),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_348),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_316),
.A2(n_247),
.B1(n_242),
.B2(n_217),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_286),
.B(n_263),
.C(n_267),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_292),
.A2(n_263),
.B(n_249),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_280),
.A2(n_245),
.B1(n_152),
.B2(n_107),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_297),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_301),
.A2(n_175),
.B1(n_152),
.B2(n_109),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_327),
.Y(n_366)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_366),
.Y(n_423)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_330),
.Y(n_367)
);

BUFx2_ASAP7_75t_SL g419 ( 
.A(n_367),
.Y(n_419)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_359),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_378),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_289),
.Y(n_375)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_337),
.B(n_283),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_377),
.B(n_383),
.Y(n_420)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_351),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_384),
.Y(n_415)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_364),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_380),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_385),
.Y(n_402)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_343),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_346),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_320),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_332),
.B(n_286),
.C(n_293),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_397),
.C(n_398),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_387),
.B(n_361),
.Y(n_422)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_389),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_358),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_391),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_331),
.B(n_306),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_392),
.B(n_395),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_393),
.A2(n_400),
.B1(n_339),
.B2(n_355),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_326),
.B(n_290),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_394),
.B(n_310),
.Y(n_427)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_349),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_325),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_326),
.B(n_313),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_328),
.B(n_308),
.Y(n_398)
);

CKINVDCx12_ASAP7_75t_R g399 ( 
.A(n_330),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_399),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_335),
.A2(n_341),
.B1(n_338),
.B2(n_333),
.Y(n_400)
);

XNOR2x2_ASAP7_75t_SL g405 ( 
.A(n_387),
.B(n_354),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_405),
.B(n_427),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_406),
.A2(n_375),
.B1(n_382),
.B2(n_366),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_369),
.A2(n_354),
.B1(n_345),
.B2(n_360),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_407),
.A2(n_369),
.B1(n_373),
.B2(n_344),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_411),
.Y(n_435)
);

A2O1A1O1Ixp25_ASAP7_75t_L g412 ( 
.A1(n_386),
.A2(n_329),
.B(n_361),
.C(n_353),
.D(n_300),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_363),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_422),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_376),
.A2(n_356),
.B(n_357),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_417),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_340),
.Y(n_418)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_376),
.A2(n_358),
.B(n_361),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_368),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_371),
.B(n_302),
.C(n_281),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_428),
.C(n_371),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_314),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_340),
.Y(n_430)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_430),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_404),
.A2(n_376),
.B1(n_400),
.B2(n_393),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_432),
.A2(n_434),
.B1(n_445),
.B2(n_450),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_403),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_438),
.Y(n_467)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_406),
.A2(n_382),
.B1(n_380),
.B2(n_391),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_443),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_362),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_442),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_416),
.A2(n_311),
.B1(n_350),
.B2(n_284),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_444),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_416),
.A2(n_324),
.B1(n_317),
.B2(n_288),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_447),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_431),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_448),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_425),
.B(n_389),
.C(n_279),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_430),
.C(n_428),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_402),
.A2(n_317),
.B1(n_312),
.B2(n_318),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_303),
.Y(n_451)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_451),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_402),
.A2(n_367),
.B1(n_291),
.B2(n_330),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_452),
.A2(n_456),
.B1(n_408),
.B2(n_429),
.Y(n_465)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_407),
.A2(n_322),
.B1(n_298),
.B2(n_287),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_462),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_437),
.A2(n_421),
.B(n_417),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_463),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_465),
.A2(n_441),
.B1(n_438),
.B2(n_434),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_403),
.C(n_427),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_470),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_453),
.B(n_422),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_472),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_414),
.C(n_424),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_405),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_412),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_476),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_413),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_437),
.C(n_436),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_479),
.B(n_484),
.Y(n_499)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_469),
.Y(n_482)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_482),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_457),
.C(n_432),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_467),
.A2(n_446),
.B1(n_435),
.B2(n_452),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_485),
.A2(n_408),
.B1(n_475),
.B2(n_471),
.Y(n_502)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_487),
.Y(n_496)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_476),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_488),
.B(n_489),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_464),
.A2(n_413),
.B1(n_446),
.B2(n_426),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_462),
.B(n_456),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_473),
.C(n_477),
.Y(n_500)
);

NAND3xp33_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_423),
.C(n_401),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_492),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_470),
.B(n_401),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_493),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_459),
.A2(n_443),
.B1(n_445),
.B2(n_450),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_495),
.A2(n_465),
.B1(n_460),
.B2(n_478),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_481),
.A2(n_463),
.B(n_459),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_498),
.A2(n_506),
.B(n_486),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_494),
.C(n_491),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_501),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_518)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_481),
.A2(n_472),
.B(n_408),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_485),
.A2(n_468),
.B(n_419),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_508),
.A2(n_506),
.B(n_498),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_503),
.A2(n_484),
.B1(n_479),
.B2(n_490),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_511),
.Y(n_519)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_496),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_512),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_491),
.C(n_486),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_513),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_515),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_497),
.A2(n_483),
.B1(n_295),
.B2(n_6),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_483),
.C(n_5),
.Y(n_516)
);

NOR2x1_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_504),
.Y(n_520)
);

NAND4xp25_ASAP7_75t_L g524 ( 
.A(n_518),
.B(n_505),
.C(n_501),
.D(n_502),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_520),
.B(n_524),
.Y(n_528)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_519),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_525),
.B(n_526),
.Y(n_529)
);

NAND5xp2_ASAP7_75t_L g526 ( 
.A(n_521),
.B(n_514),
.C(n_508),
.D(n_507),
.E(n_511),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_SL g527 ( 
.A1(n_523),
.A2(n_517),
.B(n_513),
.C(n_510),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_527),
.B(n_522),
.Y(n_530)
);

AOI322xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_523),
.A3(n_528),
.B1(n_527),
.B2(n_512),
.C1(n_516),
.C2(n_518),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_529),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_532),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_9),
.B(n_7),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_8),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_9),
.Y(n_536)
);


endmodule