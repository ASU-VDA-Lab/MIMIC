module fake_jpeg_11771_n_46 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_SL g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_14),
.Y(n_22)
);

BUFx2_ASAP7_75t_SL g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_25),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_12),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_18),
.B(n_16),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_33),
.B(n_31),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_10),
.C(n_9),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_11),
.C(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_27),
.C(n_5),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_27),
.B(n_5),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_39),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_42),
.C(n_6),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_2),
.B(n_6),
.C(n_7),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_7),
.B(n_8),
.Y(n_46)
);


endmodule