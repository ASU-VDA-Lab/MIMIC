module real_jpeg_3156_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

AO21x1_ASAP7_75t_L g10 ( 
.A1(n_2),
.A2(n_11),
.B(n_13),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_4),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_17),
.Y(n_28)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_18),
.B(n_25),
.C(n_29),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_8),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_17),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_15),
.B(n_16),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_15),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_17),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);


endmodule