module fake_jpeg_11364_n_641 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_641);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_641;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_62),
.Y(n_172)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_64),
.Y(n_182)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g203 ( 
.A(n_65),
.Y(n_203)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_66),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_68),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_69),
.Y(n_191)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g176 ( 
.A(n_70),
.Y(n_176)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_73),
.B(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_7),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_75),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g197 ( 
.A(n_76),
.Y(n_197)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_79),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_8),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_102),
.Y(n_147)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_84),
.Y(n_210)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_23),
.A2(n_18),
.B1(n_6),
.B2(n_10),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_87),
.B(n_121),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_57),
.Y(n_90)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_95),
.Y(n_212)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_97),
.Y(n_199)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_98),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_99),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_31),
.B(n_6),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_31),
.B(n_10),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_117),
.Y(n_152)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_110),
.Y(n_213)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_32),
.B(n_5),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_41),
.A2(n_5),
.B1(n_17),
.B2(n_16),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_51),
.B1(n_57),
.B2(n_53),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_32),
.A2(n_5),
.B1(n_17),
.B2(n_16),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_47),
.A2(n_5),
.B(n_17),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_127),
.Y(n_165)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_37),
.B(n_18),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_41),
.Y(n_128)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_36),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_129),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_133),
.A2(n_148),
.B(n_156),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_76),
.A2(n_29),
.B1(n_58),
.B2(n_33),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_82),
.A2(n_53),
.B1(n_51),
.B2(n_50),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_154),
.A2(n_185),
.B1(n_206),
.B2(n_220),
.Y(n_258)
);

INVx6_ASAP7_75t_SL g155 ( 
.A(n_76),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_155),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_78),
.A2(n_51),
.B1(n_56),
.B2(n_37),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_159),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_78),
.B(n_49),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_168),
.B(n_177),
.Y(n_288)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_49),
.Y(n_177)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

INVx5_ASAP7_75t_SL g232 ( 
.A(n_179),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_56),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_189),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_60),
.A2(n_46),
.B1(n_38),
.B2(n_42),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_188),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_100),
.B(n_38),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_69),
.B(n_46),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_190),
.B(n_198),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_75),
.B(n_42),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_221),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_70),
.Y(n_196)
);

BUFx4f_ASAP7_75t_SL g259 ( 
.A(n_196),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_77),
.B(n_45),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_79),
.B(n_26),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_200),
.B(n_1),
.Y(n_257)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_84),
.A2(n_19),
.B1(n_40),
.B2(n_45),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_86),
.B(n_19),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_128),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_SL g215 ( 
.A1(n_93),
.A2(n_40),
.B(n_44),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_215),
.B(n_28),
.C(n_2),
.Y(n_263)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_103),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_120),
.A2(n_19),
.B1(n_40),
.B2(n_26),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_59),
.B(n_12),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_106),
.B1(n_119),
.B2(n_113),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_222),
.A2(n_239),
.B1(n_240),
.B2(n_261),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_142),
.B(n_0),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_226),
.B(n_234),
.Y(n_310)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_229),
.B(n_263),
.Y(n_317)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_233),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_142),
.B(n_0),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_171),
.A2(n_118),
.B1(n_67),
.B2(n_72),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_235),
.A2(n_236),
.B1(n_277),
.B2(n_283),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_133),
.A2(n_80),
.B1(n_109),
.B2(n_99),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_154),
.A2(n_110),
.B1(n_95),
.B2(n_89),
.Y(n_237)
);

OA22x2_ASAP7_75t_SL g332 ( 
.A1(n_237),
.A2(n_285),
.B1(n_232),
.B2(n_236),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_146),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_193),
.A2(n_44),
.B1(n_36),
.B2(n_34),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_44),
.B1(n_34),
.B2(n_28),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_196),
.A2(n_165),
.B(n_168),
.C(n_177),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_241),
.A2(n_253),
.B(n_289),
.Y(n_327)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_162),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_243),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_197),
.A2(n_44),
.B1(n_34),
.B2(n_28),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_245),
.Y(n_341)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_134),
.Y(n_248)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_139),
.B(n_44),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_249),
.B(n_284),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_197),
.A2(n_34),
.B1(n_28),
.B2(n_14),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_250),
.A2(n_292),
.B1(n_141),
.B2(n_140),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_159),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_251),
.B(n_264),
.Y(n_322)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_145),
.Y(n_252)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_158),
.A2(n_150),
.B1(n_191),
.B2(n_151),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_255),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_257),
.B(n_265),
.Y(n_330)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_175),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_260),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_132),
.A2(n_28),
.B1(n_34),
.B2(n_14),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_165),
.B(n_1),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_262),
.B(n_267),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_196),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_152),
.B(n_14),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_189),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_266),
.B(n_270),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_147),
.B(n_1),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_169),
.Y(n_268)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_143),
.Y(n_269)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_190),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_167),
.Y(n_271)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_167),
.Y(n_272)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_272),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_147),
.B(n_2),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_161),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_152),
.B(n_2),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_274),
.B(n_282),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_164),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_275),
.A2(n_280),
.B1(n_295),
.B2(n_297),
.Y(n_331)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_183),
.Y(n_276)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_185),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_172),
.Y(n_278)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_278),
.Y(n_329)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_176),
.Y(n_279)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_279),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_130),
.A2(n_3),
.B1(n_4),
.B2(n_153),
.Y(n_280)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_176),
.Y(n_282)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_156),
.A2(n_3),
.B1(n_4),
.B2(n_148),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_198),
.Y(n_284)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_202),
.Y(n_286)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_286),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_169),
.Y(n_287)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_287),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_135),
.A2(n_4),
.B1(n_184),
.B2(n_210),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_149),
.Y(n_290)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_138),
.Y(n_291)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_201),
.A2(n_144),
.B1(n_163),
.B2(n_157),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_186),
.Y(n_293)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_200),
.B(n_182),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_181),
.C(n_206),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_163),
.A2(n_187),
.B1(n_170),
.B2(n_174),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_187),
.A2(n_213),
.B1(n_137),
.B2(n_192),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_299),
.Y(n_336)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_211),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_302),
.B(n_260),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_344),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_232),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_313),
.B(n_347),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_315),
.B(n_240),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_231),
.B(n_192),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_325),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_235),
.A2(n_217),
.B1(n_212),
.B2(n_216),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_321),
.A2(n_297),
.B1(n_295),
.B2(n_261),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_262),
.B(n_220),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_324),
.B(n_346),
.C(n_355),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_231),
.B(n_160),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_349),
.B1(n_230),
.B2(n_223),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_226),
.B(n_166),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_345),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_253),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_234),
.B(n_131),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_294),
.B(n_203),
.C(n_141),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_249),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_228),
.B(n_288),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_241),
.A2(n_178),
.B1(n_194),
.B2(n_203),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_254),
.B(n_294),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_354),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_267),
.B(n_273),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_263),
.B(n_229),
.C(n_281),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_229),
.B(n_290),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_244),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_259),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_360),
.B(n_389),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_344),
.A2(n_237),
.B1(n_258),
.B2(n_225),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_361),
.A2(n_372),
.B1(n_379),
.B2(n_385),
.Y(n_426)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_323),
.Y(n_362)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_362),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_341),
.A2(n_281),
.B1(n_244),
.B2(n_279),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_363),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_366),
.A2(n_341),
.B(n_357),
.Y(n_425)
);

O2A1O1Ixp33_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_237),
.B(n_289),
.C(n_247),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_367),
.A2(n_400),
.B(n_327),
.Y(n_419)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_304),
.Y(n_369)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_369),
.Y(n_412)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_317),
.B(n_224),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_371),
.B(n_378),
.C(n_384),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_375),
.B(n_376),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_223),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_332),
.A2(n_237),
.B1(n_293),
.B2(n_286),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_355),
.A2(n_246),
.B(n_299),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_381),
.A2(n_353),
.B(n_350),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_393),
.Y(n_411)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_304),
.Y(n_383)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_269),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_320),
.A2(n_255),
.B1(n_233),
.B2(n_243),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_301),
.Y(n_387)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_388),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_330),
.B(n_325),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_322),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_390),
.B(n_391),
.Y(n_415)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

BUFx8_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_336),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_320),
.A2(n_227),
.B1(n_242),
.B2(n_238),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_366),
.B1(n_369),
.B2(n_383),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_321),
.A2(n_268),
.B1(n_256),
.B2(n_287),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_399),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_396),
.B(n_397),
.Y(n_416)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_339),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_317),
.B(n_246),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_324),
.C(n_315),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_319),
.A2(n_291),
.B1(n_296),
.B2(n_259),
.Y(n_399)
);

NAND2x1p5_ASAP7_75t_L g400 ( 
.A(n_302),
.B(n_259),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_311),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_406),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_333),
.B(n_345),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_310),
.Y(n_430)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_403),
.B(n_329),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_311),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_352),
.Y(n_409)
);

XNOR2x1_ASAP7_75t_L g458 ( 
.A(n_409),
.B(n_422),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_328),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_424),
.C(n_434),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_405),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_418),
.B(n_423),
.Y(n_452)
);

AO21x1_ASAP7_75t_L g459 ( 
.A1(n_419),
.A2(n_400),
.B(n_365),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_376),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_310),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_367),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_393),
.B(n_307),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_427),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_432),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_370),
.Y(n_433)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_433),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_312),
.C(n_354),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_390),
.B(n_308),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_438),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_396),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_440),
.A2(n_442),
.B1(n_385),
.B2(n_372),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_384),
.B(n_312),
.C(n_337),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_443),
.C(n_362),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_394),
.A2(n_327),
.B1(n_331),
.B2(n_326),
.Y(n_442)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_380),
.B(n_329),
.C(n_353),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_419),
.Y(n_448)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_447),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_448),
.B(n_472),
.Y(n_499)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_408),
.Y(n_449)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_449),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_415),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_450),
.B(n_473),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_444),
.A2(n_400),
.B(n_364),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_453),
.B(n_476),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_381),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_465),
.C(n_474),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_455),
.A2(n_463),
.B1(n_423),
.B2(n_428),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_456),
.A2(n_459),
.B1(n_461),
.B2(n_425),
.Y(n_500)
);

O2A1O1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_364),
.B(n_375),
.C(n_365),
.Y(n_457)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_457),
.Y(n_491)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_460),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_426),
.A2(n_389),
.B1(n_377),
.B2(n_374),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_438),
.A2(n_373),
.B1(n_402),
.B2(n_360),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_462),
.A2(n_464),
.B1(n_475),
.B2(n_479),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_SL g463 ( 
.A1(n_418),
.A2(n_373),
.B(n_399),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_407),
.A2(n_371),
.B1(n_398),
.B2(n_395),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_414),
.B(n_422),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_415),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_467),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_413),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_368),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_471),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_407),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_409),
.B(n_391),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_429),
.A2(n_406),
.B1(n_401),
.B2(n_388),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_432),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_434),
.B(n_386),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_443),
.C(n_424),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_412),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_475),
.B1(n_479),
.B2(n_447),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_411),
.A2(n_342),
.B1(n_338),
.B2(n_403),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_416),
.B(n_397),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_481),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_487),
.A2(n_509),
.B1(n_478),
.B2(n_466),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_455),
.A2(n_442),
.B1(n_440),
.B2(n_431),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_488),
.A2(n_505),
.B1(n_513),
.B2(n_480),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_417),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_489),
.B(n_501),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_490),
.A2(n_392),
.B(n_359),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_480),
.Y(n_493)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_493),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_456),
.A2(n_431),
.B1(n_416),
.B2(n_441),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_494),
.A2(n_500),
.B1(n_507),
.B2(n_512),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_508),
.C(n_510),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_452),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_498),
.B(n_504),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_458),
.B(n_436),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_350),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_455),
.A2(n_420),
.B1(n_412),
.B2(n_421),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_459),
.A2(n_420),
.B1(n_421),
.B2(n_436),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_458),
.B(n_340),
.C(n_445),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_470),
.A2(n_445),
.B1(n_435),
.B2(n_433),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_451),
.B(n_340),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_454),
.B(n_356),
.C(n_435),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_514),
.C(n_515),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_471),
.A2(n_433),
.B1(n_342),
.B2(n_351),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_462),
.A2(n_439),
.B1(n_303),
.B2(n_351),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_451),
.B(n_316),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_474),
.B(n_316),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_483),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_516),
.B(n_529),
.Y(n_554)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_493),
.Y(n_517)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_517),
.Y(n_545)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_518),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_486),
.B(n_467),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_520),
.B(n_522),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_484),
.B(n_481),
.Y(n_521)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_521),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_510),
.B(n_477),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_483),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_523),
.B(n_533),
.Y(n_559)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_492),
.Y(n_526)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_526),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_R g527 ( 
.A(n_497),
.B(n_453),
.Y(n_527)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_527),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_514),
.B(n_472),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_469),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_531),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_489),
.B(n_448),
.C(n_464),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_532),
.B(n_539),
.Y(n_561)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_495),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_534),
.B(n_536),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_485),
.B(n_469),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_543),
.Y(n_550)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_502),
.Y(n_536)
);

NAND2x1_ASAP7_75t_L g537 ( 
.A(n_491),
.B(n_468),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_537),
.B(n_505),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_494),
.A2(n_457),
.B1(n_449),
.B2(n_460),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_538),
.A2(n_530),
.B1(n_482),
.B2(n_523),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_485),
.B(n_387),
.C(n_309),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g548 ( 
.A1(n_540),
.A2(n_491),
.B1(n_488),
.B2(n_512),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_309),
.C(n_356),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_541),
.B(n_544),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_300),
.C(n_338),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_548),
.Y(n_585)
);

FAx1_ASAP7_75t_SL g549 ( 
.A(n_527),
.B(n_496),
.CI(n_490),
.CON(n_549),
.SN(n_549)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_549),
.B(n_525),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_499),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_555),
.Y(n_583)
);

INVxp33_ASAP7_75t_SL g552 ( 
.A(n_534),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_552),
.A2(n_563),
.B(n_554),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_528),
.B(n_499),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_528),
.B(n_501),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_556),
.B(n_565),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_SL g558 ( 
.A(n_532),
.B(n_515),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_558),
.B(n_521),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_525),
.B(n_482),
.Y(n_565)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_566),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_567),
.A2(n_540),
.B1(n_531),
.B2(n_530),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_568),
.A2(n_547),
.B1(n_546),
.B2(n_559),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_551),
.B(n_524),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_570),
.B(n_576),
.Y(n_587)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_563),
.Y(n_571)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_571),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_553),
.B(n_519),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_575),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_558),
.B(n_550),
.Y(n_573)
);

XNOR2x1_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_577),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_574),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_555),
.B(n_524),
.C(n_539),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_550),
.B(n_565),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_556),
.B(n_544),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_561),
.B(n_541),
.C(n_538),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_557),
.C(n_566),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_579),
.B(n_580),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_SL g580 ( 
.A(n_549),
.B(n_537),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_581),
.A2(n_564),
.B(n_578),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_SL g582 ( 
.A(n_549),
.B(n_537),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_582),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_562),
.B(n_542),
.Y(n_586)
);

INVx11_ASAP7_75t_L g595 ( 
.A(n_586),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_585),
.A2(n_557),
.B1(n_569),
.B2(n_567),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_588),
.B(n_598),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_589),
.B(n_600),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_590),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_592),
.A2(n_526),
.B1(n_582),
.B2(n_502),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_585),
.A2(n_559),
.B(n_543),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_575),
.B(n_513),
.C(n_545),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_545),
.C(n_560),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_601),
.B(n_303),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_580),
.A2(n_536),
.B(n_533),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_602),
.A2(n_506),
.B(n_503),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_583),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_605),
.B(n_607),
.Y(n_623)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_606),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_587),
.B(n_601),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_596),
.A2(n_570),
.B(n_579),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_608),
.B(n_611),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_576),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_SL g617 ( 
.A(n_609),
.B(n_610),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_584),
.C(n_573),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_517),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_595),
.B(n_542),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_592),
.Y(n_619)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_614),
.Y(n_621)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_615),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_613),
.A2(n_595),
.B(n_602),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_616),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_619),
.B(n_594),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_603),
.B(n_604),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_622),
.B(n_591),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_607),
.B(n_597),
.C(n_591),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_624),
.B(n_609),
.C(n_610),
.Y(n_630)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_628),
.C(n_629),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_623),
.B(n_605),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_630),
.A2(n_617),
.B(n_624),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_613),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_L g634 ( 
.A(n_631),
.B(n_618),
.C(n_625),
.Y(n_634)
);

OAI221xp5_ASAP7_75t_L g636 ( 
.A1(n_632),
.A2(n_634),
.B1(n_620),
.B2(n_598),
.C(n_599),
.Y(n_636)
);

NAND4xp25_ASAP7_75t_L g635 ( 
.A(n_627),
.B(n_630),
.C(n_621),
.D(n_614),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_635),
.A2(n_633),
.B(n_597),
.Y(n_637)
);

OAI321xp33_ASAP7_75t_L g638 ( 
.A1(n_636),
.A2(n_637),
.A3(n_593),
.B1(n_392),
.B2(n_359),
.C(n_305),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_638),
.A2(n_300),
.B(n_392),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_639),
.B(n_318),
.C(n_593),
.Y(n_640)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_640),
.B(n_318),
.Y(n_641)
);


endmodule