module real_jpeg_24237_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_70;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_60),
.Y(n_123)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_6),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_74),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_8),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_9),
.A2(n_26),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_9),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_9),
.A2(n_26),
.B1(n_51),
.B2(n_52),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_10),
.B(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_10),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_10),
.B(n_51),
.C(n_65),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_10),
.B(n_117),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_10),
.A2(n_58),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_71),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_71),
.Y(n_144)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_15),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_20),
.B(n_87),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.C(n_76),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_21),
.A2(n_22),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_23),
.B(n_42),
.C(n_61),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_32),
.B2(n_38),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_25),
.A2(n_31),
.B1(n_79),
.B2(n_117),
.Y(n_181)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_27),
.B(n_80),
.CON(n_79),
.SN(n_79)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_34),
.C(n_36),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_27),
.A2(n_46),
.B(n_92),
.C(n_95),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_47),
.C(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_31),
.A2(n_39),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_33),
.A2(n_35),
.B(n_79),
.C(n_81),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_34),
.A2(n_35),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_35),
.B(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_61),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_44),
.A2(n_92),
.B1(n_103),
.B2(n_108),
.Y(n_102)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_45),
.B(n_104),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_46),
.A2(n_47),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_53),
.B(n_57),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_49),
.Y(n_97)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_56),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_52),
.B1(n_65),
.B2(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_52),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_53),
.B(n_84),
.Y(n_145)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_59),
.Y(n_86)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_56),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_58),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_58),
.A2(n_100),
.B1(n_150),
.B2(n_159),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_62),
.A2(n_76),
.B1(n_77),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_62),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_69),
.B(n_72),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_63),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_63),
.A2(n_68),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_63),
.A2(n_68),
.B1(n_135),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_68),
.B(n_80),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_70),
.A2(n_75),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_75),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_78),
.A2(n_82),
.B1(n_83),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

HAxp5_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_93),
.CON(n_92),
.SN(n_92)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_80),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_85),
.A2(n_149),
.B1(n_151),
.B2(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_184),
.B(n_190),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_173),
.B(n_183),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_146),
.B(n_172),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_132),
.B1(n_133),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_182)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_144),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_156),
.B(n_171),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_154),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_167),
.B(n_170),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_163),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_168),
.B(n_169),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_182),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_178),
.C(n_181),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);


endmodule