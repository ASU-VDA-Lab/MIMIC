module fake_jpeg_10329_n_143 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_32),
.Y(n_37)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_43),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_15),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_14),
.B1(n_20),
.B2(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_49),
.B1(n_19),
.B2(n_18),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_14),
.B1(n_26),
.B2(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_56),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_36),
.B1(n_29),
.B2(n_32),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_59),
.B1(n_23),
.B2(n_18),
.Y(n_71)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_32),
.B1(n_29),
.B2(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_50),
.B1(n_37),
.B2(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_43),
.B1(n_37),
.B2(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_72),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_63),
.B1(n_26),
.B2(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_76),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_41),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_47),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_49),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_89),
.B1(n_23),
.B2(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_67),
.B(n_78),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_92),
.B(n_35),
.C(n_10),
.D(n_9),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_82),
.C(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_100),
.Y(n_107)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_72),
.A3(n_65),
.B1(n_92),
.B2(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

OAI321xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_94),
.A3(n_98),
.B1(n_96),
.B2(n_95),
.C(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_113),
.Y(n_116)
);

AOI22x1_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_88),
.B1(n_87),
.B2(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_109),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_8),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_99),
.B1(n_75),
.B2(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_56),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_19),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_119),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_54),
.Y(n_120)
);

OA21x2_ASAP7_75t_SL g123 ( 
.A1(n_120),
.A2(n_111),
.B(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_75),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_122),
.C(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_0),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_127),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_35),
.C(n_31),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_31),
.C(n_30),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_121),
.B1(n_7),
.B2(n_8),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_131),
.A2(n_132),
.B1(n_0),
.B2(n_1),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_135),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_129),
.B(n_1),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_30),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_137),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C(n_30),
.Y(n_139)
);

OAI21x1_ASAP7_75t_SL g141 ( 
.A1(n_139),
.A2(n_134),
.B(n_4),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_141),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_31),
.Y(n_143)
);


endmodule