module fake_jpeg_159_n_685 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_685);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_685;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_59),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_65),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_66),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_69),
.B(n_80),
.Y(n_136)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_70),
.Y(n_199)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_73),
.Y(n_200)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_74),
.Y(n_204)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_77),
.Y(n_197)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_78),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_19),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_81),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_82),
.Y(n_206)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_18),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_106),
.Y(n_139)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_86),
.Y(n_228)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_87),
.Y(n_231)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_89),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_25),
.Y(n_90)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_90),
.Y(n_191)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_92),
.Y(n_195)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_93),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_97),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_103),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_104),
.Y(n_223)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_26),
.B(n_18),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_107),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_27),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_108),
.B(n_117),
.Y(n_164)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_26),
.B(n_17),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_129),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_30),
.Y(n_116)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_41),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_27),
.Y(n_120)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

CKINVDCx6p67_ASAP7_75t_R g178 ( 
.A(n_121),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_44),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_43),
.B(n_16),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_35),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_43),
.B(n_16),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_13),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_54),
.B1(n_56),
.B2(n_24),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_134),
.A2(n_145),
.B1(n_161),
.B2(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_138),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_35),
.B1(n_38),
.B2(n_54),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_28),
.C(n_53),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_147),
.B(n_42),
.C(n_55),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_24),
.B1(n_30),
.B2(n_33),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_150),
.A2(n_153),
.B1(n_160),
.B2(n_171),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_35),
.B1(n_38),
.B2(n_53),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_60),
.A2(n_44),
.B1(n_24),
.B2(n_56),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_65),
.A2(n_83),
.B1(n_92),
.B2(n_89),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_166),
.B(n_214),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_99),
.A2(n_57),
.B1(n_23),
.B2(n_52),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_88),
.Y(n_176)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_109),
.A2(n_57),
.B1(n_23),
.B2(n_52),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_179),
.A2(n_193),
.B1(n_212),
.B2(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_70),
.Y(n_182)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_182),
.Y(n_273)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_81),
.Y(n_183)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_183),
.Y(n_296)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_73),
.Y(n_189)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_189),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_74),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_192),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_64),
.A2(n_39),
.B1(n_28),
.B2(n_32),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_128),
.B(n_46),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_194),
.B(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_196),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_66),
.A2(n_38),
.B1(n_32),
.B2(n_46),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_98),
.A2(n_123),
.B1(n_121),
.B2(n_57),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_126),
.A2(n_52),
.B1(n_23),
.B2(n_39),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_67),
.B(n_15),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_77),
.B(n_15),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_79),
.B(n_15),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_2),
.C(n_4),
.Y(n_283)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_82),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_217),
.B(n_227),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_118),
.B(n_13),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_94),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_100),
.B(n_13),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_104),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_230),
.B(n_210),
.Y(n_316)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_232),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_235),
.Y(n_363)
);

BUFx2_ASAP7_75t_SL g237 ( 
.A(n_178),
.Y(n_237)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_237),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_151),
.Y(n_238)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_238),
.Y(n_328)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_243),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_0),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_244),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_245),
.B(n_275),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_134),
.A2(n_115),
.B1(n_55),
.B2(n_42),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_250),
.A2(n_278),
.B1(n_300),
.B2(n_312),
.Y(n_346)
);

BUFx12f_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

NAND2xp33_ASAP7_75t_R g252 ( 
.A(n_139),
.B(n_42),
.Y(n_252)
);

OR2x2_ASAP7_75t_SL g373 ( 
.A(n_252),
.B(n_259),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_140),
.A2(n_55),
.B1(n_12),
.B2(n_11),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_253),
.A2(n_269),
.B1(n_271),
.B2(n_287),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_155),
.B(n_12),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_254),
.B(n_256),
.Y(n_334)
);

AND2x2_ASAP7_75t_SL g255 ( 
.A(n_133),
.B(n_55),
.Y(n_255)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_255),
.B(n_299),
.C(n_190),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_136),
.B(n_11),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_137),
.B(n_0),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_257),
.B(n_266),
.Y(n_380)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_258),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_142),
.B(n_55),
.C(n_1),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_259),
.B(n_265),
.C(n_255),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_192),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_260),
.B(n_284),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_164),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_261),
.B(n_283),
.Y(n_355)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_262),
.Y(n_343)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_263),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_148),
.B(n_55),
.C(n_1),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_152),
.B(n_0),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_267),
.Y(n_370)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_140),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_270),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_160),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_135),
.Y(n_272)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_274),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_149),
.B(n_8),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_218),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_276),
.Y(n_356)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_132),
.Y(n_277)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_277),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_172),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_151),
.Y(n_280)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_280),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_168),
.Y(n_281)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_281),
.Y(n_366)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_205),
.Y(n_282)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_282),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_200),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_285),
.Y(n_371)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_228),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_288),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_212),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_198),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_220),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_289),
.A2(n_318),
.B1(n_220),
.B2(n_159),
.Y(n_341)
);

BUFx4f_ASAP7_75t_L g290 ( 
.A(n_211),
.Y(n_290)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_290),
.Y(n_379)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_184),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_292),
.Y(n_336)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_187),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_200),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_295),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_168),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_294),
.A2(n_315),
.B(n_150),
.Y(n_319)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_185),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_174),
.B(n_8),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_298),
.Y(n_344)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_185),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g299 ( 
.A(n_154),
.B(n_6),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_175),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_167),
.B(n_169),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_301),
.B(n_302),
.Y(n_345)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_141),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_188),
.B(n_7),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_303),
.B(n_304),
.Y(n_375)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_162),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_177),
.A2(n_8),
.B1(n_219),
.B2(n_226),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_305),
.A2(n_310),
.B1(n_271),
.B2(n_253),
.Y(n_327)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_207),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_306),
.Y(n_359)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_177),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_307),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_198),
.B(n_143),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_309),
.Y(n_325)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_219),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_213),
.A2(n_8),
.B1(n_210),
.B2(n_195),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_204),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_314),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_170),
.A2(n_181),
.B1(n_180),
.B2(n_158),
.Y(n_312)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_162),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_144),
.A2(n_225),
.B1(n_204),
.B2(n_224),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_223),
.Y(n_331)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_163),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

AND2x4_ASAP7_75t_SL g320 ( 
.A(n_240),
.B(n_224),
.Y(n_320)
);

BUFx8_ASAP7_75t_L g415 ( 
.A(n_320),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_241),
.B(n_199),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_323),
.B(n_319),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_239),
.A2(n_226),
.B1(n_206),
.B2(n_163),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_324),
.A2(n_327),
.B1(n_341),
.B2(n_342),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_331),
.B(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_332),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_179),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_338),
.B(n_347),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_234),
.A2(n_206),
.B1(n_186),
.B2(n_190),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_299),
.B(n_195),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_248),
.B(n_275),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_358),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_234),
.A2(n_186),
.B1(n_197),
.B2(n_202),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_351),
.A2(n_377),
.B1(n_381),
.B2(n_251),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_245),
.B(n_171),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_369),
.C(n_244),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_275),
.B(n_223),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_240),
.A2(n_197),
.B1(n_202),
.B2(n_146),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_361),
.A2(n_263),
.B(n_288),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_246),
.B(n_146),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_376),
.Y(n_413)
);

AOI21xp33_ASAP7_75t_L g405 ( 
.A1(n_373),
.A2(n_295),
.B(n_298),
.Y(n_405)
);

AND2x4_ASAP7_75t_SL g374 ( 
.A(n_310),
.B(n_255),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_374),
.B(n_361),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_265),
.B(n_244),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_242),
.A2(n_236),
.B1(n_264),
.B2(n_306),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_262),
.A2(n_268),
.B1(n_233),
.B2(n_309),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_325),
.Y(n_382)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_383),
.B(n_421),
.C(n_426),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_313),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_384),
.Y(n_464)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_273),
.C(n_296),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_386),
.B(n_392),
.C(n_395),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_342),
.A2(n_305),
.B1(n_294),
.B2(n_269),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_387),
.A2(n_388),
.B1(n_389),
.B2(n_412),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_351),
.A2(n_315),
.B1(n_307),
.B2(n_258),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_327),
.A2(n_321),
.B1(n_338),
.B2(n_365),
.Y(n_389)
);

AOI22x1_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_274),
.B1(n_302),
.B2(n_282),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_390),
.A2(n_408),
.B1(n_410),
.B2(n_417),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_349),
.B(n_317),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_323),
.B(n_247),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_394),
.B(n_402),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_249),
.C(n_272),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_380),
.B(n_291),
.Y(n_396)
);

NOR3xp33_ASAP7_75t_L g439 ( 
.A(n_396),
.B(n_405),
.C(n_415),
.Y(n_439)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_399),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_400),
.Y(n_437)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_336),
.Y(n_401)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_401),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_286),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_403),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_326),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_411),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_352),
.A2(n_304),
.B(n_314),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_406),
.A2(n_363),
.B(n_343),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_374),
.A2(n_232),
.B1(n_292),
.B2(n_279),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_344),
.B(n_235),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_423),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_374),
.A2(n_280),
.B1(n_318),
.B2(n_238),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_270),
.Y(n_411)
);

INVx5_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_321),
.A2(n_285),
.B1(n_251),
.B2(n_267),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_416),
.A2(n_368),
.B1(n_378),
.B2(n_339),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_346),
.A2(n_290),
.B1(n_311),
.B2(n_243),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_418),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_347),
.A2(n_320),
.B1(n_375),
.B2(n_353),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_422),
.B1(n_339),
.B2(n_359),
.Y(n_452)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_420),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_372),
.B(n_332),
.C(n_376),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_320),
.A2(n_290),
.B1(n_281),
.B2(n_277),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_332),
.B(n_345),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_358),
.B(n_331),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_356),
.Y(n_440)
);

MAJx2_ASAP7_75t_L g426 ( 
.A(n_373),
.B(n_334),
.C(n_320),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

BUFx5_ASAP7_75t_L g468 ( 
.A(n_427),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_428),
.B(n_392),
.Y(n_456)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_431),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_430),
.A2(n_339),
.B(n_362),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_354),
.Y(n_431)
);

AOI322xp5_ASAP7_75t_L g432 ( 
.A1(n_423),
.A2(n_330),
.A3(n_341),
.B1(n_362),
.B2(n_356),
.C1(n_334),
.C2(n_378),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g496 ( 
.A(n_432),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_414),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_434),
.B(n_440),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_439),
.Y(n_514)
);

AOI22x1_ASAP7_75t_SL g442 ( 
.A1(n_415),
.A2(n_368),
.B1(n_333),
.B2(n_366),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_442),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_444),
.A2(n_449),
.B1(n_452),
.B2(n_458),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_397),
.A2(n_366),
.B(n_333),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_448),
.A2(n_470),
.B(n_457),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_430),
.A2(n_398),
.B1(n_382),
.B2(n_385),
.Y(n_449)
);

OAI32xp33_ASAP7_75t_L g451 ( 
.A1(n_398),
.A2(n_360),
.A3(n_367),
.B1(n_322),
.B2(n_371),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_451),
.B(n_459),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_409),
.Y(n_454)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_454),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_455),
.A2(n_461),
.B(n_465),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_456),
.B(n_453),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_415),
.Y(n_457)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_389),
.A2(n_364),
.B1(n_328),
.B2(n_359),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_367),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_431),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_429),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_397),
.A2(n_415),
.B(n_419),
.Y(n_461)
);

AO22x1_ASAP7_75t_SL g462 ( 
.A1(n_387),
.A2(n_360),
.B1(n_364),
.B2(n_371),
.Y(n_462)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_393),
.A2(n_357),
.B1(n_370),
.B2(n_354),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_463),
.A2(n_467),
.B1(n_410),
.B2(n_422),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_413),
.A2(n_329),
.B(n_350),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_393),
.A2(n_357),
.B1(n_370),
.B2(n_350),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_471),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_476),
.B(n_478),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_471),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_421),
.C(n_413),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_479),
.B(n_481),
.C(n_489),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_435),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_440),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_482),
.B(n_502),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_461),
.A2(n_390),
.B(n_400),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_485),
.A2(n_448),
.B(n_442),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_441),
.A2(n_416),
.B1(n_412),
.B2(n_406),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_486),
.A2(n_492),
.B1(n_495),
.B2(n_504),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_487),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_450),
.B(n_383),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_490),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g531 ( 
.A1(n_491),
.A2(n_462),
.B(n_442),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_441),
.A2(n_399),
.B1(n_425),
.B2(n_401),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_469),
.Y(n_493)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_493),
.Y(n_527)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_494),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_458),
.A2(n_425),
.B1(n_394),
.B2(n_388),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_433),
.A2(n_428),
.B1(n_408),
.B2(n_407),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_498),
.A2(n_452),
.B1(n_466),
.B2(n_464),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_454),
.B(n_407),
.Y(n_499)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_499),
.Y(n_539)
);

FAx1_ASAP7_75t_SL g500 ( 
.A(n_449),
.B(n_426),
.CI(n_386),
.CON(n_500),
.SN(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_500),
.A2(n_456),
.B(n_445),
.C(n_455),
.Y(n_517)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_501),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_433),
.B(n_443),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_459),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_503),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_443),
.A2(n_390),
.B1(n_396),
.B2(n_395),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_465),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_505),
.B(n_507),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_435),
.B(n_426),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_448),
.C(n_447),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_438),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_508),
.B(n_453),
.Y(n_515)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_468),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_509),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_510),
.Y(n_534)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_451),
.Y(n_511)
);

NAND2x1_ASAP7_75t_SL g528 ( 
.A(n_511),
.B(n_462),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_438),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_513),
.A2(n_403),
.B1(n_420),
.B2(n_472),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_515),
.B(n_521),
.Y(n_556)
);

AOI21xp33_ASAP7_75t_L g572 ( 
.A1(n_517),
.A2(n_500),
.B(n_496),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_475),
.A2(n_467),
.B1(n_463),
.B2(n_437),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_519),
.A2(n_538),
.B1(n_544),
.B2(n_546),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_524),
.B1(n_535),
.B2(n_540),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_446),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_475),
.A2(n_436),
.B1(n_446),
.B2(n_445),
.Y(n_524)
);

NAND2x1_ASAP7_75t_L g525 ( 
.A(n_488),
.B(n_470),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_525),
.A2(n_529),
.B(n_487),
.Y(n_554)
);

OA22x2_ASAP7_75t_L g526 ( 
.A1(n_511),
.A2(n_444),
.B1(n_462),
.B2(n_436),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_526),
.B(n_484),
.Y(n_555)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_528),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_530),
.B(n_532),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_531),
.A2(n_484),
.B1(n_505),
.B2(n_486),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_489),
.B(n_466),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_483),
.A2(n_460),
.B1(n_434),
.B2(n_473),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_492),
.A2(n_432),
.B1(n_473),
.B2(n_472),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_479),
.B(n_481),
.C(n_506),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_541),
.B(n_548),
.C(n_552),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_512),
.A2(n_418),
.B1(n_328),
.B2(n_427),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_512),
.A2(n_328),
.B1(n_468),
.B2(n_348),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_497),
.A2(n_343),
.B(n_348),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_547),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_498),
.B(n_335),
.C(n_379),
.Y(n_548)
);

AOI32xp33_ASAP7_75t_L g549 ( 
.A1(n_514),
.A2(n_335),
.A3(n_379),
.B1(n_513),
.B2(n_507),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_480),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_483),
.A2(n_379),
.B1(n_482),
.B2(n_488),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_550),
.A2(n_477),
.B1(n_485),
.B2(n_480),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_499),
.B(n_503),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_SL g600 ( 
.A1(n_554),
.A2(n_526),
.B(n_537),
.Y(n_600)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_555),
.Y(n_598)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_557),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_502),
.Y(n_558)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_559),
.A2(n_569),
.B1(n_531),
.B2(n_529),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_534),
.B(n_476),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_573),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_532),
.B(n_497),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_565),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_495),
.C(n_478),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_570),
.C(n_576),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_521),
.B(n_504),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_542),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_566),
.B(n_575),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_518),
.B(n_515),
.C(n_541),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_520),
.B(n_477),
.Y(n_571)
);

CKINVDCx14_ASAP7_75t_R g601 ( 
.A(n_571),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_572),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_490),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_574),
.B(n_581),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_524),
.A2(n_536),
.B1(n_531),
.B2(n_516),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_530),
.B(n_517),
.C(n_551),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_538),
.A2(n_491),
.B1(n_493),
.B2(n_494),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_577),
.A2(n_582),
.B1(n_531),
.B2(n_526),
.Y(n_597)
);

CKINVDCx14_ASAP7_75t_R g578 ( 
.A(n_516),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_578),
.B(n_579),
.Y(n_603)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_543),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_542),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_580),
.Y(n_592)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_537),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_531),
.A2(n_519),
.B1(n_550),
.B2(n_544),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_547),
.Y(n_585)
);

MAJx2_ASAP7_75t_L g619 ( 
.A(n_585),
.B(n_586),
.C(n_594),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_553),
.B(n_552),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_564),
.B(n_545),
.C(n_548),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_590),
.B(n_591),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_570),
.B(n_545),
.C(n_535),
.Y(n_591)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_593),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_583),
.B(n_525),
.Y(n_594)
);

XNOR2x1_ASAP7_75t_L g595 ( 
.A(n_563),
.B(n_525),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_595),
.B(n_565),
.Y(n_610)
);

FAx1_ASAP7_75t_SL g596 ( 
.A(n_576),
.B(n_500),
.CI(n_528),
.CON(n_596),
.SN(n_596)
);

AOI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_596),
.A2(n_597),
.B1(n_598),
.B2(n_588),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_600),
.A2(n_555),
.B(n_559),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_583),
.B(n_546),
.C(n_526),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_606),
.C(n_609),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_556),
.B(n_523),
.C(n_501),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_562),
.A2(n_523),
.B1(n_522),
.B2(n_527),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g621 ( 
.A1(n_607),
.A2(n_567),
.B1(n_577),
.B2(n_582),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_556),
.B(n_533),
.C(n_509),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_610),
.B(n_613),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_586),
.B(n_568),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_612),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_554),
.Y(n_613)
);

INVx11_ASAP7_75t_L g614 ( 
.A(n_601),
.Y(n_614)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_614),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_587),
.B(n_568),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_616),
.B(n_622),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_589),
.B(n_561),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_617),
.B(n_599),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_618),
.A2(n_588),
.B(n_597),
.Y(n_644)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_621),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_584),
.B(n_560),
.C(n_580),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_602),
.A2(n_567),
.B1(n_579),
.B2(n_560),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_623),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_584),
.B(n_557),
.C(n_566),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_624),
.B(n_628),
.C(n_599),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_606),
.B(n_558),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_625),
.B(n_627),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_602),
.A2(n_581),
.B(n_608),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_626),
.B(n_595),
.Y(n_641)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_603),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_591),
.B(n_590),
.C(n_585),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g629 ( 
.A(n_609),
.B(n_594),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_629),
.B(n_592),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g638 ( 
.A1(n_630),
.A2(n_600),
.B(n_593),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_634),
.B(n_612),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_615),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_618),
.A2(n_598),
.B(n_604),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_639),
.A2(n_641),
.B(n_644),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_622),
.B(n_607),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_640),
.B(n_643),
.Y(n_657)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_642),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_628),
.B(n_624),
.C(n_611),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_645),
.B(n_648),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_630),
.A2(n_605),
.B(n_596),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_646),
.A2(n_613),
.B(n_610),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_620),
.B(n_596),
.C(n_625),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_643),
.B(n_645),
.C(n_620),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_649),
.B(n_651),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_648),
.B(n_623),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_636),
.B(n_629),
.C(n_615),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_652),
.B(n_659),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_654),
.B(n_656),
.Y(n_666)
);

XOR2xp5_ASAP7_75t_L g665 ( 
.A(n_658),
.B(n_646),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_633),
.B(n_621),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_635),
.A2(n_614),
.B1(n_616),
.B2(n_619),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_660),
.A2(n_661),
.B1(n_641),
.B2(n_637),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_632),
.B(n_619),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_649),
.B(n_642),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_662),
.B(n_664),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_652),
.B(n_635),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_665),
.B(n_667),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_657),
.B(n_631),
.C(n_644),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_669),
.B(n_663),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_650),
.B(n_647),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_SL g671 ( 
.A(n_670),
.B(n_661),
.Y(n_671)
);

NOR3xp33_ASAP7_75t_L g678 ( 
.A(n_671),
.B(n_675),
.C(n_655),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g677 ( 
.A(n_673),
.B(n_674),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_668),
.B(n_653),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_669),
.B(n_655),
.C(n_656),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_678),
.A2(n_676),
.B(n_666),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_672),
.B(n_665),
.C(n_632),
.Y(n_679)
);

AOI21x1_ASAP7_75t_L g681 ( 
.A1(n_679),
.A2(n_666),
.B(n_639),
.Y(n_681)
);

BUFx24_ASAP7_75t_SL g682 ( 
.A(n_680),
.Y(n_682)
);

MAJx2_ASAP7_75t_L g683 ( 
.A(n_682),
.B(n_681),
.C(n_677),
.Y(n_683)
);

OAI321xp33_ASAP7_75t_L g684 ( 
.A1(n_683),
.A2(n_658),
.A3(n_637),
.B1(n_660),
.B2(n_638),
.C(n_647),
.Y(n_684)
);

BUFx24_ASAP7_75t_SL g685 ( 
.A(n_684),
.Y(n_685)
);


endmodule