module real_aes_7691_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_56;
wire n_34;
wire n_55;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_33;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_51;
wire n_54;
wire n_35;
wire n_42;
wire n_45;
wire n_39;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_52;
wire n_57;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_53;
wire n_36;
NOR2xp33_ASAP7_75t_R g22 ( .A(n_0), .B(n_23), .Y(n_22) );
CKINVDCx20_ASAP7_75t_R g38 ( .A(n_0), .Y(n_38) );
NAND2xp33_ASAP7_75t_SL g52 ( .A(n_0), .B(n_53), .Y(n_52) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_1), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g37 ( .A(n_1), .B(n_15), .Y(n_37) );
NOR2xp33_ASAP7_75t_R g42 ( .A(n_1), .B(n_43), .Y(n_42) );
NAND2xp33_ASAP7_75t_SL g46 ( .A(n_1), .B(n_19), .Y(n_46) );
NAND2xp33_ASAP7_75t_SL g56 ( .A(n_1), .B(n_44), .Y(n_56) );
CKINVDCx20_ASAP7_75t_R g28 ( .A(n_2), .Y(n_28) );
NOR3xp33_ASAP7_75t_SL g26 ( .A(n_3), .B(n_11), .C(n_27), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_4), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g20 ( .A(n_5), .Y(n_20) );
NAND2xp33_ASAP7_75t_SL g33 ( .A(n_5), .B(n_34), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g44 ( .A(n_5), .B(n_21), .Y(n_44) );
CKINVDCx20_ASAP7_75t_R g55 ( .A(n_6), .Y(n_55) );
CKINVDCx20_ASAP7_75t_R g57 ( .A(n_7), .Y(n_57) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_8), .Y(n_27) );
AOI221xp5_ASAP7_75t_SL g39 ( .A1(n_9), .A2(n_13), .B1(n_40), .B2(n_45), .C(n_47), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_10), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g24 ( .A(n_12), .Y(n_24) );
NOR4xp25_ASAP7_75t_SL g32 ( .A(n_12), .B(n_33), .C(n_36), .D(n_38), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g49 ( .A(n_12), .B(n_50), .Y(n_49) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_14), .Y(n_23) );
NAND4xp25_ASAP7_75t_SL g21 ( .A(n_15), .B(n_22), .C(n_24), .D(n_25), .Y(n_21) );
OAI221xp5_ASAP7_75t_R g16 ( .A1(n_17), .A2(n_18), .B1(n_30), .B2(n_31), .C(n_39), .Y(n_16) );
NAND2xp33_ASAP7_75t_SL g18 ( .A(n_19), .B(n_29), .Y(n_18) );
NOR2xp33_ASAP7_75t_R g19 ( .A(n_20), .B(n_21), .Y(n_19) );
NAND2xp33_ASAP7_75t_SL g54 ( .A(n_20), .B(n_34), .Y(n_54) );
NAND2xp33_ASAP7_75t_SL g35 ( .A(n_23), .B(n_25), .Y(n_35) );
AND2x2_ASAP7_75t_L g25 ( .A(n_26), .B(n_28), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_32), .Y(n_31) );
CKINVDCx20_ASAP7_75t_R g34 ( .A(n_35), .Y(n_34) );
CKINVDCx20_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
NAND2xp33_ASAP7_75t_SL g50 ( .A(n_37), .B(n_51), .Y(n_50) );
CKINVDCx20_ASAP7_75t_R g40 ( .A(n_41), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_42), .Y(n_41) );
CKINVDCx16_ASAP7_75t_R g43 ( .A(n_44), .Y(n_43) );
INVx1_ASAP7_75t_SL g45 ( .A(n_46), .Y(n_45) );
OAI22xp33_ASAP7_75t_SL g47 ( .A1(n_48), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_47) );
CKINVDCx16_ASAP7_75t_R g48 ( .A(n_49), .Y(n_48) );
CKINVDCx5p33_ASAP7_75t_R g51 ( .A(n_52), .Y(n_51) );
CKINVDCx20_ASAP7_75t_R g53 ( .A(n_54), .Y(n_53) );
endmodule