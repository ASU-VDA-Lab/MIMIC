module fake_jpeg_16700_n_358 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_358);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_23),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_24),
.B1(n_38),
.B2(n_21),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_76),
.B1(n_27),
.B2(n_32),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_24),
.B1(n_22),
.B2(n_21),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_83),
.B1(n_35),
.B2(n_29),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_67),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_33),
.B(n_19),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_22),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_29),
.B1(n_38),
.B2(n_31),
.Y(n_76)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NAND2x1p5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_59),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_86),
.A2(n_90),
.B1(n_108),
.B2(n_37),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_47),
.B1(n_35),
.B2(n_27),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_27),
.B1(n_26),
.B2(n_32),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_25),
.B1(n_32),
.B2(n_26),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_104),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_25),
.B1(n_35),
.B2(n_31),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_102),
.Y(n_139)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_57),
.B1(n_68),
.B2(n_80),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_61),
.B1(n_72),
.B2(n_48),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_57),
.B1(n_68),
.B2(n_80),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_74),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_48),
.B1(n_37),
.B2(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_56),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_41),
.Y(n_116)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

OAI21x1_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_91),
.B(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_122),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_107),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_71),
.B1(n_51),
.B2(n_56),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_110),
.B1(n_114),
.B2(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_77),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_53),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_140),
.B(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_53),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_100),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_143),
.B(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_100),
.B(n_71),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_100),
.B(n_52),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_52),
.B1(n_51),
.B2(n_45),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_97),
.B1(n_104),
.B2(n_93),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_123),
.B(n_133),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_153),
.B(n_157),
.Y(n_172)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_93),
.B1(n_105),
.B2(n_109),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_103),
.B1(n_42),
.B2(n_45),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_42),
.B1(n_103),
.B2(n_36),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_160),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_63),
.C(n_37),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_133),
.C(n_142),
.Y(n_182)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_118),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_170),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_176),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_150),
.B(n_133),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_185),
.C(n_190),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_196),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_116),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_134),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_115),
.C(n_143),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_129),
.B(n_138),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_148),
.B(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_136),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_136),
.B(n_121),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_195),
.B(n_171),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_117),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_121),
.B(n_117),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_198),
.B1(n_203),
.B2(n_208),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_165),
.B1(n_148),
.B2(n_160),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_179),
.A2(n_165),
.B1(n_159),
.B2(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_220),
.B1(n_222),
.B2(n_181),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_155),
.B(n_168),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_185),
.C(n_182),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_207),
.C(n_182),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_157),
.B1(n_152),
.B2(n_146),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_192),
.B1(n_194),
.B2(n_175),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_120),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_170),
.B1(n_164),
.B2(n_126),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_164),
.B(n_141),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_213),
.B1(n_216),
.B2(n_219),
.Y(n_239)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_180),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_193),
.A2(n_37),
.B(n_34),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_187),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_141),
.B(n_34),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_145),
.B1(n_126),
.B2(n_141),
.Y(n_216)
);

NAND2x1_ASAP7_75t_SL g218 ( 
.A(n_172),
.B(n_34),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_196),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_141),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_34),
.B(n_1),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_172),
.B1(n_190),
.B2(n_189),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_215),
.B(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_227),
.B(n_238),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_214),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_241),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_197),
.B1(n_216),
.B2(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_217),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_235),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_211),
.B(n_248),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_184),
.C(n_178),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_198),
.A2(n_173),
.B1(n_184),
.B2(n_180),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_240),
.A2(n_242),
.B1(n_247),
.B2(n_220),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_202),
.B(n_39),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_37),
.C(n_36),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_213),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_0),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_39),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_222),
.A3(n_201),
.B1(n_203),
.B2(n_199),
.C1(n_207),
.C2(n_200),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_255),
.Y(n_290)
);

BUFx4f_ASAP7_75t_SL g253 ( 
.A(n_230),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_243),
.C(n_231),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_218),
.B1(n_209),
.B2(n_205),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_246),
.B1(n_234),
.B2(n_236),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_265),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_239),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_218),
.B1(n_17),
.B2(n_36),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_232),
.C(n_224),
.Y(n_272)
);

XOR2x2_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_259),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_238),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_275),
.C(n_276),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_277),
.B(n_265),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_246),
.B1(n_247),
.B2(n_229),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_278),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_241),
.B1(n_235),
.B2(n_7),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_5),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_286),
.C(n_291),
.Y(n_300)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_34),
.C(n_8),
.Y(n_286)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_253),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_269),
.B1(n_268),
.B2(n_267),
.Y(n_303)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_8),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_254),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_292),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_280),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_293),
.A2(n_304),
.B1(n_286),
.B2(n_287),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_303),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_272),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_290),
.A2(n_279),
.B(n_274),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_282),
.B(n_275),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_252),
.B(n_250),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_249),
.C(n_260),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_306),
.C(n_288),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_252),
.C(n_10),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_306),
.C(n_296),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_321),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_320),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_299),
.B(n_305),
.CI(n_300),
.CON(n_315),
.SN(n_315)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_315),
.B(n_316),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_9),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_298),
.B1(n_292),
.B2(n_14),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_307),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_292),
.A2(n_10),
.B(n_12),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_333),
.C(n_318),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_325),
.B(n_329),
.Y(n_341)
);

OA21x2_ASAP7_75t_SL g326 ( 
.A1(n_315),
.A2(n_300),
.B(n_296),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_326),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_16),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_16),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_316),
.C(n_309),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_328),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_329),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_339),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_317),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_340),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_319),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_12),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_341),
.B(n_342),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_13),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_333),
.B(n_330),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_343),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_348),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_348),
.Y(n_351)
);

AOI21x1_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_347),
.B(n_322),
.Y(n_352)
);

O2A1O1Ixp33_ASAP7_75t_SL g353 ( 
.A1(n_352),
.A2(n_350),
.B(n_345),
.C(n_344),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_353),
.A2(n_334),
.B(n_349),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_354),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_355),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_13),
.C(n_345),
.Y(n_357)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_357),
.Y(n_358)
);


endmodule