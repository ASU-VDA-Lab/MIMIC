module real_jpeg_22503_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_277, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_277;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_1),
.A2(n_2),
.B1(n_18),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_54),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_1),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_2),
.A2(n_8),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_2),
.A2(n_4),
.B1(n_18),
.B2(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_2),
.A2(n_7),
.B1(n_18),
.B2(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_2),
.A2(n_27),
.B(n_50),
.C(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_3),
.A2(n_147),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_4),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_30),
.B1(n_65),
.B2(n_66),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_50),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_7),
.A2(n_50),
.B1(n_65),
.B2(n_66),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_7),
.A2(n_25),
.B(n_26),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_7),
.B(n_28),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g185 ( 
.A1(n_7),
.A2(n_10),
.B(n_66),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_SL g208 ( 
.A1(n_7),
.A2(n_40),
.B(n_41),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_19),
.B1(n_65),
.B2(n_66),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_18),
.B(n_22),
.C(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_18),
.Y(n_22)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_10),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

BUFx3_ASAP7_75t_SL g40 ( 
.A(n_11),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_270),
.B(n_273),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_68),
.B(n_269),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_31),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_15),
.B(n_31),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_15),
.B(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_23),
.B(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_28),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_21),
.B(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_24),
.A2(n_38),
.B(n_41),
.C(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_41),
.Y(n_45)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_25),
.A2(n_42),
.B(n_50),
.C(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_28),
.A2(n_48),
.B(n_53),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_29),
.B(n_83),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_32),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_32),
.B(n_267),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_46),
.CI(n_51),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_37),
.B1(n_43),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_36),
.B(n_95),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_37),
.A2(n_94),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_38),
.A2(n_44),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_38),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_38),
.B(n_50),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_40),
.A2(n_50),
.B(n_63),
.C(n_185),
.Y(n_184)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_44),
.B(n_95),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_50),
.B(n_79),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_50),
.B(n_64),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_58),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_100),
.C(n_105),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_52),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_52),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_52),
.A2(n_92),
.B1(n_127),
.B2(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_52),
.B(n_154),
.C(n_155),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_52),
.A2(n_105),
.B1(n_127),
.B2(n_165),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_56),
.A2(n_58),
.B1(n_113),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_56),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_57),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_58),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_64),
.B1(n_67),
.B2(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_64),
.B1(n_90),
.B2(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_65),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_266),
.B(n_268),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_122),
.A3(n_133),
.B1(n_264),
.B2(n_265),
.C(n_277),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_107),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_71),
.B(n_107),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_91),
.C(n_98),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_72),
.B(n_91),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_85),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_82),
.B2(n_84),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_74),
.A2(n_75),
.B1(n_86),
.B2(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_82),
.B(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_77),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_78),
.A2(n_79),
.B1(n_148),
.B2(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_79),
.A2(n_102),
.B(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_86),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_96),
.B(n_97),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_96),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_92),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_170),
.C(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_92),
.A2(n_154),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_109),
.C(n_119),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_98),
.A2(n_99),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_100),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_101),
.A2(n_103),
.B1(n_200),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_101),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_103),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_103),
.B(n_159),
.C(n_199),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_103),
.A2(n_200),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_103),
.B(n_218),
.C(n_223),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_110),
.C(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_150),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_105),
.A2(n_140),
.B1(n_141),
.B2(n_165),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_105),
.B(n_141),
.C(n_206),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_118),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_118),
.B1(n_126),
.B2(n_131),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_118),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_110),
.A2(n_118),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_110),
.B(n_239),
.C(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_117),
.C(n_118),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_118),
.B(n_131),
.C(n_132),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_123),
.B(n_124),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_258),
.B(n_263),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_246),
.B(n_257),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_175),
.B(n_231),
.C(n_245),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_161),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_137),
.B(n_161),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_152),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_139),
.B(n_149),
.C(n_152),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_141),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_140),
.B(n_145),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_141),
.B(n_184),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

NOR2x1_ASAP7_75t_R g190 ( 
.A(n_159),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_191),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_168),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.C(n_169),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_162),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_169),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_230),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_225),
.B(n_229),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_215),
.B(n_224),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_203),
.B(n_214),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_194),
.B(n_202),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_193),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B(n_192),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_205),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_212),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_227),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_232),
.B(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_243),
.B2(n_244),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_238),
.C(n_244),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_243),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_248),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_256),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_254),
.C(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);


endmodule