module fake_netlist_5_1817_n_165 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_165);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_165;

wire n_137;
wire n_164;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_136;
wire n_86;
wire n_124;
wire n_146;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_78;
wire n_65;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_30;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVxp33_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_1),
.B(n_3),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_3),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_4),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_33),
.B1(n_51),
.B2(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_5),
.C(n_6),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_51),
.B1(n_48),
.B2(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_54),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_42),
.B1(n_43),
.B2(n_49),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_43),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_34),
.B1(n_41),
.B2(n_31),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_26),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_SL g83 ( 
.A(n_59),
.B(n_57),
.C(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_22),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_21),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_58),
.C(n_61),
.Y(n_91)
);

AOI21x1_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_73),
.B(n_56),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_73),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_64),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_64),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_60),
.B(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_58),
.B1(n_61),
.B2(n_71),
.C(n_68),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_66),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_79),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_83),
.B(n_80),
.C(n_79),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_83),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_82),
.B(n_88),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_80),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_85),
.B1(n_76),
.B2(n_80),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_76),
.B1(n_82),
.B2(n_86),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_81),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_100),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_94),
.Y(n_114)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_102),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_111),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_109),
.Y(n_126)
);

NAND4xp25_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_108),
.C(n_71),
.D(n_81),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_112),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_111),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_107),
.B1(n_110),
.B2(n_96),
.C(n_67),
.Y(n_133)
);

AOI31xp33_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_110),
.A3(n_114),
.B(n_82),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_114),
.B(n_64),
.C(n_67),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_65),
.B(n_62),
.C(n_56),
.Y(n_136)
);

AOI221xp5_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_130),
.B1(n_65),
.B2(n_62),
.C(n_129),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_130),
.B(n_132),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_122),
.B1(n_120),
.B2(n_126),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_129),
.B(n_104),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_120),
.B1(n_122),
.B2(n_129),
.Y(n_141)
);

NAND5xp2_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_124),
.C(n_89),
.D(n_90),
.E(n_92),
.Y(n_142)
);

NOR4xp25_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_124),
.C(n_128),
.D(n_10),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_82),
.B1(n_129),
.B2(n_95),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_8),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_9),
.Y(n_149)
);

NAND2x1_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_140),
.Y(n_152)
);

AOI211xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_153)
);

NAND4xp75_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_94),
.C(n_84),
.D(n_95),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_87),
.C(n_98),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

OAI211xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_147),
.B(n_151),
.C(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_156),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_157),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_160),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_158),
.B1(n_159),
.B2(n_163),
.Y(n_165)
);


endmodule