module real_jpeg_23004_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_344, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_344;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx6_ASAP7_75t_L g107 ( 
.A(n_0),
.Y(n_107)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_2),
.A2(n_42),
.B1(n_44),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_2),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_128),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_128),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_2),
.A2(n_59),
.B1(n_60),
.B2(n_128),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_3),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_61),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_61),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_61),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_42),
.B1(n_44),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_51),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_116)
);

INVx8_ASAP7_75t_SL g65 ( 
.A(n_7),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_59),
.B1(n_68),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_42),
.B1(n_44),
.B2(n_71),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_71),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_71),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_9),
.A2(n_42),
.B1(n_44),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_126),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_126),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_126),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_11),
.B(n_69),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_11),
.B(n_29),
.C(n_33),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_132),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_45),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_11),
.A2(n_106),
.B1(n_151),
.B2(n_208),
.Y(n_207)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_13),
.A2(n_131),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_13),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_42),
.B1(n_44),
.B2(n_137),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_137),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_137),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_15),
.A2(n_37),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_15),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.C(n_77),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_20),
.A2(n_72),
.B1(n_328),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_20),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_38),
.B2(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_22),
.B(n_72),
.C(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_22),
.A2(n_23),
.B1(n_78),
.B2(n_79),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_23),
.B(n_38),
.C(n_54),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_32),
.B(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_24),
.A2(n_35),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_24),
.A2(n_32),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_24),
.A2(n_32),
.B1(n_184),
.B2(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_24),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_24),
.A2(n_32),
.B1(n_114),
.B2(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_24),
.A2(n_122),
.B(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_27),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_26),
.B(n_42),
.C(n_48),
.Y(n_224)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_27),
.B(n_180),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_27),
.A2(n_47),
.B(n_223),
.C(n_224),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_32),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_32),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_32),
.B(n_132),
.Y(n_214)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_33),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_34),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_36),
.B(n_123),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_49),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_40),
.A2(n_81),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_41),
.A2(n_45),
.B(n_52),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_41),
.Y(n_268)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_44),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_42),
.A2(n_64),
.B(n_133),
.C(n_154),
.Y(n_153)
);

HAxp5_ASAP7_75t_SL g223 ( 
.A(n_42),
.B(n_132),
.CON(n_223),
.SN(n_223)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_44),
.B(n_60),
.C(n_65),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_45),
.B(n_50),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_45),
.A2(n_52),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_45),
.A2(n_52),
.B1(n_164),
.B2(n_223),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_45),
.A2(n_52),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_46),
.A2(n_81),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_46),
.A2(n_49),
.B(n_298),
.Y(n_297)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_63),
.B(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_70),
.B(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_62),
.A2(n_69),
.B1(n_130),
.B2(n_134),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_62),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_62),
.A2(n_69),
.B1(n_144),
.B2(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_63),
.A2(n_135),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_69),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_72),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_72),
.Y(n_328)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_75),
.B(n_132),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_77),
.B(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_82),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_80),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_81),
.A2(n_82),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_89),
.A2(n_142),
.B(n_314),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_325),
.A3(n_336),
.B1(n_341),
.B2(n_342),
.C(n_344),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_303),
.B(n_324),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_280),
.B(n_302),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_172),
.B(n_256),
.C(n_279),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_156),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_101),
.B(n_156),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_138),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_118),
.B2(n_119),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_103),
.B(n_119),
.C(n_138),
.Y(n_257)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_113),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_105),
.B(n_113),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_108),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_112),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_106),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_106),
.A2(n_111),
.B1(n_201),
.B2(n_208),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_106),
.A2(n_107),
.B(n_287),
.Y(n_286)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_107),
.Y(n_170)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_107),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_110),
.A2(n_195),
.B(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_115),
.B(n_246),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_117),
.A2(n_123),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.C(n_129),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_125),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_158),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B(n_133),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_147),
.B2(n_155),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_141),
.B(n_145),
.C(n_155),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_142),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_153),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_161),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_157),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_160),
.B(n_161),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_162),
.B(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_171),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_255),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_250),
.B(n_254),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_235),
.B(n_249),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_219),
.B(n_234),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_196),
.B(n_218),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_185),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_181),
.B1(n_182),
.B2(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_194),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_195),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_205),
.B(n_217),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_203),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_213),
.B(n_216),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_233),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_233),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_228),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_229),
.C(n_232),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_222),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_231),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_236),
.B(n_237),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_244),
.C(n_247),
.Y(n_253)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_258),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_278),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_269),
.B1(n_276),
.B2(n_277),
.Y(n_259)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_264),
.C(n_266),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_265),
.Y(n_294)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_276),
.C(n_278),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_274),
.Y(n_299)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_282),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_301),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_290),
.C(n_301),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_286),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_285),
.A2(n_309),
.B(n_313),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_288),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_299),
.B2(n_300),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_297),
.C(n_300),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_296),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_298),
.Y(n_320)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_305),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_323),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_316),
.B2(n_317),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_316),
.C(n_323),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_315),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_311),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B(n_322),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_322),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_327),
.B1(n_331),
.B2(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_333),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_333),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.C(n_332),
.Y(n_326)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_327),
.Y(n_340)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_337),
.B(n_338),
.Y(n_341)
);


endmodule