module real_jpeg_4706_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_0),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_0),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_0),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_0),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_0),
.B(n_250),
.Y(n_249)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_2),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_2),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_2),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_2),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_2),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_36),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_4),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_5),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_5),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_6),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_7),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_7),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_7),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_7),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_7),
.B(n_54),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_7),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_7),
.B(n_66),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_7),
.B(n_287),
.Y(n_286)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_9),
.Y(n_136)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_9),
.Y(n_232)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_12),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_12),
.B(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_13),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_13),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_14),
.B(n_80),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_14),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_14),
.B(n_56),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_14),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_14),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_14),
.B(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_15),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_15),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_16),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_16),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_17),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_17),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_17),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_17),
.B(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_17),
.B(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_203),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_202),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_174),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_22),
.B(n_174),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_106),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_67),
.C(n_83),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_24),
.B(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_46),
.C(n_57),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_25),
.A2(n_26),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_27),
.B(n_34),
.C(n_45),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_28),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_32),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_40),
.B2(n_45),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_39),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_39),
.Y(n_216)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_47),
.B(n_58),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_48),
.B(n_53),
.Y(n_308)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_56),
.Y(n_147)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJx2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_65),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_59),
.B(n_61),
.CI(n_65),
.CON(n_305),
.SN(n_305)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_64),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_64),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_67),
.B(n_83),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_75),
.C(n_79),
.Y(n_123)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_73),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_96),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_85),
.B(n_91),
.C(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_95),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_96),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.C(n_103),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_97),
.B(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_99),
.Y(n_198)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_102),
.Y(n_219)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_138),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_121),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_158),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.C(n_157),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_140),
.A2(n_141),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_146),
.C(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_150),
.B(n_153),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_161),
.B1(n_172),
.B2(n_173),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_170),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_168),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_199),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_176),
.B(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_178),
.B(n_199),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_194),
.C(n_195),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_179),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.C(n_192),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_180),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_280)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_188),
.B(n_193),
.Y(n_302)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_194),
.Y(n_322)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

AOI21x1_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_326),
.B(n_330),
.Y(n_203)
);

OAI21x1_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_313),
.B(n_325),
.Y(n_204)
);

AOI21x1_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_298),
.B(n_312),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_270),
.B(n_297),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_245),
.B(n_269),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_223),
.B(n_244),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_220),
.B(n_222),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_218),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_217),
.Y(n_224)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_225),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_236),
.C(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_231),
.Y(n_257)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_240),
.B2(n_241),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_268),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_268),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_258),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_257),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_257),
.C(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_254),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_283),
.C(n_284),
.Y(n_282)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_273),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_281),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_282),
.C(n_285),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_277),
.C(n_280),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_292),
.C(n_295),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_288)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_292),
.Y(n_296)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_311),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_311),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_303),
.C(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_308),
.C(n_309),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_305),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_323),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_323),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_317),
.C(n_320),
.Y(n_329)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_329),
.Y(n_330)
);


endmodule