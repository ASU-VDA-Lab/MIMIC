module fake_jpeg_30939_n_427 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_427);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_427;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_9),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_55),
.B(n_74),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_32),
.B(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_82),
.Y(n_93)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_80),
.Y(n_104)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_18),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_81),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_33),
.B(n_18),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_87),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_24),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_8),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_24),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_37),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_34),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_92),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_56),
.B1(n_68),
.B2(n_59),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_116),
.B1(n_66),
.B2(n_73),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_50),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_117),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_42),
.B(n_25),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_76),
.C(n_52),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_22),
.B1(n_24),
.B2(n_38),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_50),
.Y(n_117)
);

HAxp5_ASAP7_75t_SL g121 ( 
.A(n_71),
.B(n_37),
.CON(n_121),
.SN(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_36),
.B(n_43),
.C(n_41),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_43),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_127),
.B(n_130),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_47),
.B(n_41),
.Y(n_130)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_93),
.B(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_135),
.B(n_144),
.Y(n_197)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_142),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_167),
.B1(n_169),
.B2(n_98),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_97),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_34),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_150),
.CI(n_151),
.CON(n_170),
.SN(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

OR2x2_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_166),
.Y(n_183)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g195 ( 
.A(n_149),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_19),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_23),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_23),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_155),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_36),
.B(n_26),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_26),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_67),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_163),
.B1(n_107),
.B2(n_96),
.Y(n_180)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_131),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_99),
.A2(n_79),
.B1(n_75),
.B2(n_77),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_126),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_151),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_172),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_103),
.B1(n_115),
.B2(n_120),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_180),
.B1(n_184),
.B2(n_143),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_96),
.B1(n_115),
.B2(n_120),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_175),
.B1(n_157),
.B2(n_180),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_103),
.B1(n_123),
.B2(n_98),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_202),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_150),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_204),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_145),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_208),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_147),
.B1(n_161),
.B2(n_158),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_153),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_139),
.C(n_140),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

OR2x4_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_148),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_154),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_122),
.B1(n_187),
.B2(n_159),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_177),
.A2(n_149),
.B1(n_169),
.B2(n_125),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_152),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_189),
.Y(n_216)
);

CKINVDCx11_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_217),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_184),
.B(n_16),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_174),
.B(n_137),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_134),
.B(n_165),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_195),
.B(n_194),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_223),
.A2(n_230),
.B(n_179),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_239),
.B1(n_244),
.B2(n_192),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_222),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_231),
.B1(n_216),
.B2(n_221),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_195),
.B(n_194),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_219),
.B1(n_214),
.B2(n_212),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_241),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_201),
.A2(n_187),
.B1(n_186),
.B2(n_190),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_194),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_186),
.B1(n_190),
.B2(n_185),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_198),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_199),
.A2(n_156),
.B1(n_193),
.B2(n_196),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_271),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_242),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

AO22x1_ASAP7_75t_SL g250 ( 
.A1(n_245),
.A2(n_206),
.B1(n_208),
.B2(n_207),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_252),
.Y(n_279)
);

AOI22x1_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_238),
.B1(n_231),
.B2(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_251),
.Y(n_300)
);

OA22x2_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_205),
.B1(n_213),
.B2(n_215),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_233),
.B(n_202),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_254),
.B(n_257),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_255),
.A2(n_265),
.B1(n_239),
.B2(n_236),
.Y(n_290)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_240),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_234),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_260),
.B(n_261),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_235),
.A2(n_204),
.B(n_182),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_269),
.B(n_271),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_182),
.B(n_195),
.C(n_146),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_264),
.A2(n_266),
.B(n_268),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_209),
.B1(n_193),
.B2(n_196),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_192),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_267),
.B(n_275),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_179),
.B(n_167),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_225),
.B(n_246),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_277),
.B1(n_141),
.B2(n_48),
.Y(n_295)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_192),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_38),
.B1(n_27),
.B2(n_39),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_292),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_240),
.C(n_247),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_302),
.C(n_251),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_252),
.B1(n_274),
.B2(n_253),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_291),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_263),
.B(n_203),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_266),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_259),
.A2(n_236),
.B(n_164),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_294),
.A2(n_118),
.B(n_124),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_295),
.A2(n_265),
.B1(n_276),
.B2(n_262),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_160),
.Y(n_298)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_273),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_90),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_131),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_124),
.C(n_118),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_269),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_304),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_325),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_307),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_250),
.C(n_266),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_320),
.C(n_282),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_309),
.A2(n_316),
.B1(n_327),
.B2(n_305),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_317),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_315),
.A2(n_313),
.B1(n_318),
.B2(n_310),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_273),
.B1(n_252),
.B2(n_256),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_252),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_294),
.B1(n_282),
.B2(n_286),
.Y(n_331)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_94),
.C(n_105),
.Y(n_320)
);

FAx1_ASAP7_75t_L g321 ( 
.A(n_279),
.B(n_300),
.CI(n_301),
.CON(n_321),
.SN(n_321)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_279),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_293),
.A2(n_11),
.B(n_16),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_322),
.A2(n_283),
.B(n_8),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_0),
.Y(n_323)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_39),
.B1(n_94),
.B2(n_27),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_325),
.Y(n_362)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_336),
.B(n_321),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_302),
.C(n_297),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_342),
.C(n_351),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_316),
.B1(n_309),
.B2(n_327),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_297),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_341),
.B(n_347),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_317),
.C(n_320),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_344),
.A2(n_350),
.B1(n_285),
.B2(n_286),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_323),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_295),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_348),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_305),
.Y(n_351)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_353),
.A2(n_337),
.B1(n_38),
.B2(n_27),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_354),
.A2(n_366),
.B1(n_331),
.B2(n_346),
.Y(n_370)
);

AO221x1_ASAP7_75t_L g355 ( 
.A1(n_334),
.A2(n_326),
.B1(n_287),
.B2(n_289),
.C(n_296),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_329),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_357),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_363),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_328),
.C(n_296),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_343),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_364),
.B(n_365),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_289),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_287),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_109),
.C(n_57),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_368),
.B(n_369),
.C(n_342),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_341),
.Y(n_369)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_370),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_367),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_359),
.A2(n_338),
.B(n_351),
.Y(n_372)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

AOI211xp5_ASAP7_75t_L g375 ( 
.A1(n_360),
.A2(n_347),
.B(n_337),
.C(n_49),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_375),
.B(n_377),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_376),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_81),
.C(n_128),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_128),
.C(n_72),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_378),
.B(n_379),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_54),
.C(n_22),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_78),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_382),
.B(n_358),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_380),
.Y(n_384)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_385),
.B(n_379),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_362),
.C(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_387),
.B(n_388),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_357),
.Y(n_390)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_357),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_395),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_361),
.C(n_101),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_396),
.B(n_400),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_374),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_402),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_390),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_381),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_381),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_404),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_361),
.Y(n_405)
);

NOR4xp25_ASAP7_75t_L g408 ( 
.A(n_405),
.B(n_382),
.C(n_13),
.D(n_14),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_392),
.B(n_378),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_391),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_410),
.Y(n_415)
);

AOI21x1_ASAP7_75t_L g416 ( 
.A1(n_408),
.A2(n_412),
.B(n_401),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_64),
.C(n_101),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_403),
.A2(n_90),
.B1(n_7),
.B2(n_11),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_6),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_400),
.B(n_7),
.Y(n_412)
);

AOI322xp5_ASAP7_75t_L g420 ( 
.A1(n_416),
.A2(n_418),
.A3(n_419),
.B1(n_413),
.B2(n_409),
.C1(n_14),
.C2(n_6),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_413),
.A2(n_399),
.B(n_396),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_417),
.A2(n_13),
.B(n_15),
.Y(n_421)
);

OAI321xp33_ASAP7_75t_L g419 ( 
.A1(n_414),
.A2(n_6),
.A3(n_17),
.B1(n_15),
.B2(n_4),
.C(n_5),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_420),
.B(n_421),
.C(n_422),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_415),
.A2(n_17),
.B(n_1),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_423),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_424),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_90),
.Y(n_426)
);

OAI321xp33_ASAP7_75t_L g427 ( 
.A1(n_426),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_217),
.C(n_400),
.Y(n_427)
);


endmodule