module fake_jpeg_19313_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx24_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g10 ( 
.A1(n_1),
.A2(n_5),
.B(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_0),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_8),
.C(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_5),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_15),
.B(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_0),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_8),
.A2(n_10),
.B1(n_11),
.B2(n_9),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_8),
.B1(n_11),
.B2(n_6),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_10),
.B(n_1),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_8),
.B1(n_13),
.B2(n_9),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_1),
.C(n_2),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_25),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_17),
.B1(n_12),
.B2(n_14),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_24),
.B1(n_19),
.B2(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_25),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_1),
.B(n_2),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_3),
.C(n_4),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_26),
.C(n_3),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.A3(n_3),
.B1(n_4),
.B2(n_30),
.C1(n_14),
.C2(n_29),
.Y(n_33)
);


endmodule