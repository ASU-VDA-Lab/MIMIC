module fake_jpeg_15942_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_14),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_29),
.B1(n_31),
.B2(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_63),
.B1(n_17),
.B2(n_40),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_22),
.C(n_26),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_62),
.C(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_22),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_31),
.B1(n_29),
.B2(n_17),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_40),
.B1(n_34),
.B2(n_23),
.Y(n_83)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_21),
.C(n_24),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_64),
.A2(n_43),
.B1(n_20),
.B2(n_23),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_21),
.B1(n_20),
.B2(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_77),
.B1(n_83),
.B2(n_52),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_25),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_73),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_42),
.B1(n_37),
.B2(n_38),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_46),
.B1(n_61),
.B2(n_52),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_21),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_27),
.B(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_86),
.B(n_104),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_58),
.B1(n_53),
.B2(n_59),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_54),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_103),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_62),
.B(n_54),
.Y(n_92)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_99),
.B(n_107),
.C(n_77),
.D(n_76),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_95),
.B1(n_83),
.B2(n_80),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_24),
.B(n_1),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_43),
.B1(n_53),
.B2(n_27),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_43),
.B1(n_44),
.B2(n_27),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_81),
.Y(n_120)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_69),
.A2(n_44),
.B(n_25),
.C(n_16),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_107),
.B(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_114),
.B(n_117),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_119),
.B1(n_90),
.B2(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_85),
.B1(n_68),
.B2(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_123),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_68),
.B1(n_75),
.B2(n_70),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_125),
.B1(n_102),
.B2(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_16),
.B(n_15),
.C(n_75),
.D(n_67),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_124),
.A2(n_107),
.B(n_88),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_67),
.B1(n_15),
.B2(n_65),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_15),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_0),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_130),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_1),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_95),
.B(n_86),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_138),
.B(n_139),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_146),
.C(n_151),
.Y(n_152)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_102),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_108),
.B1(n_100),
.B2(n_3),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_157),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_2),
.Y(n_184)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_122),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_149),
.C(n_132),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_183),
.C(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_141),
.B1(n_139),
.B2(n_131),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_172),
.A2(n_174),
.B1(n_178),
.B2(n_181),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_127),
.B(n_144),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_166),
.A2(n_138),
.B(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_177),
.B(n_182),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_140),
.B1(n_122),
.B2(n_137),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_124),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_155),
.B1(n_164),
.B2(n_159),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_125),
.B1(n_146),
.B2(n_133),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_161),
.A2(n_129),
.B(n_142),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_151),
.C(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_174),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_154),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_194),
.Y(n_199)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_158),
.B(n_180),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_154),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_168),
.C(n_162),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_196),
.C(n_172),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_162),
.C(n_160),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_180),
.B1(n_178),
.B2(n_182),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_193),
.B1(n_158),
.B2(n_108),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_200),
.C(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_181),
.C(n_160),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_206),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_205),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_213),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_201),
.A2(n_189),
.B1(n_187),
.B2(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_200),
.B(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_204),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_202),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_218),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

AOI31xp33_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_198),
.A3(n_169),
.B(n_163),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_209),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_223),
.B1(n_3),
.B2(n_4),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_215),
.B(n_211),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_226),
.A3(n_227),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_213),
.B(n_163),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_229),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_226),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_229)
);

AOI321xp33_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.C(n_13),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_9),
.Y(n_232)
);


endmodule