module fake_jpeg_16132_n_186 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_40),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_1),
.B(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_24),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_49),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_47),
.Y(n_94)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_27),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_55),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_4),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_23),
.B1(n_16),
.B2(n_26),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_60),
.B(n_17),
.Y(n_80)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_59),
.Y(n_79)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_28),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_83),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_34),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_75),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_78),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_31),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_42),
.B1(n_32),
.B2(n_16),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_85),
.B1(n_78),
.B2(n_92),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_26),
.B1(n_23),
.B2(n_74),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_29),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_44),
.B1(n_66),
.B2(n_32),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_86),
.B1(n_18),
.B2(n_22),
.Y(n_97)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_26),
.B1(n_16),
.B2(n_15),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_31),
.C(n_20),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_88),
.B(n_9),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_22),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_4),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_47),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_5),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_6),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_100),
.B1(n_86),
.B2(n_76),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_106),
.B1(n_7),
.B2(n_8),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_113),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_15),
.B1(n_20),
.B2(n_19),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_62),
.B1(n_19),
.B2(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_70),
.B(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_112),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_116),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_7),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_121),
.B1(n_127),
.B2(n_98),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_84),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_116),
.B1(n_99),
.B2(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_94),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_134),
.C(n_94),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_8),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_138),
.A2(n_139),
.B1(n_145),
.B2(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_108),
.B1(n_97),
.B2(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_98),
.B1(n_105),
.B2(n_69),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_105),
.B(n_94),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_118),
.B(n_132),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_154),
.C(n_159),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_152),
.A2(n_157),
.B1(n_136),
.B2(n_137),
.Y(n_163)
);

NOR4xp25_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_134),
.C(n_117),
.D(n_119),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_138),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_131),
.C(n_124),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_146),
.B(n_148),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_124),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_163),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_150),
.B(n_156),
.Y(n_169)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_145),
.B(n_148),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_144),
.B(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_168),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_144),
.B1(n_135),
.B2(n_143),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_142),
.C(n_143),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_169),
.A2(n_170),
.B(n_121),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_120),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_177),
.B(n_81),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_161),
.B1(n_154),
.B2(n_168),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_178),
.A3(n_173),
.B1(n_162),
.B2(n_13),
.C1(n_14),
.C2(n_11),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_162),
.C(n_160),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_144),
.B(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_179),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_175),
.B(n_183),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_182),
.Y(n_186)
);


endmodule