module real_aes_6284_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_516;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g463 ( .A1(n_0), .A2(n_143), .B(n_464), .C(n_467), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_1), .B(n_458), .Y(n_469) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g181 ( .A(n_3), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_4), .B(n_144), .Y(n_541) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_5), .A2(n_122), .B1(n_123), .B2(n_429), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_5), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_5), .A2(n_95), .B1(n_429), .B2(n_733), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_6), .A2(n_443), .B(n_490), .Y(n_489) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_7), .A2(n_150), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_8), .A2(n_36), .B1(n_147), .B2(n_199), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_9), .B(n_150), .Y(n_167) );
AND2x6_ASAP7_75t_L g152 ( .A(n_10), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_11), .A2(n_152), .B(n_446), .C(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_12), .B(n_38), .Y(n_113) );
INVx1_ASAP7_75t_L g134 ( .A(n_13), .Y(n_134) );
INVx1_ASAP7_75t_L g173 ( .A(n_14), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_15), .B(n_140), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_16), .B(n_144), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_17), .B(n_130), .Y(n_129) );
AO32x2_ASAP7_75t_L g210 ( .A1(n_18), .A2(n_150), .A3(n_151), .B1(n_170), .B2(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_19), .B(n_147), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_20), .B(n_130), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_21), .A2(n_54), .B1(n_147), .B2(n_199), .Y(n_213) );
AOI22xp33_ASAP7_75t_SL g207 ( .A1(n_22), .A2(n_79), .B1(n_140), .B2(n_147), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_23), .B(n_147), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_24), .A2(n_151), .B(n_446), .C(n_448), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_25), .A2(n_151), .B(n_446), .C(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_26), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_27), .A2(n_96), .B1(n_117), .B2(n_118), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_27), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_28), .B(n_189), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_29), .A2(n_443), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_30), .B(n_189), .Y(n_226) );
INVx2_ASAP7_75t_L g142 ( .A(n_31), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_32), .A2(n_478), .B(n_479), .C(n_483), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_33), .B(n_147), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_34), .B(n_189), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_35), .B(n_195), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_37), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_39), .B(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_40), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_41), .B(n_144), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_42), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_43), .B(n_443), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_44), .A2(n_478), .B(n_483), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_45), .B(n_147), .Y(n_160) );
INVx1_ASAP7_75t_L g465 ( .A(n_46), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_47), .A2(n_731), .B1(n_734), .B2(n_735), .Y(n_730) );
INVx1_ASAP7_75t_L g735 ( .A(n_47), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_48), .A2(n_89), .B1(n_199), .B2(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g504 ( .A(n_49), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_50), .B(n_147), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_51), .B(n_147), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_52), .B(n_443), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_53), .B(n_165), .Y(n_164) );
AOI22xp33_ASAP7_75t_SL g146 ( .A1(n_55), .A2(n_59), .B1(n_140), .B2(n_147), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_56), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_57), .B(n_147), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_58), .B(n_147), .Y(n_246) );
INVx1_ASAP7_75t_L g153 ( .A(n_60), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_61), .B(n_443), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_62), .B(n_458), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_63), .A2(n_165), .B(n_176), .C(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_64), .B(n_147), .Y(n_182) );
INVx1_ASAP7_75t_L g133 ( .A(n_65), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_66), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_67), .B(n_144), .Y(n_481) );
AO32x2_ASAP7_75t_L g203 ( .A1(n_68), .A2(n_150), .A3(n_151), .B1(n_204), .B2(n_208), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_69), .B(n_145), .Y(n_515) );
INVx1_ASAP7_75t_L g245 ( .A(n_70), .Y(n_245) );
INVx1_ASAP7_75t_L g221 ( .A(n_71), .Y(n_221) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_72), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_73), .B(n_450), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_74), .A2(n_446), .B(n_483), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_75), .B(n_140), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_76), .Y(n_491) );
INVx1_ASAP7_75t_L g107 ( .A(n_77), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_78), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_80), .B(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_81), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_82), .B(n_140), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_83), .A2(n_103), .B1(n_114), .B2(n_742), .Y(n_102) );
INVx2_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_85), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_86), .B(n_137), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_87), .B(n_140), .Y(n_161) );
OR2x2_ASAP7_75t_L g109 ( .A(n_88), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g432 ( .A(n_88), .B(n_111), .Y(n_432) );
INVx2_ASAP7_75t_L g718 ( .A(n_88), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_90), .A2(n_101), .B1(n_140), .B2(n_141), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_91), .B(n_443), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_92), .Y(n_480) );
INVxp67_ASAP7_75t_L g494 ( .A(n_93), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_94), .B(n_140), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_95), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_96), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_97), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g511 ( .A(n_98), .Y(n_511) );
INVx1_ASAP7_75t_L g540 ( .A(n_99), .Y(n_540) );
AND2x2_ASAP7_75t_L g506 ( .A(n_100), .B(n_189), .Y(n_506) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g743 ( .A(n_104), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_108), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g741 ( .A(n_109), .Y(n_741) );
NOR2x2_ASAP7_75t_L g725 ( .A(n_110), .B(n_718), .Y(n_725) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g717 ( .A(n_111), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AO221x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_726), .B1(n_729), .B2(n_736), .C(n_738), .Y(n_114) );
OAI222xp33_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_119), .B1(n_719), .B2(n_720), .C1(n_723), .C2(n_724), .Y(n_115) );
INVx1_ASAP7_75t_L g719 ( .A(n_116), .Y(n_719) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_430), .B1(n_433), .B2(n_715), .Y(n_120) );
INVx1_ASAP7_75t_L g722 ( .A(n_121), .Y(n_722) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
XNOR2xp5_ASAP7_75t_L g731 ( .A(n_123), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_363), .Y(n_123) );
NOR5xp2_ASAP7_75t_L g124 ( .A(n_125), .B(n_276), .C(n_322), .D(n_335), .E(n_347), .Y(n_124) );
OAI211xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_184), .B(n_230), .C(n_257), .Y(n_125) );
INVx1_ASAP7_75t_SL g358 ( .A(n_126), .Y(n_358) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_154), .Y(n_126) );
AND2x2_ASAP7_75t_L g282 ( .A(n_127), .B(n_155), .Y(n_282) );
AND2x2_ASAP7_75t_L g310 ( .A(n_127), .B(n_256), .Y(n_310) );
AND2x2_ASAP7_75t_L g318 ( .A(n_127), .B(n_261), .Y(n_318) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g248 ( .A(n_128), .B(n_156), .Y(n_248) );
INVx2_ASAP7_75t_L g260 ( .A(n_128), .Y(n_260) );
AND2x2_ASAP7_75t_L g385 ( .A(n_128), .B(n_327), .Y(n_385) );
OR2x2_ASAP7_75t_L g387 ( .A(n_128), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_135), .Y(n_128) );
INVx1_ASAP7_75t_L g254 ( .A(n_129), .Y(n_254) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_130), .Y(n_150) );
INVx1_ASAP7_75t_L g170 ( .A(n_130), .Y(n_170) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_131), .B(n_132), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
NAND3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_149), .C(n_151), .Y(n_135) );
AO21x1_ASAP7_75t_L g253 ( .A1(n_136), .A2(n_149), .B(n_254), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_139), .B1(n_143), .B2(n_146), .Y(n_136) );
INVx2_ASAP7_75t_L g200 ( .A(n_137), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g204 ( .A1(n_137), .A2(n_145), .B1(n_205), .B2(n_207), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_137), .A2(n_143), .B1(n_212), .B2(n_213), .Y(n_211) );
INVx4_ASAP7_75t_L g466 ( .A(n_137), .Y(n_466) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
INVx1_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
AND2x2_ASAP7_75t_L g444 ( .A(n_138), .B(n_166), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_138), .Y(n_447) );
INVx2_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx1_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_143), .A2(n_163), .B(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_143), .A2(n_180), .B(n_181), .C(n_182), .Y(n_179) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_144), .A2(n_160), .B(n_161), .Y(n_159) );
O2A1O1Ixp5_ASAP7_75t_SL g219 ( .A1(n_144), .A2(n_220), .B(n_221), .C(n_222), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_144), .A2(n_242), .B(n_243), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_144), .B(n_494), .Y(n_493) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx3_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_147), .Y(n_542) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
BUFx3_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
AND2x6_ASAP7_75t_L g446 ( .A(n_148), .B(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g458 ( .A(n_149), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_149), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_149), .A2(n_510), .B(n_517), .Y(n_509) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_149), .A2(n_537), .B(n_544), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_149), .B(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_150), .A2(n_158), .B(n_167), .Y(n_157) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_150), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_150), .A2(n_522), .B(n_523), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_151), .A2(n_241), .B(n_244), .Y(n_240) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g158 ( .A1(n_152), .A2(n_159), .B(n_162), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_152), .A2(n_172), .B(n_179), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_152), .A2(n_191), .B(n_196), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_152), .A2(n_219), .B(n_223), .Y(n_218) );
AND2x4_ASAP7_75t_L g443 ( .A(n_152), .B(n_444), .Y(n_443) );
INVx4_ASAP7_75t_SL g468 ( .A(n_152), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_152), .B(n_444), .Y(n_512) );
INVx2_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g298 ( .A(n_155), .B(n_270), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_155), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g412 ( .A(n_155), .B(n_252), .Y(n_412) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_168), .Y(n_155) );
AND2x2_ASAP7_75t_L g255 ( .A(n_156), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g302 ( .A(n_156), .Y(n_302) );
AND2x2_ASAP7_75t_L g327 ( .A(n_156), .B(n_239), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_156), .B(n_360), .Y(n_397) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g261 ( .A(n_157), .B(n_239), .Y(n_261) );
AND2x2_ASAP7_75t_L g275 ( .A(n_157), .B(n_238), .Y(n_275) );
AND2x2_ASAP7_75t_L g292 ( .A(n_157), .B(n_168), .Y(n_292) );
AND2x2_ASAP7_75t_L g349 ( .A(n_157), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_157), .B(n_256), .Y(n_362) );
AND2x2_ASAP7_75t_L g414 ( .A(n_157), .B(n_339), .Y(n_414) );
INVx2_ASAP7_75t_L g180 ( .A(n_165), .Y(n_180) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g237 ( .A(n_168), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g256 ( .A(n_168), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_168), .B(n_239), .Y(n_333) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_183), .Y(n_168) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_169), .A2(n_240), .B(n_247), .Y(n_239) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_170), .B(n_518), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_176), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_174), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_174), .A2(n_525), .B(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_176), .A2(n_540), .B(n_541), .C(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_177), .A2(n_224), .B(n_225), .Y(n_223) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g450 ( .A(n_178), .Y(n_450) );
O2A1O1Ixp5_ASAP7_75t_L g244 ( .A1(n_180), .A2(n_200), .B(n_245), .C(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_180), .A2(n_449), .B(n_451), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_214), .B(n_227), .Y(n_184) );
INVx1_ASAP7_75t_SL g346 ( .A(n_185), .Y(n_346) );
AND2x4_ASAP7_75t_L g185 ( .A(n_186), .B(n_202), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_187), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g229 ( .A(n_188), .Y(n_229) );
INVx1_ASAP7_75t_L g266 ( .A(n_188), .Y(n_266) );
AND2x2_ASAP7_75t_L g287 ( .A(n_188), .B(n_209), .Y(n_287) );
AND2x2_ASAP7_75t_L g321 ( .A(n_188), .B(n_210), .Y(n_321) );
OR2x2_ASAP7_75t_L g340 ( .A(n_188), .B(n_216), .Y(n_340) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_188), .Y(n_354) );
AND2x2_ASAP7_75t_L g367 ( .A(n_188), .B(n_368), .Y(n_367) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_201), .Y(n_188) );
INVx2_ASAP7_75t_L g208 ( .A(n_189), .Y(n_208) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_189), .A2(n_218), .B(n_226), .Y(n_217) );
INVx1_ASAP7_75t_L g456 ( .A(n_189), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_189), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_189), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_191) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_200), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_202), .A2(n_289), .B1(n_290), .B2(n_299), .Y(n_288) );
AND2x2_ASAP7_75t_L g372 ( .A(n_202), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_209), .Y(n_202) );
INVx1_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_203), .Y(n_270) );
INVx1_ASAP7_75t_L g281 ( .A(n_203), .Y(n_281) );
AND2x2_ASAP7_75t_L g296 ( .A(n_203), .B(n_210), .Y(n_296) );
INVx2_ASAP7_75t_L g467 ( .A(n_206), .Y(n_467) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_206), .Y(n_482) );
INVx1_ASAP7_75t_L g453 ( .A(n_208), .Y(n_453) );
OR2x2_ASAP7_75t_L g250 ( .A(n_209), .B(n_235), .Y(n_250) );
AND2x2_ASAP7_75t_L g280 ( .A(n_209), .B(n_281), .Y(n_280) );
NOR2xp67_ASAP7_75t_L g368 ( .A(n_209), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g228 ( .A(n_210), .B(n_229), .Y(n_228) );
BUFx2_ASAP7_75t_L g337 ( .A(n_210), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_214), .B(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g315 ( .A(n_215), .B(n_281), .Y(n_315) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g227 ( .A(n_216), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g286 ( .A(n_216), .Y(n_286) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g235 ( .A(n_217), .Y(n_235) );
OR2x2_ASAP7_75t_L g265 ( .A(n_217), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_217), .Y(n_320) );
AOI32xp33_ASAP7_75t_L g357 ( .A1(n_227), .A2(n_287), .A3(n_358), .B1(n_359), .B2(n_361), .Y(n_357) );
AND2x2_ASAP7_75t_L g283 ( .A(n_228), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_228), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_228), .B(n_315), .Y(n_401) );
INVx1_ASAP7_75t_L g406 ( .A(n_228), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_236), .B1(n_249), .B2(n_251), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
AND2x2_ASAP7_75t_L g336 ( .A(n_232), .B(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_233), .B(n_235), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_234), .A2(n_258), .B1(n_262), .B2(n_272), .Y(n_257) );
AND2x2_ASAP7_75t_L g279 ( .A(n_234), .B(n_280), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g330 ( .A1(n_234), .A2(n_248), .B(n_296), .C(n_331), .Y(n_330) );
OAI332xp33_ASAP7_75t_L g335 ( .A1(n_234), .A2(n_336), .A3(n_338), .B1(n_340), .B2(n_341), .B3(n_343), .C1(n_344), .C2(n_346), .Y(n_335) );
INVx2_ASAP7_75t_L g376 ( .A(n_234), .Y(n_376) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_235), .Y(n_294) );
INVx1_ASAP7_75t_L g369 ( .A(n_235), .Y(n_369) );
AND2x2_ASAP7_75t_L g423 ( .A(n_235), .B(n_287), .Y(n_423) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_248), .Y(n_236) );
AND2x2_ASAP7_75t_L g303 ( .A(n_238), .B(n_253), .Y(n_303) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g252 ( .A(n_239), .B(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g351 ( .A(n_239), .B(n_253), .Y(n_351) );
INVx1_ASAP7_75t_L g360 ( .A(n_239), .Y(n_360) );
INVx1_ASAP7_75t_L g334 ( .A(n_248), .Y(n_334) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g418 ( .A(n_250), .B(n_270), .Y(n_418) );
INVx1_ASAP7_75t_SL g329 ( .A(n_251), .Y(n_329) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
AND2x2_ASAP7_75t_L g356 ( .A(n_252), .B(n_314), .Y(n_356) );
INVx1_ASAP7_75t_L g375 ( .A(n_252), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_252), .B(n_342), .Y(n_377) );
INVx1_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
AND2x2_ASAP7_75t_L g278 ( .A(n_255), .B(n_259), .Y(n_278) );
AND2x2_ASAP7_75t_L g345 ( .A(n_255), .B(n_303), .Y(n_345) );
INVx2_ASAP7_75t_L g388 ( .A(n_255), .Y(n_388) );
INVx2_ASAP7_75t_L g271 ( .A(n_256), .Y(n_271) );
AND2x2_ASAP7_75t_L g273 ( .A(n_256), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
INVx1_ASAP7_75t_L g289 ( .A(n_259), .Y(n_289) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_260), .B(n_333), .Y(n_339) );
OR2x2_ASAP7_75t_L g403 ( .A(n_260), .B(n_362), .Y(n_403) );
INVx1_ASAP7_75t_L g427 ( .A(n_260), .Y(n_427) );
INVx1_ASAP7_75t_L g383 ( .A(n_261), .Y(n_383) );
AND2x2_ASAP7_75t_L g428 ( .A(n_261), .B(n_271), .Y(n_428) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_265), .A2(n_291), .B1(n_293), .B2(n_297), .Y(n_290) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI322xp33_ASAP7_75t_SL g374 ( .A1(n_268), .A2(n_375), .A3(n_376), .B1(n_377), .B2(n_378), .C1(n_381), .C2(n_383), .Y(n_374) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x2_ASAP7_75t_L g371 ( .A(n_269), .B(n_287), .Y(n_371) );
OR2x2_ASAP7_75t_L g405 ( .A(n_269), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g408 ( .A(n_269), .B(n_340), .Y(n_408) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g353 ( .A(n_270), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g409 ( .A(n_270), .B(n_340), .Y(n_409) );
INVx3_ASAP7_75t_L g342 ( .A(n_271), .Y(n_342) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_L g398 ( .A(n_273), .Y(n_398) );
AOI222xp33_ASAP7_75t_L g277 ( .A1(n_275), .A2(n_278), .B1(n_279), .B2(n_282), .C1(n_283), .C2(n_285), .Y(n_277) );
INVx1_ASAP7_75t_L g308 ( .A(n_275), .Y(n_308) );
NAND3xp33_ASAP7_75t_SL g276 ( .A(n_277), .B(n_288), .C(n_305), .Y(n_276) );
AND2x2_ASAP7_75t_L g393 ( .A(n_280), .B(n_294), .Y(n_393) );
BUFx2_ASAP7_75t_L g284 ( .A(n_281), .Y(n_284) );
INVx1_ASAP7_75t_L g325 ( .A(n_281), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_282), .A2(n_318), .B1(n_371), .B2(n_372), .C(n_374), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_284), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_287), .Y(n_311) );
AND2x2_ASAP7_75t_L g324 ( .A(n_287), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_292), .B(n_303), .Y(n_304) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
OAI21xp33_ASAP7_75t_L g299 ( .A1(n_294), .A2(n_300), .B(n_304), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_294), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g391 ( .A(n_296), .B(n_373), .Y(n_391) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g314 ( .A(n_302), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_303), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g420 ( .A(n_303), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_311), .B1(n_312), .B2(n_315), .C(n_316), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_307), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g416 ( .A(n_315), .B(n_321), .Y(n_416) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OAI31xp33_ASAP7_75t_SL g384 ( .A1(n_319), .A2(n_358), .A3(n_385), .B(n_386), .Y(n_384) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g373 ( .A(n_320), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_321), .B(n_325), .Y(n_424) );
OAI221xp5_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_326), .B1(n_328), .B2(n_329), .C(n_330), .Y(n_322) );
INVx1_ASAP7_75t_L g328 ( .A(n_324), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_327), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g343 ( .A(n_336), .Y(n_343) );
INVx2_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g365 ( .A(n_342), .B(n_351), .Y(n_365) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_342), .A2(n_359), .B(n_416), .C(n_417), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g347 ( .A1(n_343), .A2(n_348), .B1(n_352), .B2(n_355), .C(n_357), .Y(n_347) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_346), .A2(n_411), .B(n_413), .C(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_349), .A2(n_400), .B1(n_402), .B2(n_404), .C(n_407), .Y(n_399) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NOR4xp25_ASAP7_75t_L g363 ( .A(n_364), .B(n_389), .C(n_410), .D(n_421), .Y(n_363) );
OAI211xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_366), .B(n_370), .C(n_384), .Y(n_364) );
INVx1_ASAP7_75t_SL g419 ( .A(n_371), .Y(n_419) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_SL g382 ( .A(n_380), .Y(n_382) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_387), .A2(n_396), .B1(n_408), .B2(n_409), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_394), .C(n_399), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI31xp33_ASAP7_75t_L g421 ( .A1(n_392), .A2(n_422), .A3(n_424), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_432), .A2(n_434), .B1(n_717), .B2(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_SL g434 ( .A(n_435), .B(n_651), .Y(n_434) );
NOR5xp2_ASAP7_75t_L g435 ( .A(n_436), .B(n_582), .C(n_611), .D(n_631), .E(n_638), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_470), .B(n_527), .C(n_569), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_438), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_653) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_457), .Y(n_438) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_439), .Y(n_530) );
AND2x4_ASAP7_75t_L g562 ( .A(n_439), .B(n_563), .Y(n_562) );
INVx5_ASAP7_75t_L g580 ( .A(n_439), .Y(n_580) );
AND2x2_ASAP7_75t_L g589 ( .A(n_439), .B(n_581), .Y(n_589) );
AND2x2_ASAP7_75t_L g601 ( .A(n_439), .B(n_474), .Y(n_601) );
AND2x2_ASAP7_75t_L g697 ( .A(n_439), .B(n_565), .Y(n_697) );
OR2x6_ASAP7_75t_L g439 ( .A(n_440), .B(n_454), .Y(n_439) );
AOI21xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_445), .B(n_453), .Y(n_440) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx5_ASAP7_75t_L g462 ( .A(n_446), .Y(n_462) );
INVx2_ASAP7_75t_L g452 ( .A(n_450), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_452), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_452), .A2(n_482), .B(n_504), .C(n_505), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx2_ASAP7_75t_L g563 ( .A(n_457), .Y(n_563) );
AND2x2_ASAP7_75t_L g581 ( .A(n_457), .B(n_536), .Y(n_581) );
AND2x2_ASAP7_75t_L g600 ( .A(n_457), .B(n_535), .Y(n_600) );
AND2x2_ASAP7_75t_L g640 ( .A(n_457), .B(n_580), .Y(n_640) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_459), .B(n_469), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_462), .B(n_463), .C(n_468), .Y(n_460) );
INVx2_ASAP7_75t_L g478 ( .A(n_462), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_462), .A2(n_468), .B(n_491), .C(n_492), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g483 ( .A(n_468), .Y(n_483) );
INVxp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_496), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AOI322xp5_ASAP7_75t_L g699 ( .A1(n_473), .A2(n_507), .A3(n_554), .B1(n_562), .B2(n_616), .C1(n_700), .C2(n_703), .Y(n_699) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_486), .Y(n_473) );
INVx5_ASAP7_75t_L g532 ( .A(n_474), .Y(n_532) );
AND2x2_ASAP7_75t_L g548 ( .A(n_474), .B(n_534), .Y(n_548) );
BUFx2_ASAP7_75t_L g626 ( .A(n_474), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_474), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g703 ( .A(n_474), .B(n_610), .Y(n_703) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_486), .B(n_498), .Y(n_557) );
INVx1_ASAP7_75t_L g584 ( .A(n_486), .Y(n_584) );
AND2x2_ASAP7_75t_L g597 ( .A(n_486), .B(n_519), .Y(n_597) );
AND2x2_ASAP7_75t_L g698 ( .A(n_486), .B(n_616), .Y(n_698) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g552 ( .A(n_487), .B(n_498), .Y(n_552) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
OR2x2_ASAP7_75t_L g567 ( .A(n_487), .B(n_519), .Y(n_567) );
AND2x2_ASAP7_75t_L g577 ( .A(n_487), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_487), .B(n_509), .Y(n_606) );
INVxp67_ASAP7_75t_L g630 ( .A(n_487), .Y(n_630) );
AND2x2_ASAP7_75t_L g637 ( .A(n_487), .B(n_507), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_487), .B(n_519), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_487), .B(n_508), .Y(n_663) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_498), .B(n_520), .Y(n_607) );
OR2x2_ASAP7_75t_L g629 ( .A(n_498), .B(n_508), .Y(n_629) );
AND2x2_ASAP7_75t_L g642 ( .A(n_498), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_498), .B(n_597), .Y(n_648) );
OAI211xp5_ASAP7_75t_SL g652 ( .A1(n_498), .A2(n_653), .B(n_658), .C(n_667), .Y(n_652) );
AND2x2_ASAP7_75t_L g713 ( .A(n_498), .B(n_519), .Y(n_713) );
INVx5_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g566 ( .A(n_499), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_499), .B(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_499), .B(n_561), .Y(n_573) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_499), .Y(n_575) );
OR2x2_ASAP7_75t_L g586 ( .A(n_499), .B(n_508), .Y(n_586) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_499), .B(n_577), .Y(n_591) );
AND2x2_ASAP7_75t_L g616 ( .A(n_499), .B(n_508), .Y(n_616) );
AND2x2_ASAP7_75t_L g636 ( .A(n_499), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g674 ( .A(n_499), .B(n_507), .Y(n_674) );
OR2x2_ASAP7_75t_L g677 ( .A(n_499), .B(n_663), .Y(n_677) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_519), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_508), .A2(n_621), .B(n_624), .C(n_630), .Y(n_620) );
INVx5_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_509), .B(n_519), .Y(n_551) );
AND2x2_ASAP7_75t_L g555 ( .A(n_509), .B(n_520), .Y(n_555) );
OR2x2_ASAP7_75t_L g561 ( .A(n_509), .B(n_519), .Y(n_561) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_513), .Y(n_510) );
INVx1_ASAP7_75t_SL g578 ( .A(n_519), .Y(n_578) );
OR2x2_ASAP7_75t_L g706 ( .A(n_519), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_546), .B(n_549), .C(n_558), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AOI31xp33_ASAP7_75t_L g631 ( .A1(n_529), .A2(n_632), .A3(n_634), .B(n_635), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_530), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_531), .B(n_562), .Y(n_568) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_532), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g588 ( .A(n_532), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g593 ( .A(n_532), .B(n_563), .Y(n_593) );
AND2x2_ASAP7_75t_L g603 ( .A(n_532), .B(n_562), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_532), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g623 ( .A(n_532), .B(n_580), .Y(n_623) );
AND2x2_ASAP7_75t_L g628 ( .A(n_532), .B(n_600), .Y(n_628) );
OR2x2_ASAP7_75t_L g647 ( .A(n_532), .B(n_534), .Y(n_647) );
OR2x2_ASAP7_75t_L g649 ( .A(n_532), .B(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_532), .Y(n_696) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g596 ( .A(n_534), .B(n_563), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_534), .B(n_580), .Y(n_619) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g565 ( .A(n_536), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_543), .Y(n_537) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g656 ( .A(n_548), .B(n_580), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g658 ( .A1(n_548), .A2(n_562), .A3(n_600), .B1(n_659), .B2(n_660), .C1(n_661), .C2(n_664), .Y(n_658) );
INVx1_ASAP7_75t_L g666 ( .A(n_548), .Y(n_666) );
NAND2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_SL g660 ( .A(n_550), .Y(n_660) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OR2x2_ASAP7_75t_L g612 ( .A(n_551), .B(n_557), .Y(n_612) );
INVx1_ASAP7_75t_L g643 ( .A(n_551), .Y(n_643) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .A3(n_564), .B1(n_566), .B2(n_568), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AOI21xp33_ASAP7_75t_SL g598 ( .A1(n_561), .A2(n_576), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_SL g613 ( .A(n_562), .Y(n_613) );
AND2x4_ASAP7_75t_L g610 ( .A(n_563), .B(n_580), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_563), .B(n_646), .Y(n_645) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_564), .A2(n_591), .A3(n_610), .B1(n_643), .B2(n_676), .C1(n_678), .C2(n_679), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_564), .A2(n_641), .B1(n_705), .B2(n_706), .C(n_708), .Y(n_704) );
AND2x2_ASAP7_75t_L g592 ( .A(n_565), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g572 ( .A(n_567), .Y(n_572) );
OR2x2_ASAP7_75t_L g644 ( .A(n_567), .B(n_629), .Y(n_644) );
OAI31xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_573), .A3(n_574), .B(n_579), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_570), .A2(n_603), .B1(n_604), .B2(n_608), .Y(n_602) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g615 ( .A(n_572), .B(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_574), .A2(n_615), .B1(n_668), .B2(n_671), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g657 ( .A(n_577), .B(n_626), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_577), .B(n_616), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_578), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g691 ( .A(n_578), .B(n_629), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_579), .A2(n_674), .B1(n_687), .B2(n_690), .Y(n_686) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx2_ASAP7_75t_L g595 ( .A(n_580), .Y(n_595) );
AND2x2_ASAP7_75t_L g678 ( .A(n_580), .B(n_600), .Y(n_678) );
OR2x2_ASAP7_75t_L g680 ( .A(n_580), .B(n_647), .Y(n_680) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_580), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_581), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_581), .B(n_626), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_587), .B(n_590), .C(n_602), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_594), .B2(n_597), .C(n_598), .Y(n_590) );
INVxp67_ASAP7_75t_L g702 ( .A(n_593), .Y(n_702) );
INVx1_ASAP7_75t_L g669 ( .A(n_594), .Y(n_669) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g633 ( .A(n_595), .B(n_600), .Y(n_633) );
INVx1_ASAP7_75t_L g650 ( .A(n_596), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_596), .B(n_623), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g665 ( .A(n_600), .Y(n_665) );
AND2x2_ASAP7_75t_L g671 ( .A(n_600), .B(n_626), .Y(n_671) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_SL g659 ( .A(n_607), .Y(n_659) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_610), .B(n_646), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B1(n_614), .B2(n_617), .C(n_620), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g707 ( .A(n_616), .Y(n_707) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g625 ( .A(n_619), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_623), .B(n_682), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_629), .Y(n_624) );
OAI211xp5_ASAP7_75t_SL g672 ( .A1(n_627), .A2(n_673), .B(n_675), .C(n_681), .Y(n_672) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g684 ( .A(n_629), .Y(n_684) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI222xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B1(n_644), .B2(n_645), .C1(n_648), .C2(n_649), .Y(n_638) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g714 ( .A(n_645), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_646), .B(n_689), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_646), .A2(n_693), .B1(n_695), .B2(n_698), .Y(n_692) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
NOR4xp25_ASAP7_75t_L g651 ( .A(n_652), .B(n_672), .C(n_685), .D(n_704), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_654), .B(n_684), .Y(n_694) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g661 ( .A(n_659), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_662), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_692), .C(n_699), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx2_ASAP7_75t_L g701 ( .A(n_697), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_711), .B(n_714), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g737 ( .A(n_727), .Y(n_737) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g734 ( .A(n_731), .Y(n_734) );
BUFx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
endmodule