module fake_jpeg_22401_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_0),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_20),
.B1(n_25),
.B2(n_37),
.Y(n_76)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_62),
.Y(n_98)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_37),
.B1(n_20),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_72),
.B1(n_85),
.B2(n_90),
.Y(n_101)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_70),
.B(n_77),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_30),
.B1(n_23),
.B2(n_24),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_33),
.B1(n_31),
.B2(n_93),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_37),
.B1(n_20),
.B2(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_53),
.B(n_19),
.Y(n_115)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_25),
.B1(n_24),
.B2(n_28),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_89),
.B1(n_35),
.B2(n_32),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_32),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_9),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_25),
.B1(n_34),
.B2(n_35),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_22),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_19),
.Y(n_109)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_90),
.B1(n_55),
.B2(n_57),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_43),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_94),
.B(n_107),
.C(n_111),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_103),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_97),
.A2(n_116),
.B1(n_117),
.B2(n_127),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_31),
.B(n_38),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_114),
.Y(n_136)
);

NAND2xp67_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_26),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_46),
.C(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_13),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_53),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_53),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_115),
.A2(n_126),
.B1(n_27),
.B2(n_21),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_46),
.B1(n_51),
.B2(n_42),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_51),
.B1(n_42),
.B2(n_17),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_38),
.C(n_33),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_75),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_129),
.B1(n_59),
.B2(n_39),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_0),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_80),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_60),
.A2(n_17),
.B1(n_27),
.B2(n_21),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_75),
.A2(n_39),
.B1(n_27),
.B2(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_130),
.B(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_95),
.B(n_13),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_95),
.B(n_13),
.Y(n_134)
);

AO22x1_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_69),
.B1(n_67),
.B2(n_83),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_135),
.A2(n_96),
.B1(n_110),
.B2(n_106),
.Y(n_180)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_137),
.B(n_142),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_139),
.A2(n_140),
.B1(n_151),
.B2(n_163),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_59),
.B1(n_67),
.B2(n_69),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_9),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_11),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_147),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_94),
.B(n_39),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_113),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_152),
.B1(n_121),
.B2(n_108),
.Y(n_179)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_157),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_151)
);

AO21x2_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_112),
.B(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_6),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_119),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_109),
.B(n_6),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_156),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_97),
.A2(n_6),
.B1(n_14),
.B2(n_12),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_162),
.B1(n_118),
.B2(n_108),
.Y(n_172)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_159),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_161),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_111),
.A2(n_123),
.B1(n_124),
.B2(n_121),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_94),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_94),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_163),
.B1(n_151),
.B2(n_134),
.Y(n_184)
);

NAND2x1_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_124),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_171),
.B(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_173),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_152),
.A2(n_113),
.B(n_114),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_125),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_177),
.B(n_182),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_190),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_125),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_110),
.B1(n_106),
.B2(n_99),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_197),
.B1(n_136),
.B2(n_14),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_152),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_114),
.B(n_3),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_141),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_189),
.B(n_193),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_160),
.B1(n_161),
.B2(n_152),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_138),
.A2(n_99),
.B1(n_96),
.B2(n_11),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

NAND2x1_ASAP7_75t_SL g192 ( 
.A(n_132),
.B(n_4),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_141),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_140),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_4),
.B1(n_5),
.B2(n_11),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_153),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_198),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_165),
.A2(n_144),
.B(n_138),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_207),
.B(n_171),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_204),
.B(n_228),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_187),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_132),
.B1(n_156),
.B2(n_137),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_220),
.B1(n_226),
.B2(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_175),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_215),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_132),
.B1(n_136),
.B2(n_150),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_221),
.B1(n_174),
.B2(n_179),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_158),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_217),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_165),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_225),
.C(n_199),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_167),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_185),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_227),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_227),
.B(n_177),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_242),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_166),
.B1(n_200),
.B2(n_224),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_219),
.B1(n_210),
.B2(n_208),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_222),
.C(n_208),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_197),
.CI(n_188),
.CON(n_241),
.SN(n_241)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_241),
.B(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_170),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_215),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_170),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_252),
.A2(n_261),
.B1(n_270),
.B2(n_258),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_262),
.C(n_267),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_238),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_236),
.A2(n_219),
.B1(n_166),
.B2(n_203),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_225),
.C(n_205),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_200),
.B1(n_168),
.B2(n_180),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_250),
.B1(n_234),
.B2(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_207),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_242),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_269),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_198),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_259),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_283),
.Y(n_300)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_281),
.B(n_282),
.Y(n_291)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_254),
.A2(n_234),
.B(n_250),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_248),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_241),
.B1(n_230),
.B2(n_251),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_SL g296 ( 
.A1(n_284),
.A2(n_267),
.B(n_241),
.C(n_261),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_280),
.B1(n_287),
.B2(n_265),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_252),
.A2(n_244),
.B(n_212),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_287),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_256),
.C(n_255),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_294),
.C(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_284),
.A2(n_224),
.B1(n_264),
.B2(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_258),
.C(n_257),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_297),
.B1(n_286),
.B2(n_231),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_257),
.C(n_260),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_249),
.B(n_265),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_299),
.A2(n_277),
.B(n_271),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_302),
.B(n_304),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_273),
.B(n_232),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_253),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_306),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_232),
.B(n_285),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_283),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_275),
.C(n_245),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_312),
.Y(n_320)
);

OAI21x1_ASAP7_75t_SL g311 ( 
.A1(n_307),
.A2(n_296),
.B(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_286),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_247),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_209),
.B(n_229),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_288),
.B1(n_298),
.B2(n_296),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_317),
.B1(n_296),
.B2(n_272),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_317),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_241),
.B(n_300),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_316),
.C(n_314),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_310),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_325),
.B(n_318),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_320),
.B(n_322),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_209),
.B(n_176),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_178),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_178),
.B1(n_169),
.B2(n_191),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_169),
.B1(n_207),
.B2(n_192),
.Y(n_332)
);


endmodule