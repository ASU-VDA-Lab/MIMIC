module real_aes_2337_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_755;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_0), .B(n_139), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_1), .A2(n_148), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_2), .B(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_3), .B(n_155), .Y(n_218) );
INVx1_ASAP7_75t_L g146 ( .A(n_4), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_5), .B(n_155), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_6), .B(n_159), .Y(n_478) );
INVx1_ASAP7_75t_L g512 ( .A(n_7), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g809 ( .A(n_8), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_9), .Y(n_550) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_10), .B(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g136 ( .A(n_11), .Y(n_136) );
AOI221x1_ASAP7_75t_L g234 ( .A1(n_12), .A2(n_24), .B1(n_139), .B2(n_148), .C(n_235), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_13), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g807 ( .A(n_13), .B(n_808), .C(n_810), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_14), .B(n_139), .Y(n_138) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_15), .A2(n_134), .B(n_137), .Y(n_133) );
INVx1_ASAP7_75t_L g487 ( .A(n_16), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_17), .B(n_173), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_18), .B(n_155), .Y(n_182) );
AO21x1_ASAP7_75t_L g213 ( .A1(n_19), .A2(n_139), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g117 ( .A(n_20), .Y(n_117) );
INVx1_ASAP7_75t_L g485 ( .A(n_21), .Y(n_485) );
INVx1_ASAP7_75t_SL g495 ( .A(n_22), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_23), .B(n_140), .Y(n_578) );
NAND2x1_ASAP7_75t_L g204 ( .A(n_25), .B(n_155), .Y(n_204) );
AOI33xp33_ASAP7_75t_L g524 ( .A1(n_26), .A2(n_52), .A3(n_462), .B1(n_467), .B2(n_525), .B3(n_526), .Y(n_524) );
NAND2x1_ASAP7_75t_L g192 ( .A(n_27), .B(n_157), .Y(n_192) );
INVx1_ASAP7_75t_L g544 ( .A(n_28), .Y(n_544) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_29), .A2(n_85), .B(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g160 ( .A(n_29), .B(n_85), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_30), .B(n_470), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_31), .B(n_157), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_32), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_33), .B(n_157), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_34), .A2(n_148), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g145 ( .A(n_35), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g149 ( .A(n_35), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g461 ( .A(n_35), .Y(n_461) );
OR2x6_ASAP7_75t_L g115 ( .A(n_36), .B(n_116), .Y(n_115) );
INVxp67_ASAP7_75t_L g810 ( .A(n_36), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_37), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_38), .B(n_139), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_39), .B(n_470), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_40), .A2(n_159), .B1(n_166), .B2(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_41), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_42), .B(n_140), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_43), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_44), .B(n_157), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_45), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_46), .B(n_134), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_47), .B(n_140), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_48), .A2(n_148), .B(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_49), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_50), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_51), .B(n_157), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_53), .B(n_140), .Y(n_536) );
INVx1_ASAP7_75t_L g142 ( .A(n_54), .Y(n_142) );
INVx1_ASAP7_75t_L g152 ( .A(n_54), .Y(n_152) );
AND2x2_ASAP7_75t_L g537 ( .A(n_55), .B(n_173), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_56), .A2(n_73), .B1(n_459), .B2(n_470), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_57), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_58), .B(n_155), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_59), .B(n_166), .Y(n_552) );
AOI21xp5_ASAP7_75t_SL g458 ( .A1(n_60), .A2(n_459), .B(n_464), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_61), .A2(n_148), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g481 ( .A(n_62), .Y(n_481) );
AO21x1_ASAP7_75t_L g215 ( .A1(n_63), .A2(n_148), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_64), .B(n_139), .Y(n_168) );
INVx1_ASAP7_75t_L g535 ( .A(n_65), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_66), .B(n_139), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_67), .A2(n_459), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g228 ( .A(n_68), .B(n_174), .Y(n_228) );
INVx1_ASAP7_75t_L g144 ( .A(n_69), .Y(n_144) );
INVx1_ASAP7_75t_L g150 ( .A(n_69), .Y(n_150) );
AND2x2_ASAP7_75t_L g196 ( .A(n_70), .B(n_165), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_71), .B(n_470), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_72), .A2(n_121), .B1(n_784), .B2(n_788), .Y(n_783) );
AND2x2_ASAP7_75t_L g497 ( .A(n_74), .B(n_165), .Y(n_497) );
INVx1_ASAP7_75t_L g482 ( .A(n_75), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_76), .A2(n_459), .B(n_494), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g576 ( .A1(n_77), .A2(n_459), .B(n_519), .C(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g118 ( .A(n_78), .Y(n_118) );
AND2x2_ASAP7_75t_L g164 ( .A(n_79), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_80), .B(n_139), .Y(n_184) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_81), .B(n_165), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_82), .A2(n_459), .B1(n_522), .B2(n_523), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g795 ( .A1(n_83), .A2(n_796), .B1(n_797), .B2(n_798), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_83), .Y(n_797) );
AND2x2_ASAP7_75t_L g214 ( .A(n_84), .B(n_159), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_86), .B(n_157), .Y(n_183) );
AND2x2_ASAP7_75t_L g208 ( .A(n_87), .B(n_165), .Y(n_208) );
INVx1_ASAP7_75t_L g465 ( .A(n_88), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_89), .B(n_155), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_90), .A2(n_148), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_91), .B(n_157), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_92), .Y(n_121) );
AND2x2_ASAP7_75t_L g528 ( .A(n_93), .B(n_165), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_94), .B(n_155), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_95), .A2(n_542), .B(n_543), .C(n_545), .Y(n_541) );
BUFx2_ASAP7_75t_L g105 ( .A(n_96), .Y(n_105) );
BUFx2_ASAP7_75t_SL g793 ( .A(n_96), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_97), .A2(n_148), .B(n_153), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_98), .B(n_140), .Y(n_468) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_803), .B(n_811), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_120), .B(n_790), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_106), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVxp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_107), .A2(n_795), .B(n_800), .Y(n_794) );
NOR2xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_119), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_R g802 ( .A(n_112), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x6_ASAP7_75t_SL g125 ( .A(n_113), .B(n_115), .Y(n_125) );
OR2x6_ASAP7_75t_SL g782 ( .A(n_113), .B(n_114), .Y(n_782) );
OR2x2_ASAP7_75t_L g789 ( .A(n_113), .B(n_115), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g806 ( .A(n_116), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B(n_783), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_126), .B1(n_449), .B2(n_782), .Y(n_123) );
INVx3_ASAP7_75t_SL g786 ( .A(n_124), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g784 ( .A1(n_127), .A2(n_782), .B1(n_785), .B2(n_787), .Y(n_784) );
INVx1_ASAP7_75t_L g796 ( .A(n_127), .Y(n_796) );
INVx2_ASAP7_75t_L g799 ( .A(n_127), .Y(n_799) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_370), .Y(n_127) );
NOR3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_282), .C(n_322), .Y(n_128) );
OAI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_197), .B1(n_246), .B2(n_261), .C(n_264), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_161), .Y(n_131) );
INVx2_ASAP7_75t_L g279 ( .A(n_132), .Y(n_279) );
AND2x2_ASAP7_75t_L g309 ( .A(n_132), .B(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g247 ( .A(n_133), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g254 ( .A(n_133), .B(n_187), .Y(n_254) );
INVx2_ASAP7_75t_L g260 ( .A(n_133), .Y(n_260) );
AND2x2_ASAP7_75t_L g269 ( .A(n_133), .B(n_163), .Y(n_269) );
INVx1_ASAP7_75t_L g285 ( .A(n_133), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_133), .B(n_331), .Y(n_330) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_134), .A2(n_510), .B(n_514), .Y(n_509) );
INVx2_ASAP7_75t_SL g519 ( .A(n_134), .Y(n_519) );
BUFx4f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
AND2x4_ASAP7_75t_L g159 ( .A(n_136), .B(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_136), .B(n_160), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_147), .B(n_159), .Y(n_137) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
INVx1_ASAP7_75t_L g483 ( .A(n_140), .Y(n_483) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
AND2x6_ASAP7_75t_L g157 ( .A(n_141), .B(n_150), .Y(n_157) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g155 ( .A(n_143), .B(n_152), .Y(n_155) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx5_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_145), .Y(n_545) );
AND2x2_ASAP7_75t_L g151 ( .A(n_146), .B(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_146), .Y(n_472) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
BUFx3_ASAP7_75t_L g473 ( .A(n_149), .Y(n_473) );
INVx2_ASAP7_75t_L g463 ( .A(n_150), .Y(n_463) );
AND2x4_ASAP7_75t_L g459 ( .A(n_151), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g467 ( .A(n_152), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_158), .Y(n_153) );
INVxp67_ASAP7_75t_L g488 ( .A(n_155), .Y(n_488) );
INVxp67_ASAP7_75t_L g486 ( .A(n_157), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_158), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_158), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_158), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_158), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_158), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_158), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_158), .A2(n_236), .B(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_158), .A2(n_465), .B(n_466), .C(n_468), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_158), .B(n_159), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g494 ( .A1(n_158), .A2(n_466), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_158), .A2(n_466), .B(n_512), .C(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g522 ( .A(n_158), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_158), .A2(n_466), .B(n_535), .C(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_158), .A2(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_SL g178 ( .A(n_159), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_159), .B(n_220), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_159), .A2(n_458), .B(n_469), .Y(n_457) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_162), .B(n_175), .Y(n_161) );
INVx4_ASAP7_75t_L g250 ( .A(n_162), .Y(n_250) );
AND2x2_ASAP7_75t_L g281 ( .A(n_162), .B(n_188), .Y(n_281) );
AND2x2_ASAP7_75t_L g357 ( .A(n_162), .B(n_331), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g399 ( .A(n_162), .B(n_187), .Y(n_399) );
INVx5_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_163), .B(n_187), .Y(n_286) );
AND2x2_ASAP7_75t_L g310 ( .A(n_163), .B(n_188), .Y(n_310) );
BUFx2_ASAP7_75t_L g326 ( .A(n_163), .Y(n_326) );
NOR2x1_ASAP7_75t_SL g429 ( .A(n_163), .B(n_331), .Y(n_429) );
OR2x6_ASAP7_75t_L g163 ( .A(n_164), .B(n_167), .Y(n_163) );
INVx3_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_165), .A2(n_207), .B1(n_541), .B2(n_546), .Y(n_540) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_166), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_173), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_173), .Y(n_195) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_173), .A2(n_234), .B(n_238), .Y(n_233) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_173), .A2(n_234), .B(n_238), .Y(n_296) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g306 ( .A(n_175), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_175), .A2(n_373), .B1(n_375), .B2(n_377), .C(n_382), .Y(n_372) );
AND2x2_ASAP7_75t_L g392 ( .A(n_175), .B(n_285), .Y(n_392) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_187), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g248 ( .A(n_177), .Y(n_248) );
INVx1_ASAP7_75t_L g301 ( .A(n_177), .Y(n_301) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_185), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_178), .B(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_178), .A2(n_179), .B(n_185), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_184), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_187), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g270 ( .A(n_187), .B(n_258), .Y(n_270) );
INVx2_ASAP7_75t_L g312 ( .A(n_187), .Y(n_312) );
AND2x2_ASAP7_75t_L g445 ( .A(n_187), .B(n_260), .Y(n_445) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_188), .Y(n_302) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_195), .A2(n_491), .B(n_497), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_229), .C(n_244), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_209), .Y(n_198) );
INVx2_ASAP7_75t_L g359 ( .A(n_199), .Y(n_359) );
AND2x2_ASAP7_75t_L g404 ( .A(n_199), .B(n_281), .Y(n_404) );
BUFx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g349 ( .A(n_200), .Y(n_349) );
AND2x4_ASAP7_75t_SL g364 ( .A(n_200), .B(n_276), .Y(n_364) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_207), .B(n_208), .Y(n_200) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_201), .A2(n_207), .B(n_208), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_206), .Y(n_201) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_207), .A2(n_222), .B(n_228), .Y(n_221) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_207), .A2(n_222), .B(n_228), .Y(n_241) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_207), .A2(n_531), .B(n_537), .Y(n_530) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_207), .A2(n_531), .B(n_537), .Y(n_560) );
INVx2_ASAP7_75t_L g318 ( .A(n_209), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_209), .B(n_348), .Y(n_374) );
AND2x4_ASAP7_75t_L g407 ( .A(n_209), .B(n_354), .Y(n_407) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
AND2x2_ASAP7_75t_L g245 ( .A(n_210), .B(n_240), .Y(n_245) );
OR2x2_ASAP7_75t_L g275 ( .A(n_210), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_210), .B(n_296), .Y(n_344) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
BUFx2_ASAP7_75t_L g289 ( .A(n_211), .Y(n_289) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
OAI21x1_ASAP7_75t_SL g212 ( .A1(n_213), .A2(n_215), .B(n_219), .Y(n_212) );
INVx1_ASAP7_75t_L g220 ( .A(n_214), .Y(n_220) );
INVx2_ASAP7_75t_L g276 ( .A(n_221), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_227), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_229), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_239), .Y(n_230) );
AND2x2_ASAP7_75t_L g244 ( .A(n_231), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g317 ( .A(n_231), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g402 ( .A(n_231), .Y(n_402) );
BUFx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_L g262 ( .A(n_232), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g381 ( .A(n_232), .B(n_241), .Y(n_381) );
AND2x2_ASAP7_75t_L g385 ( .A(n_232), .B(n_251), .Y(n_385) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g354 ( .A(n_233), .Y(n_354) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_233), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_239), .B(n_262), .Y(n_338) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_240), .B(n_263), .Y(n_448) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g252 ( .A(n_241), .B(n_243), .Y(n_252) );
AND2x2_ASAP7_75t_L g334 ( .A(n_241), .B(n_296), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_241), .B(n_242), .Y(n_353) );
BUFx2_ASAP7_75t_L g274 ( .A(n_242), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_242), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx3_ASAP7_75t_L g251 ( .A(n_243), .Y(n_251) );
INVxp67_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
INVx1_ASAP7_75t_L g267 ( .A(n_245), .Y(n_267) );
AND2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_274), .Y(n_303) );
NAND2xp33_ASAP7_75t_L g384 ( .A(n_245), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g421 ( .A(n_245), .B(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B1(n_252), .B2(n_253), .C(n_255), .Y(n_246) );
AND2x2_ASAP7_75t_L g350 ( .A(n_247), .B(n_250), .Y(n_350) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_247), .B(n_310), .Y(n_369) );
AND2x2_ASAP7_75t_L g387 ( .A(n_247), .B(n_312), .Y(n_387) );
AND2x2_ASAP7_75t_L g442 ( .A(n_247), .B(n_281), .Y(n_442) );
INVx1_ASAP7_75t_L g258 ( .A(n_248), .Y(n_258) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_248), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_249), .Y(n_394) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_250), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_250), .B(n_301), .Y(n_376) );
AND2x2_ASAP7_75t_L g343 ( .A(n_251), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g379 ( .A(n_251), .Y(n_379) );
AND2x2_ASAP7_75t_L g288 ( .A(n_252), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_252), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g430 ( .A(n_252), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_252), .B(n_354), .Y(n_440) );
AND2x4_ASAP7_75t_L g356 ( .A(n_253), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g427 ( .A(n_254), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
OR2x2_ASAP7_75t_L g298 ( .A(n_259), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g305 ( .A(n_260), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g336 ( .A(n_260), .B(n_310), .Y(n_336) );
AND2x2_ASAP7_75t_L g410 ( .A(n_260), .B(n_331), .Y(n_410) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g358 ( .A(n_262), .B(n_359), .Y(n_358) );
OAI32xp33_ASAP7_75t_L g423 ( .A1(n_262), .A2(n_424), .A3(n_426), .B1(n_427), .B2(n_430), .Y(n_423) );
AND2x4_ASAP7_75t_L g295 ( .A(n_263), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g393 ( .A(n_263), .B(n_296), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .B1(n_271), .B2(n_277), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_SL g382 ( .A1(n_266), .A2(n_280), .B(n_383), .C(n_384), .Y(n_382) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g366 ( .A(n_267), .B(n_294), .Y(n_366) );
INVx1_ASAP7_75t_SL g437 ( .A(n_268), .Y(n_437) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x4_ASAP7_75t_L g340 ( .A(n_270), .B(n_279), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_270), .A2(n_419), .B1(n_420), .B2(n_421), .C(n_423), .Y(n_418) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_275), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_278), .A2(n_308), .B1(n_361), .B2(n_362), .Y(n_360) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_279), .A2(n_397), .B(n_405), .C(n_418), .Y(n_396) );
INVx2_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g316 ( .A(n_281), .B(n_285), .Y(n_316) );
OAI211xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_287), .B(n_290), .C(n_319), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g313 ( .A(n_285), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g433 ( .A(n_285), .B(n_429), .Y(n_433) );
OAI32xp33_ASAP7_75t_L g390 ( .A1(n_286), .A2(n_391), .A3(n_393), .B1(n_394), .B2(n_395), .Y(n_390) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_289), .B(n_381), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B1(n_303), .B2(n_304), .C(n_307), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g447 ( .A(n_294), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_295), .B(n_359), .Y(n_361) );
A2O1A1O1Ixp25_ASAP7_75t_L g432 ( .A1(n_295), .A2(n_364), .B(n_380), .C(n_426), .D(n_433), .Y(n_432) );
AOI31xp33_ASAP7_75t_L g434 ( .A1(n_295), .A2(n_316), .A3(n_426), .B(n_433), .Y(n_434) );
AND2x2_ASAP7_75t_L g348 ( .A(n_296), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_298), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx2_ASAP7_75t_L g425 ( .A(n_300), .Y(n_425) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g420 ( .A(n_301), .B(n_312), .Y(n_420) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
AND2x2_ASAP7_75t_L g320 ( .A(n_304), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AOI31xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .A3(n_315), .B(n_317), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_310), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g443 ( .A(n_310), .B(n_389), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g388 ( .A(n_312), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g414 ( .A(n_312), .Y(n_414) );
INVxp67_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g321 ( .A(n_317), .Y(n_321) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND3xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_339), .C(n_355), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_332), .B1(n_336), .B2(n_337), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx2_ASAP7_75t_L g409 ( .A(n_326), .Y(n_409) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_330), .Y(n_389) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_330), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_330), .B(n_399), .Y(n_416) );
NAND2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g367 ( .A(n_334), .Y(n_367) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_350), .B2(n_351), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_342), .B(n_345), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_348), .A2(n_353), .B1(n_387), .B2(n_388), .C(n_390), .Y(n_386) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2x1_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g426 ( .A(n_353), .Y(n_426) );
AND2x2_ASAP7_75t_L g363 ( .A(n_354), .B(n_364), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_SL g411 ( .A1(n_354), .A2(n_412), .B(n_416), .C(n_417), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B(n_360), .C(n_365), .Y(n_355) );
AND2x2_ASAP7_75t_L g406 ( .A(n_359), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g417 ( .A(n_364), .Y(n_417) );
AOI21xp33_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_368), .Y(n_365) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NOR3xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_396), .C(n_431), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_372), .B(n_386), .Y(n_371) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g395 ( .A(n_380), .Y(n_395) );
INVxp67_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g403 ( .A(n_393), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B1(n_403), .B2(n_404), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B(n_411), .Y(n_405) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g444 ( .A(n_429), .B(n_445), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_435), .B2(n_438), .C(n_441), .Y(n_431) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI31xp33_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_443), .A3(n_444), .B(n_446), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g787 ( .A(n_449), .Y(n_787) );
NAND3x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_669), .C(n_746), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_621), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_452), .B(n_561), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_498), .B1(n_505), .B2(n_554), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_474), .Y(n_453) );
NOR2xp67_ASAP7_75t_SL g604 ( .A(n_454), .B(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g619 ( .A(n_454), .B(n_620), .Y(n_619) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_454), .B(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_SL g676 ( .A(n_454), .B(n_677), .Y(n_676) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_455), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_455), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g611 ( .A(n_455), .Y(n_611) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_455), .Y(n_616) );
AND2x2_ASAP7_75t_L g645 ( .A(n_455), .B(n_585), .Y(n_645) );
OR2x2_ASAP7_75t_L g649 ( .A(n_455), .B(n_490), .Y(n_649) );
AND2x4_ASAP7_75t_L g662 ( .A(n_455), .B(n_620), .Y(n_662) );
NOR2x1_ASAP7_75t_SL g664 ( .A(n_455), .B(n_477), .Y(n_664) );
AND2x2_ASAP7_75t_L g692 ( .A(n_455), .B(n_570), .Y(n_692) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
INVxp67_ASAP7_75t_L g551 ( .A(n_459), .Y(n_551) );
NOR2x1p5_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g526 ( .A(n_462), .Y(n_526) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x6_ASAP7_75t_L g466 ( .A(n_463), .B(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_466), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_480) );
INVxp67_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
INVx2_ASAP7_75t_L g580 ( .A(n_466), .Y(n_580) );
AND2x2_ASAP7_75t_L g471 ( .A(n_467), .B(n_472), .Y(n_471) );
INVxp33_ASAP7_75t_L g525 ( .A(n_467), .Y(n_525) );
INVx1_ASAP7_75t_L g553 ( .A(n_470), .Y(n_553) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g573 ( .A(n_471), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_473), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_474), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_475), .A2(n_750), .B1(n_752), .B2(n_755), .Y(n_749) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_490), .Y(n_475) );
INVx1_ASAP7_75t_L g504 ( .A(n_476), .Y(n_504) );
AND2x2_ASAP7_75t_L g607 ( .A(n_476), .B(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g612 ( .A(n_476), .B(n_570), .Y(n_612) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g569 ( .A(n_477), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g585 ( .A(n_477), .Y(n_585) );
AND2x2_ASAP7_75t_L g618 ( .A(n_477), .B(n_490), .Y(n_618) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_484), .B(n_489), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_483), .B(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_484) );
INVx2_ASAP7_75t_L g502 ( .A(n_490), .Y(n_502) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_490), .Y(n_587) );
INVx1_ASAP7_75t_L g606 ( .A(n_490), .Y(n_606) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_490), .Y(n_675) );
INVx1_ASAP7_75t_L g687 ( .A(n_490), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI31xp33_ASAP7_75t_SL g741 ( .A1(n_499), .A2(n_742), .A3(n_743), .B(n_744), .Y(n_741) );
NOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g666 ( .A(n_501), .B(n_568), .Y(n_666) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g582 ( .A(n_502), .Y(n_582) );
AND2x4_ASAP7_75t_SL g702 ( .A(n_504), .B(n_606), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_505), .A2(n_623), .B(n_626), .Y(n_622) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
INVx2_ASAP7_75t_L g595 ( .A(n_506), .Y(n_595) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2x1p5_ASAP7_75t_L g722 ( .A(n_507), .B(n_630), .Y(n_722) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g632 ( .A(n_508), .B(n_538), .Y(n_632) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVxp67_ASAP7_75t_L g557 ( .A(n_509), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_509), .B(n_518), .Y(n_592) );
AND2x4_ASAP7_75t_L g602 ( .A(n_509), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g647 ( .A(n_509), .B(n_539), .Y(n_647) );
INVx2_ASAP7_75t_L g655 ( .A(n_509), .Y(n_655) );
INVx1_ASAP7_75t_L g754 ( .A(n_509), .Y(n_754) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_509), .Y(n_763) );
INVx1_ASAP7_75t_L g700 ( .A(n_515), .Y(n_700) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_516), .B(n_529), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g556 ( .A(n_517), .B(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g695 ( .A(n_517), .B(n_630), .Y(n_695) );
AND2x2_ASAP7_75t_L g712 ( .A(n_517), .B(n_530), .Y(n_712) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_518), .B(n_560), .Y(n_735) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_528), .Y(n_518) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_519), .A2(n_520), .B(n_528), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_521), .B(n_527), .Y(n_520) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g658 ( .A(n_529), .B(n_556), .Y(n_658) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_538), .Y(n_529) );
INVx2_ASAP7_75t_L g564 ( .A(n_530), .Y(n_564) );
NOR2xp67_ASAP7_75t_L g745 ( .A(n_530), .B(n_538), .Y(n_745) );
NOR2x1_ASAP7_75t_L g753 ( .A(n_530), .B(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g661 ( .A(n_538), .B(n_565), .Y(n_661) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_539), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g590 ( .A(n_539), .Y(n_590) );
AND2x4_ASAP7_75t_L g654 ( .A(n_539), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g684 ( .A(n_539), .Y(n_684) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_547), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_551), .B1(n_552), .B2(n_553), .Y(n_547) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g705 ( .A1(n_555), .A2(n_568), .B1(n_706), .B2(n_707), .C(n_708), .Y(n_705) );
NAND2x1p5_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
AND2x2_ASAP7_75t_L g682 ( .A(n_556), .B(n_683), .Y(n_682) );
BUFx2_ASAP7_75t_L g725 ( .A(n_556), .Y(n_725) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g668 ( .A(n_559), .B(n_592), .Y(n_668) );
INVx3_ASAP7_75t_L g630 ( .A(n_560), .Y(n_630) );
AND2x2_ASAP7_75t_L g762 ( .A(n_560), .B(n_763), .Y(n_762) );
NAND3xp33_ASAP7_75t_SL g561 ( .A(n_562), .B(n_593), .C(n_609), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .B1(n_583), .B2(n_588), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_563), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g693 ( .A(n_563), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g704 ( .A(n_563), .B(n_599), .Y(n_704) );
AND2x2_ASAP7_75t_L g774 ( .A(n_563), .B(n_647), .Y(n_774) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g603 ( .A(n_565), .Y(n_603) );
INVx1_ASAP7_75t_L g652 ( .A(n_565), .Y(n_652) );
INVxp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI222xp33_ASAP7_75t_L g719 ( .A1(n_567), .A2(n_720), .B1(n_721), .B2(n_723), .C1(n_724), .C2(n_726), .Y(n_719) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_581), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_568), .B(n_595), .Y(n_594) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_568), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g686 ( .A(n_569), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g742 ( .A(n_569), .B(n_616), .Y(n_742) );
INVx2_ASAP7_75t_L g608 ( .A(n_570), .Y(n_608) );
INVx1_ASAP7_75t_L g620 ( .A(n_570), .Y(n_620) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_570), .Y(n_677) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_576), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .C(n_575), .Y(n_572) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_582), .Y(n_625) );
INVx3_ASAP7_75t_L g644 ( .A(n_582), .Y(n_644) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g710 ( .A(n_584), .Y(n_710) );
NAND2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g697 ( .A(n_586), .Y(n_697) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g698 ( .A(n_589), .Y(n_698) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g599 ( .A(n_590), .Y(n_599) );
AND2x2_ASAP7_75t_L g717 ( .A(n_590), .B(n_602), .Y(n_717) );
AND2x2_ASAP7_75t_L g780 ( .A(n_590), .B(n_712), .Y(n_780) );
AND2x2_ASAP7_75t_L g709 ( .A(n_591), .B(n_629), .Y(n_709) );
INVx1_ASAP7_75t_L g720 ( .A(n_591), .Y(n_720) );
AND2x2_ASAP7_75t_L g737 ( .A(n_591), .B(n_684), .Y(n_737) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .B1(n_600), .B2(n_604), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g609 ( .A1(n_596), .A2(n_610), .B(n_613), .Y(n_609) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g641 ( .A(n_599), .B(n_602), .Y(n_641) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g744 ( .A(n_602), .B(n_745), .Y(n_744) );
BUFx2_ASAP7_75t_L g707 ( .A(n_605), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_606), .Y(n_635) );
AND2x2_ASAP7_75t_SL g615 ( .A(n_607), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g680 ( .A(n_607), .Y(n_680) );
AND2x2_ASAP7_75t_L g778 ( .A(n_607), .B(n_675), .Y(n_778) );
INVx1_ASAP7_75t_L g733 ( .A(n_608), .Y(n_733) );
INVx1_ASAP7_75t_L g639 ( .A(n_610), .Y(n_639) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g728 ( .A(n_611), .Y(n_728) );
INVx4_ASAP7_75t_L g637 ( .A(n_612), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI32xp33_ASAP7_75t_L g708 ( .A1(n_615), .A2(n_709), .A3(n_710), .B1(n_711), .B2(n_712), .Y(n_708) );
AND2x2_ASAP7_75t_L g703 ( .A(n_616), .B(n_618), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_SL g766 ( .A1(n_616), .A2(n_767), .B(n_768), .C(n_770), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_SL g731 ( .A(n_618), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g770 ( .A(n_618), .Y(n_770) );
AND2x2_ASAP7_75t_L g624 ( .A(n_619), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g751 ( .A(n_619), .Y(n_751) );
AND2x2_ASAP7_75t_L g757 ( .A(n_619), .B(n_644), .Y(n_757) );
NOR3x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_638), .C(n_656), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_633), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
AND2x2_ASAP7_75t_L g646 ( .A(n_629), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g689 ( .A(n_629), .B(n_654), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_629), .B(n_675), .Y(n_716) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_637), .B(n_644), .Y(n_743) );
INVx2_ASAP7_75t_L g765 ( .A(n_637), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_642), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_639), .A2(n_730), .B1(n_734), .B2(n_736), .C(n_741), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_640), .A2(n_760), .B1(n_761), .B2(n_764), .Y(n_759) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_648), .B2(n_650), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g688 ( .A(n_644), .B(n_664), .Y(n_688) );
INVx1_ASAP7_75t_L g694 ( .A(n_644), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_644), .B(n_662), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_647), .B(n_715), .Y(n_781) );
NAND2x1_ASAP7_75t_L g764 ( .A(n_648), .B(n_765), .Y(n_764) );
INVx2_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_649), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2x1_ASAP7_75t_SL g767 ( .A(n_652), .B(n_654), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_652), .B(n_752), .Y(n_773) );
OR2x2_ASAP7_75t_L g734 ( .A(n_653), .B(n_735), .Y(n_734) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g769 ( .A(n_654), .B(n_695), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_657), .B(n_663), .Y(n_656) );
OAI21xp33_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_659), .B(n_662), .Y(n_657) );
OR2x2_ASAP7_75t_L g721 ( .A(n_660), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g755 ( .A(n_661), .B(n_753), .Y(n_755) );
AND2x2_ASAP7_75t_SL g701 ( .A(n_662), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g711 ( .A(n_662), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_667), .Y(n_663) );
AND2x2_ASAP7_75t_L g696 ( .A(n_664), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_713), .Y(n_670) );
NOR3xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_690), .C(n_705), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_678), .B(n_681), .C(n_685), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g739 ( .A(n_684), .Y(n_739) );
AND2x2_ASAP7_75t_L g752 ( .A(n_684), .B(n_753), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g760 ( .A(n_686), .Y(n_760) );
OAI21xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_698), .B(n_699), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_695), .B2(n_696), .Y(n_691) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_692), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_703), .B2(n_704), .Y(n_699) );
INVx1_ASAP7_75t_SL g706 ( .A(n_704), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_710), .B(n_751), .Y(n_750) );
OAI22xp33_ASAP7_75t_SL g776 ( .A1(n_711), .A2(n_777), .B1(n_779), .B2(n_781), .Y(n_776) );
AOI211x1_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_718), .B(n_719), .C(n_729), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_731), .A2(n_772), .B(n_774), .Y(n_771) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g740 ( .A(n_735), .Y(n_740) );
NOR2xp67_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_738), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_758), .C(n_771), .D(n_775), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_756), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_766), .Y(n_758) );
INVxp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx4_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
INVx3_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
INVx3_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_805), .B(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_SL g805 ( .A(n_806), .B(n_807), .Y(n_805) );
endmodule