module fake_jpeg_196_n_415 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_415);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_415;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_45),
.A2(n_37),
.B1(n_29),
.B2(n_26),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_48),
.Y(n_134)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_50),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_13),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_53),
.B(n_59),
.Y(n_139)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_10),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx12f_ASAP7_75t_SL g68 ( 
.A(n_23),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_79),
.Y(n_143)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_82),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_11),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_86),
.Y(n_122)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx16f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_89),
.Y(n_147)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_9),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_21),
.B(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_90),
.B(n_0),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_18),
.B(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_1),
.Y(n_150)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_96),
.Y(n_125)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_34),
.B1(n_40),
.B2(n_43),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_97),
.A2(n_100),
.B1(n_129),
.B2(n_74),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_34),
.B1(n_40),
.B2(n_43),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_21),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_48),
.B(n_38),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_127),
.B(n_86),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_34),
.B1(n_41),
.B2(n_18),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_146),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_43),
.B1(n_40),
.B2(n_38),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_117),
.A2(n_124),
.B1(n_146),
.B2(n_114),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_47),
.B(n_18),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_80),
.A2(n_37),
.B1(n_29),
.B2(n_26),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_123),
.A2(n_137),
.B1(n_149),
.B2(n_72),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_54),
.B(n_9),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_39),
.B1(n_1),
.B2(n_3),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_95),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_56),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_65),
.B(n_5),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_154),
.B(n_161),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_155),
.A2(n_165),
.B1(n_168),
.B2(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_122),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_157),
.B(n_170),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_158),
.B(n_167),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_160),
.B(n_180),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_75),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_101),
.A2(n_49),
.B1(n_66),
.B2(n_85),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_47),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_171),
.B(n_174),
.Y(n_219)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_71),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_81),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_175),
.B(n_178),
.Y(n_223)
);

OR2x2_ASAP7_75t_SL g176 ( 
.A(n_101),
.B(n_67),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_58),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_189),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_51),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_67),
.B(n_50),
.C(n_51),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_185),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_125),
.A2(n_78),
.B1(n_81),
.B2(n_50),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_103),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_188),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_107),
.B(n_7),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_98),
.B(n_8),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_115),
.B(n_140),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_117),
.Y(n_211)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_196),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_97),
.A2(n_100),
.B1(n_129),
.B2(n_123),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_198),
.B1(n_199),
.B2(n_104),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_195),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_121),
.B(n_110),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_104),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_197),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_144),
.A2(n_137),
.B1(n_133),
.B2(n_114),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_160),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_210),
.B(n_222),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_232),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_231),
.B1(n_157),
.B2(n_197),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_152),
.B1(n_110),
.B2(n_118),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_214),
.A2(n_218),
.B1(n_185),
.B2(n_170),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_182),
.A2(n_152),
.B1(n_118),
.B2(n_128),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_166),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_190),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_149),
.B1(n_142),
.B2(n_128),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_142),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_177),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_245),
.C(n_250),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_164),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_236),
.B(n_240),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_154),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_163),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_242),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_178),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_243),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_213),
.A2(n_159),
.B1(n_199),
.B2(n_194),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_249),
.B1(n_251),
.B2(n_257),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_184),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_191),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_217),
.A2(n_155),
.B1(n_181),
.B2(n_173),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_176),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_162),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_253),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_156),
.B1(n_192),
.B2(n_179),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_214),
.B1(n_218),
.B2(n_222),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_219),
.B(n_187),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_211),
.A2(n_195),
.B1(n_179),
.B2(n_186),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_172),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_193),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_204),
.A2(n_195),
.B1(n_99),
.B2(n_136),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_209),
.B1(n_225),
.B2(n_230),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_262),
.A2(n_269),
.B1(n_257),
.B2(n_258),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_252),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_265),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_259),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_274),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_216),
.B(n_209),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_268),
.A2(n_279),
.B(n_282),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_251),
.A2(n_237),
.B1(n_248),
.B2(n_244),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_260),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_275),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_236),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_241),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_247),
.A2(n_220),
.B(n_225),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_216),
.B1(n_215),
.B2(n_225),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_280),
.A2(n_242),
.B1(n_253),
.B2(n_238),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_255),
.A2(n_210),
.B(n_227),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_250),
.A2(n_227),
.B(n_200),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_234),
.B(n_224),
.Y(n_302)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_300),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_281),
.B(n_245),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_290),
.B(n_294),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_292),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_267),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_235),
.C(n_239),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_297),
.C(n_301),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_268),
.B(n_261),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_295),
.A2(n_284),
.B1(n_274),
.B2(n_283),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_200),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_299),
.A2(n_303),
.B1(n_270),
.B2(n_278),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_221),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_234),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_269),
.A2(n_201),
.B1(n_228),
.B2(n_224),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_263),
.A2(n_201),
.B1(n_228),
.B2(n_221),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_262),
.B1(n_295),
.B2(n_287),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_273),
.B(n_202),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_308),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_280),
.C(n_279),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_284),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_286),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_323),
.B1(n_325),
.B2(n_329),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_322),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_327),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_321),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_266),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_296),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_332),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_283),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_326),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_272),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_328),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_299),
.A2(n_284),
.B1(n_275),
.B2(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_331),
.Y(n_350)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_296),
.B1(n_308),
.B2(n_288),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_333),
.A2(n_342),
.B1(n_351),
.B2(n_315),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_324),
.A2(n_309),
.B(n_302),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_338),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_301),
.C(n_294),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_310),
.B(n_327),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_169),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_332),
.A2(n_305),
.B1(n_297),
.B2(n_303),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_272),
.Y(n_343)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_343),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_323),
.A2(n_272),
.B1(n_270),
.B2(n_278),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_345),
.A2(n_314),
.B1(n_312),
.B2(n_320),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_282),
.C(n_212),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_169),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_233),
.Y(n_349)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_314),
.A2(n_233),
.B1(n_202),
.B2(n_111),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_344),
.B(n_311),
.Y(n_352)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_354),
.A2(n_341),
.B1(n_340),
.B2(n_366),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_347),
.B(n_317),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_363),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_350),
.A2(n_329),
.B1(n_321),
.B2(n_320),
.Y(n_356)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_356),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_357),
.Y(n_374)
);

INVx13_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_358),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_350),
.A2(n_315),
.B1(n_310),
.B2(n_233),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_359),
.B(n_364),
.Y(n_369)
);

AOI21xp33_ASAP7_75t_L g376 ( 
.A1(n_361),
.A2(n_337),
.B(n_334),
.Y(n_376)
);

NAND4xp25_ASAP7_75t_SL g362 ( 
.A(n_349),
.B(n_169),
.C(n_148),
.D(n_136),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_362),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_333),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_148),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_338),
.C(n_346),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_356),
.A2(n_340),
.B(n_336),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_376),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_348),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_353),
.C(n_355),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_382),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_365),
.Y(n_380)
);

AOI21xp33_ASAP7_75t_L g392 ( 
.A1(n_380),
.A2(n_386),
.B(n_388),
.Y(n_392)
);

INVx11_ASAP7_75t_L g383 ( 
.A(n_377),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_384),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_359),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_372),
.B(n_360),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_374),
.B(n_343),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_389),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_372),
.B(n_341),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_385),
.A2(n_368),
.B(n_369),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_391),
.A2(n_335),
.B(n_345),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_374),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_394),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_371),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_373),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_395),
.B(n_369),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_397),
.B(n_371),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_398),
.B(n_399),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_388),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_390),
.C(n_392),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_396),
.A2(n_354),
.B1(n_358),
.B2(n_367),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_402),
.Y(n_406)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_405),
.Y(n_409)
);

O2A1O1Ixp33_ASAP7_75t_SL g407 ( 
.A1(n_400),
.A2(n_377),
.B(n_339),
.C(n_351),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_402),
.B(n_403),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_408),
.A2(n_410),
.B(n_406),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_404),
.B(n_377),
.C(n_362),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_409),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_411),
.A2(n_412),
.B(n_377),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_413),
.B(n_105),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_105),
.Y(n_415)
);


endmodule