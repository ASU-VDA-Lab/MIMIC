module real_jpeg_7848_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_0),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_0),
.A2(n_1),
.B1(n_27),
.B2(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_1),
.A2(n_31),
.B(n_32),
.C(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_4),
.A2(n_20),
.B1(n_23),
.B2(n_55),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_4),
.A2(n_8),
.B(n_20),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_6),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_5),
.A2(n_28),
.B(n_38),
.C(n_42),
.Y(n_41)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_5),
.B(n_28),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_5),
.A2(n_6),
.A3(n_28),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_6),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_6),
.B(n_55),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_8),
.B1(n_24),
.B2(n_40),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_6),
.A2(n_24),
.B(n_55),
.C(n_83),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g29 ( 
.A(n_7),
.B(n_24),
.CON(n_29),
.SN(n_29)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_28),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_8),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_38),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_77),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_76),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_66),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_13),
.B(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_65),
.Y(n_13)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_34),
.B2(n_35),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_25),
.B2(n_33),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_17),
.A2(n_18),
.B1(n_45),
.B2(n_46),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_17),
.A2(n_18),
.B1(n_85),
.B2(n_88),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_17),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_17),
.A2(n_18),
.B1(n_73),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_36),
.C(n_45),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_18),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_18),
.B(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_18),
.B(n_53),
.C(n_86),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_21),
.B(n_22),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_21),
.B(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_23),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_24),
.B(n_57),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_29),
.B(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_59),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_40),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_51),
.A2(n_63),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_53),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_53),
.B1(n_82),
.B2(n_98),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_59),
.B(n_105),
.C(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_59),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_52),
.A2(n_53),
.B1(n_71),
.B2(n_72),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_67),
.C(n_71),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_57),
.B(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_67),
.A2(n_68),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_73),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_107),
.B(n_114),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_100),
.B(n_106),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_99),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_84),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);


endmodule