module fake_jpeg_9353_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_28),
.B1(n_32),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_58),
.B1(n_16),
.B2(n_18),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_28),
.B1(n_32),
.B2(n_29),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_64),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_27),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_32),
.B1(n_29),
.B2(n_26),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_16),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_69),
.B(n_73),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_45),
.B1(n_38),
.B2(n_39),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_95),
.B1(n_20),
.B2(n_18),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_29),
.B1(n_33),
.B2(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_84),
.B1(n_88),
.B2(n_20),
.Y(n_112)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_83),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_78),
.A2(n_79),
.B1(n_51),
.B2(n_60),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_47),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_17),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_81),
.B(n_90),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_25),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_17),
.B1(n_33),
.B2(n_25),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_91),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_17),
.B1(n_33),
.B2(n_31),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_16),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_27),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_0),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_122),
.B1(n_127),
.B2(n_89),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_53),
.C(n_45),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_117),
.C(n_119),
.Y(n_149)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_109),
.Y(n_152)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_121),
.B1(n_89),
.B2(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_93),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_51),
.B1(n_60),
.B2(n_53),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_74),
.B1(n_99),
.B2(n_79),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_38),
.C(n_54),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_54),
.C(n_56),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_73),
.A2(n_75),
.B1(n_84),
.B2(n_92),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_13),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_100),
.Y(n_159)
);

XOR2x2_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_31),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_95),
.B(n_90),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_81),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_56),
.C(n_47),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_85),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_142),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_90),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_133),
.A2(n_135),
.B(n_148),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_70),
.B(n_59),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_140),
.A2(n_144),
.B(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_70),
.Y(n_141)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_121),
.B(n_88),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_102),
.B1(n_105),
.B2(n_108),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_101),
.A2(n_59),
.B1(n_74),
.B2(n_99),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_160),
.B1(n_114),
.B2(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_155),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_22),
.B(n_26),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_0),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_96),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_150),
.C(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_158),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_96),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_119),
.B1(n_110),
.B2(n_100),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_107),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_15),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_169),
.B1(n_178),
.B2(n_147),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_160),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_173),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_167),
.B(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_155),
.A2(n_104),
.B1(n_107),
.B2(n_105),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_181),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_131),
.Y(n_171)
);

CKINVDCx10_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_85),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_131),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_174),
.B(n_177),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_190),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_176),
.A2(n_185),
.B1(n_1),
.B2(n_2),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_102),
.B1(n_87),
.B2(n_24),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_138),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_24),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_129),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_188),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_130),
.B(n_109),
.C(n_23),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_23),
.B1(n_30),
.B2(n_19),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_146),
.B1(n_161),
.B2(n_19),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_195),
.A2(n_220),
.B1(n_181),
.B2(n_162),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_144),
.B1(n_134),
.B2(n_140),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_205),
.B1(n_208),
.B2(n_179),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_182),
.A2(n_135),
.B1(n_132),
.B2(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_201),
.B(n_211),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_158),
.B1(n_157),
.B2(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_153),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_1),
.B(n_3),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_151),
.B1(n_142),
.B2(n_143),
.Y(n_204)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_143),
.B1(n_148),
.B2(n_30),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_148),
.B1(n_22),
.B2(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_210),
.Y(n_240)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_215),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_221),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_219),
.A2(n_223),
.B(n_165),
.Y(n_231)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_1),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_224),
.A2(n_234),
.B1(n_245),
.B2(n_246),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_168),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_225),
.B(n_237),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_166),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_204),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_230),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_170),
.B1(n_177),
.B2(n_162),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_214),
.A2(n_163),
.B1(n_175),
.B2(n_164),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_195),
.A2(n_167),
.B1(n_164),
.B2(n_186),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_197),
.A2(n_190),
.B1(n_186),
.B2(n_168),
.Y(n_236)
);

XNOR2x2_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_173),
.Y(n_237)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_239),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_223),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_208),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_202),
.A2(n_3),
.B(n_5),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_212),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_199),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_196),
.C(n_222),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_252),
.C(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_222),
.C(n_210),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_259),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_209),
.C(n_203),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_203),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_217),
.C(n_205),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_264),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_245),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_213),
.C(n_207),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_11),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_241),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_11),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_247),
.B(n_246),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_269),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_244),
.B1(n_227),
.B2(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_253),
.A2(n_227),
.B1(n_242),
.B2(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_226),
.B(n_231),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_258),
.B(n_259),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_224),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_282),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_242),
.B1(n_267),
.B2(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_286),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_295),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_298),
.Y(n_312)
);

NOR4xp25_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_266),
.C(n_249),
.D(n_270),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_277),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_251),
.B(n_282),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_257),
.B(n_251),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_272),
.B(n_279),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_12),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_306),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_8),
.C2(n_5),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_303),
.B(n_304),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_232),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_284),
.C(n_280),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_309),
.C(n_13),
.Y(n_316)
);

AOI21x1_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_280),
.B(n_284),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_11),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_15),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_9),
.C(n_14),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_300),
.B1(n_289),
.B2(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_319),
.Y(n_322)
);

AOI31xp67_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_320),
.A3(n_321),
.B(n_8),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_6),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_302),
.A2(n_6),
.B(n_7),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_6),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_315),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_324),
.B(n_325),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_308),
.B(n_312),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_327),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_328),
.C(n_322),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_330),
.C(n_317),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_8),
.Y(n_334)
);


endmodule