module fake_ibex_1114_n_921 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_921);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_921;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_433;
wire n_262;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_206;
wire n_179;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_285;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_298;
wire n_231;
wire n_202;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_9),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_19),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

BUFx2_ASAP7_75t_SL g181 ( 
.A(n_50),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_37),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_26),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_55),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_32),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_92),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_67),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_63),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_44),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_70),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_54),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_53),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_57),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_76),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_77),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_19),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_21),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_164),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_33),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_30),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_117),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_129),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_64),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_140),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_46),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_82),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_105),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_147),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_51),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_48),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_119),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_95),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_22),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_71),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_99),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_69),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_22),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_78),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_37),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_145),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_134),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_91),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_52),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_66),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_100),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_79),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_143),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_26),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_72),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_125),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_8),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_2),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_59),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_155),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_0),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_49),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_86),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_165),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_38),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_35),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_45),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_133),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_39),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_18),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_56),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_94),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_131),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_120),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_16),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_21),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_43),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_146),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_154),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_30),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_41),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_80),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_132),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_29),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_191),
.B(n_0),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_199),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_210),
.B(n_1),
.Y(n_282)
);

AOI22x1_ASAP7_75t_SL g283 ( 
.A1(n_170),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_217),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_175),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_175),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_182),
.B(n_40),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_221),
.B(n_4),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_221),
.B(n_5),
.Y(n_291)
);

AOI22x1_ASAP7_75t_SL g292 ( 
.A1(n_170),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_182),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_6),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_268),
.B(n_10),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_11),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_172),
.B(n_42),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_190),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g302 ( 
.A(n_172),
.B(n_47),
.Y(n_302)
);

OA21x2_ASAP7_75t_L g303 ( 
.A1(n_190),
.A2(n_88),
.B(n_163),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_192),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_184),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_192),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_206),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_171),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_200),
.B(n_11),
.Y(n_310)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_200),
.B(n_58),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_197),
.B(n_60),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_223),
.B(n_12),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_177),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_197),
.B(n_13),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_14),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_213),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_218),
.B(n_15),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_216),
.B(n_16),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_216),
.B(n_17),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_177),
.B(n_17),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_169),
.A2(n_93),
.B(n_161),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_186),
.Y(n_323)
);

AOI22x1_ASAP7_75t_SL g324 ( 
.A1(n_186),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_229),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_20),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_235),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_199),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_250),
.B(n_23),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_176),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_251),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_257),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_178),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_171),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_261),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_227),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_24),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_180),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_24),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_264),
.B(n_25),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_227),
.Y(n_343)
);

CKINVDCx11_ASAP7_75t_R g344 ( 
.A(n_255),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_265),
.Y(n_345)
);

BUFx8_ASAP7_75t_L g346 ( 
.A(n_183),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_187),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_271),
.Y(n_348)
);

CKINVDCx8_ASAP7_75t_R g349 ( 
.A(n_181),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_193),
.Y(n_350)
);

OAI21x1_ASAP7_75t_L g351 ( 
.A1(n_195),
.A2(n_98),
.B(n_160),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_199),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_201),
.B(n_25),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_203),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_281),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_337),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_284),
.B(n_173),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_294),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_284),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_304),
.B(n_173),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_174),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_344),
.Y(n_367)
);

BUFx10_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g369 ( 
.A(n_287),
.B(n_208),
.C(n_205),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_310),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_294),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_321),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_349),
.B(n_174),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_310),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_185),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_315),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_266),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_309),
.B(n_209),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_306),
.B(n_215),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_346),
.B(n_188),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_346),
.B(n_188),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_353),
.B(n_256),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_298),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_298),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_319),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_282),
.B(n_290),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_353),
.B(n_258),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_280),
.B(n_297),
.C(n_353),
.Y(n_392)
);

NOR2x1p5_ASAP7_75t_L g393 ( 
.A(n_338),
.B(n_253),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_308),
.B(n_222),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_326),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_320),
.B(n_259),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_320),
.B(n_260),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_291),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_331),
.B(n_260),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_320),
.B(n_263),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_299),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_317),
.B(n_224),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_334),
.B(n_340),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_330),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_339),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_325),
.B(n_225),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_286),
.Y(n_417)
);

INVx8_ASAP7_75t_L g418 ( 
.A(n_299),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_334),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_303),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_327),
.B(n_329),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_L g422 ( 
.A(n_299),
.B(n_302),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_340),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_303),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_286),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_309),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_332),
.B(n_333),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_336),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_288),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_345),
.B(n_269),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_288),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_313),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_301),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_348),
.B(n_274),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_293),
.B(n_228),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_301),
.B(n_274),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_305),
.B(n_276),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_305),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_307),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_307),
.B(n_276),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_295),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_299),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_300),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_312),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_318),
.B(n_194),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_341),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_312),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_302),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_312),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_318),
.B(n_196),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_296),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_312),
.Y(n_453)
);

INVxp33_ASAP7_75t_L g454 ( 
.A(n_344),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_365),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_372),
.B(n_342),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_449),
.B(n_342),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_434),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_357),
.B(n_316),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_449),
.B(n_316),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_L g463 ( 
.A1(n_398),
.A2(n_285),
.B1(n_314),
.B2(n_335),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_364),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_409),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_302),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_418),
.B(n_302),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_398),
.B(n_338),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_366),
.B(n_343),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_359),
.A2(n_302),
.B1(n_311),
.B2(n_312),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_429),
.B(n_311),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_366),
.B(n_311),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_362),
.B(n_343),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_412),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_365),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_356),
.A2(n_296),
.B1(n_311),
.B2(n_324),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_375),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_356),
.B(n_289),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_204),
.Y(n_482)
);

AO22x2_ASAP7_75t_L g483 ( 
.A1(n_392),
.A2(n_283),
.B1(n_292),
.B2(n_267),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_390),
.B(n_207),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_368),
.B(n_211),
.Y(n_485)
);

O2A1O1Ixp33_ASAP7_75t_L g486 ( 
.A1(n_358),
.A2(n_244),
.B(n_245),
.C(n_278),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_390),
.B(n_212),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_368),
.B(n_214),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_374),
.B(n_220),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_444),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_418),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_362),
.B(n_230),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_L g493 ( 
.A(n_443),
.B(n_234),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_406),
.B(n_428),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_363),
.B(n_179),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_446),
.B(n_231),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_452),
.B(n_236),
.Y(n_497)
);

OAI221xp5_ASAP7_75t_L g498 ( 
.A1(n_433),
.A2(n_202),
.B1(n_246),
.B2(n_272),
.C(n_262),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_421),
.B(n_237),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_404),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_404),
.B(n_240),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

OR2x6_ASAP7_75t_SL g503 ( 
.A(n_379),
.B(n_241),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_239),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

NOR3xp33_ASAP7_75t_L g506 ( 
.A(n_369),
.B(n_198),
.C(n_226),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_374),
.B(n_242),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_378),
.B(n_243),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_417),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_433),
.B(n_232),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_401),
.B(n_248),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_385),
.B(n_273),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_402),
.A2(n_277),
.B1(n_254),
.B2(n_252),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_414),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_426),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_414),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_407),
.B(n_249),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_391),
.B(n_322),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_425),
.B(n_322),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_426),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_430),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_360),
.B(n_351),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_374),
.B(n_97),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_371),
.B(n_27),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_420),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_381),
.B(n_28),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_389),
.B(n_28),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_370),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_431),
.B(n_102),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_370),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_396),
.B(n_359),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_367),
.B(n_34),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_432),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_359),
.A2(n_36),
.B1(n_61),
.B2(n_62),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_377),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_377),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_377),
.A2(n_36),
.B1(n_65),
.B2(n_68),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_386),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_386),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_382),
.B(n_74),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_464),
.B(n_373),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_464),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_475),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_519),
.A2(n_422),
.B(n_453),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_L g548 ( 
.A(n_478),
.B(n_384),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_537),
.Y(n_549)
);

CKINVDCx14_ASAP7_75t_R g550 ( 
.A(n_503),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_523),
.A2(n_422),
.B(n_450),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_455),
.A2(n_393),
.B1(n_435),
.B2(n_437),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_494),
.B(n_380),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_460),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_491),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_479),
.B(n_394),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_465),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_468),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_491),
.B(n_445),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_518),
.A2(n_450),
.B(n_448),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_480),
.B(n_410),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_476),
.B(n_454),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_481),
.B(n_456),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_466),
.A2(n_424),
.B(n_420),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_465),
.Y(n_565)
);

CKINVDCx10_ASAP7_75t_R g566 ( 
.A(n_483),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_471),
.A2(n_441),
.B(n_438),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_472),
.A2(n_424),
.B(n_420),
.Y(n_568)
);

A2O1A1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_461),
.A2(n_486),
.B(n_538),
.C(n_540),
.Y(n_569)
);

O2A1O1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_498),
.A2(n_416),
.B(n_439),
.C(n_436),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_467),
.A2(n_424),
.B(n_420),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_533),
.A2(n_424),
.B(n_440),
.Y(n_572)
);

OAI21xp33_ASAP7_75t_L g573 ( 
.A1(n_481),
.A2(n_379),
.B(n_424),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_461),
.B(n_411),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_473),
.A2(n_376),
.B(n_411),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_510),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_534),
.B(n_81),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_469),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_500),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_482),
.B(n_427),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_462),
.A2(n_376),
.B(n_408),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_484),
.B(n_487),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_474),
.B(n_427),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_541),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_496),
.B(n_504),
.Y(n_585)
);

AO21x1_ASAP7_75t_L g586 ( 
.A1(n_524),
.A2(n_405),
.B(n_403),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_501),
.B(n_83),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_471),
.A2(n_388),
.B(n_403),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_492),
.B(n_84),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_529),
.B(n_85),
.Y(n_590)
);

O2A1O1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_463),
.A2(n_400),
.B(n_399),
.C(n_397),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_492),
.B(n_87),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_463),
.B(n_499),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_457),
.A2(n_388),
.B(n_400),
.Y(n_594)
);

AOI21x1_ASAP7_75t_L g595 ( 
.A1(n_514),
.A2(n_516),
.B(n_543),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_525),
.A2(n_387),
.B(n_399),
.Y(n_596)
);

A2O1A1Ixp33_ASAP7_75t_L g597 ( 
.A1(n_522),
.A2(n_383),
.B(n_397),
.C(n_395),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_527),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_528),
.A2(n_383),
.B(n_395),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_531),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_512),
.B(n_89),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_495),
.B(n_90),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_483),
.B(n_101),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_477),
.B(n_104),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_490),
.B(n_108),
.Y(n_605)
);

O2A1O1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_506),
.A2(n_361),
.B(n_355),
.C(n_111),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_458),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_459),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_483),
.B(n_109),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_502),
.B(n_110),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_506),
.B(n_112),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_508),
.B(n_511),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_517),
.B(n_114),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_513),
.B(n_115),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_521),
.A2(n_413),
.B(n_116),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_505),
.A2(n_413),
.B(n_118),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_532),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_470),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_509),
.A2(n_413),
.B(n_126),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_485),
.B(n_121),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_515),
.B(n_520),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_535),
.A2(n_413),
.B(n_139),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_521),
.A2(n_166),
.B(n_141),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_530),
.A2(n_144),
.B(n_148),
.C(n_151),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_526),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_542),
.Y(n_626)
);

A2O1A1Ixp33_ASAP7_75t_L g627 ( 
.A1(n_497),
.A2(n_153),
.B(n_156),
.C(n_539),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_488),
.B(n_489),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_507),
.B(n_493),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_545),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_546),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_555),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_554),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_563),
.B(n_536),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_600),
.Y(n_635)
);

AO32x2_ASAP7_75t_L g636 ( 
.A1(n_554),
.A2(n_526),
.A3(n_536),
.B1(n_539),
.B2(n_591),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_553),
.B(n_556),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_569),
.A2(n_568),
.B(n_547),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_562),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_606),
.B(n_627),
.C(n_573),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_617),
.A2(n_593),
.B1(n_582),
.B2(n_585),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_558),
.B(n_576),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_551),
.A2(n_572),
.B(n_560),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_578),
.B(n_580),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_572),
.A2(n_574),
.B(n_612),
.Y(n_645)
);

AO31x2_ASAP7_75t_L g646 ( 
.A1(n_586),
.A2(n_624),
.A3(n_615),
.B(n_623),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_561),
.B(n_548),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_621),
.A2(n_567),
.B(n_575),
.Y(n_648)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_616),
.A2(n_622),
.B(n_619),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_579),
.B(n_583),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_544),
.B(n_552),
.Y(n_651)
);

OAI21x1_ASAP7_75t_SL g652 ( 
.A1(n_555),
.A2(n_629),
.B(n_602),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_625),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_615),
.A2(n_570),
.B(n_598),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_628),
.B(n_608),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_626),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_550),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_607),
.B(n_618),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_590),
.B(n_609),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_625),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_603),
.B(n_549),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_589),
.A2(n_592),
.B1(n_601),
.B2(n_577),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_588),
.A2(n_597),
.B(n_581),
.Y(n_664)
);

BUFx8_ASAP7_75t_L g665 ( 
.A(n_566),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_587),
.A2(n_614),
.B(n_620),
.C(n_611),
.Y(n_666)
);

OAI21x1_ASAP7_75t_SL g667 ( 
.A1(n_613),
.A2(n_595),
.B(n_604),
.Y(n_667)
);

AO31x2_ASAP7_75t_L g668 ( 
.A1(n_596),
.A2(n_599),
.A3(n_610),
.B(n_605),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_594),
.A2(n_599),
.B(n_559),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_565),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_565),
.A2(n_546),
.B1(n_553),
.B2(n_593),
.Y(n_671)
);

AND2x6_ASAP7_75t_L g672 ( 
.A(n_557),
.B(n_546),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_557),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_625),
.A2(n_449),
.B(n_627),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_563),
.B(n_546),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_563),
.B(n_546),
.Y(n_676)
);

AO31x2_ASAP7_75t_L g677 ( 
.A1(n_571),
.A2(n_627),
.A3(n_586),
.B(n_564),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_545),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_563),
.B(n_546),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_563),
.B(n_546),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_563),
.B(n_546),
.Y(n_681)
);

OA22x2_ASAP7_75t_L g682 ( 
.A1(n_558),
.A2(n_379),
.B1(n_338),
.B2(n_343),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_563),
.B(n_546),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_545),
.B(n_335),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_564),
.A2(n_422),
.B(n_467),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_554),
.Y(n_686)
);

NOR2xp67_ASAP7_75t_L g687 ( 
.A(n_555),
.B(n_546),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_569),
.A2(n_518),
.B(n_519),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_545),
.B(n_464),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_563),
.B(n_546),
.Y(n_690)
);

AO31x2_ASAP7_75t_L g691 ( 
.A1(n_571),
.A2(n_627),
.A3(n_586),
.B(n_564),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_555),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_555),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_563),
.B(n_546),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_563),
.B(n_546),
.Y(n_695)
);

NOR2x1_ASAP7_75t_SL g696 ( 
.A(n_555),
.B(n_546),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_612),
.A2(n_591),
.B(n_461),
.C(n_518),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_554),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_563),
.B(n_546),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_545),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_625),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_545),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_555),
.Y(n_703)
);

CKINVDCx6p67_ASAP7_75t_R g704 ( 
.A(n_566),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_569),
.A2(n_518),
.B(n_519),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_546),
.A2(n_553),
.B1(n_593),
.B2(n_563),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_612),
.A2(n_591),
.B(n_461),
.C(n_518),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_563),
.B(n_546),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_545),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_555),
.Y(n_710)
);

CKINVDCx6p67_ASAP7_75t_R g711 ( 
.A(n_566),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_593),
.B(n_464),
.Y(n_712)
);

BUFx2_ASAP7_75t_SL g713 ( 
.A(n_554),
.Y(n_713)
);

BUFx2_ASAP7_75t_L g714 ( 
.A(n_545),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_555),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_612),
.A2(n_591),
.B(n_461),
.C(n_518),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_697),
.A2(n_716),
.B(n_707),
.Y(n_717)
);

AO22x2_ASAP7_75t_L g718 ( 
.A1(n_706),
.A2(n_671),
.B1(n_660),
.B2(n_652),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_633),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_657),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_637),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_713),
.B(n_693),
.Y(n_722)
);

NOR2x1_ASAP7_75t_SL g723 ( 
.A(n_693),
.B(n_710),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_665),
.Y(n_724)
);

AO21x1_ASAP7_75t_L g725 ( 
.A1(n_654),
.A2(n_645),
.B(n_663),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_710),
.B(n_715),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_669),
.A2(n_638),
.B(n_685),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_642),
.B(n_689),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_712),
.A2(n_644),
.B1(n_682),
.B2(n_641),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_641),
.A2(n_650),
.B1(n_678),
.B2(n_714),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_675),
.A2(n_694),
.B1(n_679),
.B2(n_708),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_658),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_676),
.B(n_680),
.Y(n_733)
);

NAND2x1p5_ASAP7_75t_L g734 ( 
.A(n_715),
.B(n_670),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_681),
.A2(n_695),
.B1(n_683),
.B2(n_690),
.Y(n_735)
);

AOI21xp33_ASAP7_75t_L g736 ( 
.A1(n_654),
.A2(n_634),
.B(n_640),
.Y(n_736)
);

AO21x2_ASAP7_75t_L g737 ( 
.A1(n_643),
.A2(n_640),
.B(n_667),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_687),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_699),
.A2(n_666),
.B1(n_662),
.B2(n_635),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_688),
.B(n_705),
.C(n_647),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_700),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_709),
.B(n_651),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_630),
.B(n_702),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_655),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_704),
.A2(n_711),
.B1(n_684),
.B2(n_656),
.Y(n_745)
);

OAI21xp5_ASAP7_75t_L g746 ( 
.A1(n_648),
.A2(n_664),
.B(n_674),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_656),
.A2(n_659),
.B1(n_670),
.B2(n_703),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_639),
.B(n_698),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_673),
.Y(n_749)
);

AO31x2_ASAP7_75t_L g750 ( 
.A1(n_636),
.A2(n_677),
.A3(n_691),
.B(n_646),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_653),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_686),
.Y(n_752)
);

INVx3_ASAP7_75t_SL g753 ( 
.A(n_632),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_692),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_649),
.A2(n_701),
.B(n_661),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_672),
.A2(n_636),
.B(n_691),
.Y(n_756)
);

OAI21x1_ASAP7_75t_L g757 ( 
.A1(n_677),
.A2(n_691),
.B(n_646),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_672),
.B(n_653),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_701),
.B(n_653),
.Y(n_759)
);

AOI211xp5_ASAP7_75t_L g760 ( 
.A1(n_636),
.A2(n_661),
.B(n_701),
.C(n_646),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_668),
.A2(n_716),
.B(n_707),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_712),
.A2(n_583),
.B1(n_573),
.B2(n_617),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_641),
.A2(n_309),
.B1(n_343),
.B2(n_338),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_697),
.A2(n_716),
.B(n_707),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_637),
.B(n_696),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_637),
.B(n_464),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_SL g767 ( 
.A1(n_706),
.A2(n_309),
.B1(n_343),
.B2(n_338),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_637),
.B(n_464),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_637),
.B(n_455),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_706),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_637),
.B(n_641),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_693),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_706),
.A2(n_641),
.B1(n_637),
.B2(n_634),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_712),
.B(n_506),
.C(n_583),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_706),
.A2(n_641),
.B1(n_637),
.B2(n_634),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_SL g776 ( 
.A(n_706),
.B(n_670),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_637),
.B(n_455),
.Y(n_777)
);

CKINVDCx11_ASAP7_75t_R g778 ( 
.A(n_704),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_631),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_740),
.Y(n_780)
);

AND2x4_ASAP7_75t_SL g781 ( 
.A(n_722),
.B(n_765),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_SL g782 ( 
.A1(n_776),
.A2(n_770),
.B1(n_765),
.B2(n_726),
.Y(n_782)
);

BUFx12f_ASAP7_75t_L g783 ( 
.A(n_778),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_732),
.B(n_771),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_722),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_761),
.A2(n_727),
.B(n_757),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_722),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_739),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_774),
.A2(n_735),
.B(n_731),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_758),
.B(n_772),
.Y(n_790)
);

OAI21xp33_ASAP7_75t_L g791 ( 
.A1(n_767),
.A2(n_729),
.B(n_762),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_741),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_779),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_733),
.B(n_732),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_771),
.B(n_721),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_769),
.B(n_777),
.Y(n_796)
);

AO21x2_ASAP7_75t_L g797 ( 
.A1(n_746),
.A2(n_727),
.B(n_717),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_738),
.Y(n_798)
);

AO31x2_ASAP7_75t_L g799 ( 
.A1(n_725),
.A2(n_775),
.A3(n_773),
.B(n_755),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_772),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_773),
.B(n_775),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_719),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_738),
.B(n_734),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_767),
.A2(n_763),
.B1(n_742),
.B2(n_730),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_766),
.B(n_768),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_744),
.B(n_743),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_723),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_749),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_747),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_747),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_745),
.B(n_728),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_717),
.Y(n_812)
);

AO21x2_ASAP7_75t_L g813 ( 
.A1(n_764),
.A2(n_736),
.B(n_756),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_764),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_753),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_718),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_749),
.B(n_750),
.Y(n_817)
);

NAND4xp25_ASAP7_75t_SL g818 ( 
.A(n_724),
.B(n_752),
.C(n_760),
.D(n_754),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_750),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_781),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_781),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_798),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_797),
.B(n_756),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_819),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_797),
.B(n_737),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_798),
.Y(n_826)
);

BUFx2_ASAP7_75t_SL g827 ( 
.A(n_785),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_813),
.B(n_751),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_813),
.B(n_759),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_801),
.B(n_784),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_784),
.B(n_748),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_788),
.B(n_720),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_795),
.B(n_812),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_814),
.B(n_786),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_SL g835 ( 
.A1(n_789),
.A2(n_785),
.B1(n_787),
.B2(n_794),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_808),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_826),
.Y(n_837)
);

INVx5_ASAP7_75t_L g838 ( 
.A(n_820),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_823),
.B(n_809),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_823),
.B(n_809),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_824),
.Y(n_841)
);

NOR2x1_ASAP7_75t_SL g842 ( 
.A(n_820),
.B(n_803),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_823),
.B(n_810),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_834),
.B(n_810),
.Y(n_844)
);

NAND2x1p5_ASAP7_75t_L g845 ( 
.A(n_820),
.B(n_787),
.Y(n_845)
);

OR2x2_ASAP7_75t_SL g846 ( 
.A(n_822),
.B(n_817),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_834),
.B(n_816),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_836),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_834),
.B(n_816),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_825),
.B(n_799),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_833),
.B(n_780),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_839),
.B(n_828),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_848),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_840),
.B(n_830),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_841),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_851),
.B(n_836),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_843),
.B(n_825),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_843),
.B(n_829),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_851),
.B(n_830),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_844),
.B(n_847),
.Y(n_860)
);

OR2x6_ASAP7_75t_L g861 ( 
.A(n_845),
.B(n_820),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_860),
.B(n_857),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_858),
.B(n_837),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_860),
.B(n_844),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_857),
.B(n_847),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_852),
.B(n_849),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_853),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_854),
.B(n_846),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_852),
.B(n_850),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_855),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_855),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_867),
.B(n_835),
.C(n_856),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_870),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_863),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_864),
.B(n_865),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_868),
.A2(n_842),
.B(n_861),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_871),
.Y(n_877)
);

OAI32xp33_ASAP7_75t_L g878 ( 
.A1(n_862),
.A2(n_854),
.A3(n_845),
.B1(n_821),
.B2(n_859),
.Y(n_878)
);

OAI32xp33_ASAP7_75t_L g879 ( 
.A1(n_866),
.A2(n_845),
.A3(n_821),
.B1(n_822),
.B2(n_832),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_863),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_869),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_874),
.B(n_869),
.Y(n_882)
);

OAI221xp5_ASAP7_75t_L g883 ( 
.A1(n_872),
.A2(n_874),
.B1(n_876),
.B2(n_880),
.C(n_835),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_873),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_877),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_SL g886 ( 
.A1(n_883),
.A2(n_807),
.B(n_782),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_882),
.A2(n_879),
.B(n_878),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_882),
.B(n_881),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_887),
.B(n_783),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_888),
.B(n_884),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_890),
.B(n_886),
.Y(n_891)
);

NOR3x1_ASAP7_75t_L g892 ( 
.A(n_889),
.B(n_783),
.C(n_832),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_891),
.B(n_885),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_892),
.B(n_802),
.C(n_792),
.Y(n_894)
);

NAND4xp75_ASAP7_75t_L g895 ( 
.A(n_893),
.B(n_811),
.C(n_884),
.D(n_805),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_894),
.Y(n_896)
);

AOI22x1_ASAP7_75t_L g897 ( 
.A1(n_896),
.A2(n_815),
.B1(n_800),
.B2(n_875),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_895),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_896),
.A2(n_861),
.B1(n_804),
.B2(n_838),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_897),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_898),
.Y(n_901)
);

OR2x4_ASAP7_75t_L g902 ( 
.A(n_899),
.B(n_832),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_898),
.Y(n_903)
);

AO21x2_ASAP7_75t_L g904 ( 
.A1(n_898),
.A2(n_791),
.B(n_806),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_901),
.Y(n_905)
);

AOI31xp33_ASAP7_75t_L g906 ( 
.A1(n_901),
.A2(n_802),
.A3(n_790),
.B(n_796),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_903),
.A2(n_815),
.B(n_800),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_903),
.B(n_863),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_900),
.A2(n_904),
.B(n_902),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_901),
.A2(n_818),
.B1(n_815),
.B2(n_827),
.Y(n_910)
);

OAI22x1_ASAP7_75t_L g911 ( 
.A1(n_901),
.A2(n_800),
.B1(n_838),
.B2(n_790),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_908),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_911),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_905),
.B(n_793),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_909),
.A2(n_842),
.B(n_861),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_912),
.A2(n_907),
.B1(n_910),
.B2(n_906),
.Y(n_916)
);

NOR2x1p5_ASAP7_75t_L g917 ( 
.A(n_913),
.B(n_831),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_917),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_916),
.Y(n_919)
);

NAND2x1_ASAP7_75t_SL g920 ( 
.A(n_918),
.B(n_914),
.Y(n_920)
);

AOI21xp33_ASAP7_75t_SL g921 ( 
.A1(n_920),
.A2(n_919),
.B(n_915),
.Y(n_921)
);


endmodule