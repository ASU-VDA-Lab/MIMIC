module fake_ariane_3038_n_180 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_180);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_180;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_128;
wire n_105;
wire n_44;
wire n_82;
wire n_178;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_121;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_168;
wire n_43;
wire n_87;
wire n_81;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVxp33_ASAP7_75t_SL g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_0),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_1),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_34),
.A2(n_53),
.B1(n_51),
.B2(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_34),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_53),
.B1(n_51),
.B2(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_1),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_2),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_42),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_41),
.B1(n_32),
.B2(n_37),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_58),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_74),
.B(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_75),
.B1(n_59),
.B2(n_61),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_64),
.B(n_65),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_64),
.B(n_72),
.Y(n_96)
);

AO21x2_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_73),
.B(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_70),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_70),
.B(n_66),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_68),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_2),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_63),
.B(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_100),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_80),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_80),
.Y(n_109)
);

AOI21x1_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_82),
.B(n_86),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_87),
.B1(n_78),
.B2(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_100),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_117),
.A2(n_109),
.B(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_117),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_118),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_115),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_113),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_130),
.Y(n_141)
);

OAI21x1_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_110),
.B(n_124),
.Y(n_142)
);

AOI321xp33_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_111),
.A3(n_94),
.B1(n_131),
.B2(n_102),
.C(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NAND4xp75_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_130),
.C(n_128),
.D(n_125),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_111),
.C(n_103),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_113),
.Y(n_147)
);

OAI211xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_129),
.B(n_128),
.C(n_116),
.Y(n_148)
);

O2A1O1Ixp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_114),
.B(n_116),
.C(n_112),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_85),
.B(n_104),
.C(n_112),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_79),
.C(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_3),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_4),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_96),
.B(n_5),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_4),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_5),
.Y(n_159)
);

NAND4xp25_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_156),
.C(n_158),
.D(n_154),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_146),
.C(n_149),
.Y(n_161)
);

NOR4xp75_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_162)
);

OR3x1_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_110),
.C(n_84),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_7),
.Y(n_164)
);

NAND4xp75_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_84),
.C(n_79),
.D(n_77),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_85),
.C(n_77),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_164),
.B1(n_167),
.B2(n_166),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_8),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_83),
.B1(n_81),
.B2(n_105),
.C(n_93),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_SL g171 ( 
.A1(n_162),
.A2(n_10),
.B1(n_95),
.B2(n_83),
.C(n_81),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_81),
.Y(n_172)
);

OAI22x1_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_165),
.B1(n_105),
.B2(n_83),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_14),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_176),
.B(n_174),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_178),
.B1(n_177),
.B2(n_173),
.C(n_97),
.Y(n_180)
);


endmodule