module fake_jpeg_27377_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_31),
.Y(n_62)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_31),
.Y(n_66)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_21),
.B1(n_25),
.B2(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_55),
.B1(n_28),
.B2(n_19),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_21),
.B1(n_25),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_21),
.B1(n_25),
.B2(n_19),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_51),
.B(n_66),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_21),
.B1(n_25),
.B2(n_24),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_31),
.B1(n_16),
.B2(n_18),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_59),
.Y(n_108)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_18),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_39),
.C(n_36),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_45),
.C(n_27),
.Y(n_76)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_70),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_71),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_95),
.B1(n_101),
.B2(n_64),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_77),
.B1(n_99),
.B2(n_96),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_84),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_17),
.B1(n_20),
.B2(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_17),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_16),
.B(n_18),
.C(n_27),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_33),
.B1(n_27),
.B2(n_16),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_43),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_62),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_94),
.C(n_42),
.Y(n_126)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_17),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_33),
.B(n_20),
.C(n_35),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_30),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_19),
.B1(n_35),
.B2(n_28),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_0),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_102),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_33),
.B(n_20),
.C(n_35),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_32),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_65),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_26),
.B1(n_32),
.B2(n_23),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_50),
.B1(n_68),
.B2(n_60),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_100),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_54),
.B1(n_60),
.B2(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_28),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_34),
.B(n_26),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_11),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_56),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_119),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_134),
.B1(n_107),
.B2(n_105),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_115),
.B1(n_123),
.B2(n_135),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_54),
.B1(n_64),
.B2(n_46),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_29),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_29),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_73),
.A2(n_46),
.A3(n_42),
.B1(n_43),
.B2(n_34),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_94),
.B(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_43),
.B1(n_42),
.B2(n_26),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_34),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_126),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g128 ( 
.A1(n_73),
.A2(n_34),
.A3(n_26),
.B1(n_29),
.B2(n_23),
.Y(n_128)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_70),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_26),
.B1(n_32),
.B2(n_57),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_80),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_84),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_142),
.B(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_87),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_145),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_87),
.B1(n_76),
.B2(n_95),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_146),
.B1(n_166),
.B2(n_129),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_91),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_158),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_97),
.B(n_81),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_160),
.Y(n_182)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_169),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_102),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_157),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_72),
.Y(n_157)
);

NAND2x1p5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_94),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_101),
.B1(n_83),
.B2(n_88),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_165),
.B1(n_167),
.B2(n_120),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_106),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_71),
.B(n_100),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_163),
.B(n_170),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_75),
.B(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_164),
.B(n_168),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_114),
.A2(n_79),
.B1(n_92),
.B2(n_75),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_79),
.B1(n_78),
.B2(n_82),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_114),
.A2(n_78),
.B1(n_82),
.B2(n_85),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_115),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_180),
.B(n_185),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_172),
.B(n_175),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_181),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_179),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_109),
.C(n_127),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_168),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_125),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_192),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_161),
.B1(n_57),
.B2(n_32),
.Y(n_221)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_146),
.Y(n_191)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_109),
.Y(n_192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_129),
.B(n_128),
.C(n_135),
.D(n_127),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_148),
.B(n_152),
.C(n_130),
.D(n_137),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_23),
.B(n_1),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_141),
.B(n_129),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_142),
.Y(n_212)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_200),
.B1(n_130),
.B2(n_119),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_163),
.B1(n_147),
.B2(n_155),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_150),
.B(n_137),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_147),
.A3(n_140),
.B1(n_153),
.B2(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_221),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_143),
.B1(n_151),
.B2(n_155),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_213),
.B1(n_223),
.B2(n_227),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_214),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_143),
.B1(n_135),
.B2(n_152),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_145),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_198),
.C(n_194),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_86),
.B1(n_23),
.B2(n_14),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_225),
.B(n_1),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_0),
.B(n_1),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_197),
.B1(n_177),
.B2(n_180),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_171),
.A2(n_86),
.B1(n_23),
.B2(n_13),
.Y(n_229)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_232),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_207),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_212),
.C(n_214),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_241),
.C(n_246),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_236),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_245),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_192),
.C(n_196),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_198),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_244),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_210),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_178),
.C(n_176),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_182),
.B1(n_208),
.B2(n_190),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_178),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_254),
.B(n_255),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_205),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_250),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_233),
.A2(n_216),
.B1(n_227),
.B2(n_217),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_270),
.B1(n_243),
.B2(n_244),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_213),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_266),
.C(n_267),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_223),
.B1(n_221),
.B2(n_229),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_239),
.B1(n_231),
.B2(n_247),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_219),
.C(n_176),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_219),
.C(n_176),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_233),
.B(n_215),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_269),
.C(n_225),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_188),
.C(n_183),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_231),
.A2(n_216),
.B1(n_206),
.B2(n_224),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_247),
.B(n_259),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_285),
.B(n_184),
.Y(n_296)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_279),
.C(n_283),
.Y(n_290)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_243),
.B(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_249),
.C(n_237),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_282),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_228),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_236),
.B(n_184),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_264),
.B(n_257),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_288),
.B1(n_295),
.B2(n_275),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_267),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_294),
.B(n_281),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_255),
.B(n_254),
.Y(n_294)
);

OAI22x1_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_261),
.B1(n_268),
.B2(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_295),
.A2(n_279),
.B1(n_276),
.B2(n_273),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_300),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_288),
.A3(n_286),
.B1(n_297),
.B2(n_287),
.C1(n_6),
.C2(n_7),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_271),
.C(n_252),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_304),
.B(n_2),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_291),
.A2(n_271),
.B(n_252),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_303),
.B(n_305),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_281),
.C(n_23),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_13),
.B(n_12),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_86),
.C(n_11),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_307),
.A2(n_309),
.B1(n_311),
.B2(n_8),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_312),
.B(n_8),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_300),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_309),
.B(n_310),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_8),
.C(n_9),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_317),
.B(n_8),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_9),
.B(n_315),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_9),
.Y(n_321)
);


endmodule