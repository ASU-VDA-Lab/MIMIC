module fake_jpeg_20768_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_25),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_45),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_20),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_30),
.B1(n_18),
.B2(n_24),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_52),
.B1(n_61),
.B2(n_75),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_24),
.B1(n_28),
.B2(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_63),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_42),
.C(n_44),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_34),
.A2(n_24),
.B1(n_28),
.B2(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_18),
.B1(n_32),
.B2(n_25),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_72),
.B1(n_73),
.B2(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_36),
.A2(n_18),
.B1(n_21),
.B2(n_19),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_29),
.B1(n_21),
.B2(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_74),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_29),
.B1(n_16),
.B2(n_17),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_82),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_55),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_89),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_44),
.B1(n_16),
.B2(n_20),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_98),
.B1(n_83),
.B2(n_99),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_0),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_69),
.B1(n_64),
.B2(n_60),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_1),
.C(n_2),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_101),
.C(n_91),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_103),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_3),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_59),
.B1(n_49),
.B2(n_8),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_5),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_54),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_54),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_6),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_69),
.B(n_57),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_111),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_85),
.B1(n_8),
.B2(n_9),
.Y(n_153)
);

NOR2x1_ASAP7_75t_R g117 ( 
.A(n_99),
.B(n_74),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_88),
.B(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_128),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_125),
.B1(n_130),
.B2(n_79),
.Y(n_148)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_64),
.B1(n_71),
.B2(n_60),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_131),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_84),
.A2(n_59),
.B1(n_49),
.B2(n_9),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_13),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_152),
.C(n_117),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_80),
.C(n_78),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_141),
.C(n_144),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_140),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_78),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_147),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_87),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_106),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_104),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_123),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_87),
.B1(n_85),
.B2(n_89),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_115),
.B1(n_107),
.B2(n_126),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_85),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_7),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_10),
.Y(n_185)
);

AOI221xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_124),
.B1(n_118),
.B2(n_105),
.C(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_172),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_165),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_120),
.C(n_112),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_141),
.C(n_144),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_129),
.B(n_110),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_168),
.B(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_15),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_122),
.B(n_108),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_109),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_170),
.A2(n_148),
.B1(n_151),
.B2(n_138),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_161),
.B1(n_159),
.B2(n_155),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_181),
.C(n_158),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_185),
.B(n_163),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_135),
.C(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_181),
.C(n_176),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_179),
.A2(n_157),
.B1(n_162),
.B2(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_161),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_169),
.B1(n_168),
.B2(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_166),
.B1(n_167),
.B2(n_109),
.Y(n_196)
);

OAI22x1_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_180),
.B1(n_173),
.B2(n_178),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_185),
.B(n_174),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_206),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_204),
.A2(n_205),
.B1(n_191),
.B2(n_193),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_197),
.A2(n_175),
.B1(n_186),
.B2(n_185),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_182),
.C(n_13),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_208),
.B1(n_205),
.B2(n_202),
.Y(n_214)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_210),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_192),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_212),
.A2(n_201),
.B(n_198),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_213),
.A2(n_210),
.B(n_209),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_199),
.B(n_188),
.Y(n_218)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_215),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_217),
.B(n_218),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_216),
.C(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.C(n_10),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_14),
.Y(n_223)
);


endmodule