module fake_jpeg_24431_n_179 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_24),
.B1(n_18),
.B2(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g33 ( 
.A(n_23),
.B(n_0),
.CON(n_33),
.SN(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_46),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_42),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_21),
.Y(n_42)
);

CKINVDCx12_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_17),
.C(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_53),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_57),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_65),
.Y(n_82)
);

OA21x2_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_27),
.B(n_35),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_66),
.B1(n_44),
.B2(n_40),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_35),
.B(n_30),
.C(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_70),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_66),
.B(n_52),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_42),
.B1(n_40),
.B2(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_42),
.B1(n_26),
.B2(n_36),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_76),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_26),
.B1(n_43),
.B2(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_66),
.B1(n_54),
.B2(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_66),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_65),
.B(n_83),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_85),
.B(n_35),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_90),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_93),
.B(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_97),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_30),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_94),
.A2(n_79),
.B1(n_73),
.B2(n_71),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_94),
.B1(n_91),
.B2(n_85),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_72),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_112),
.Y(n_121)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_108),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_115),
.B(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_63),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_64),
.C(n_43),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_122),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_107),
.B(n_112),
.Y(n_134)
);

OAI322xp33_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_91),
.A3(n_93),
.B1(n_22),
.B2(n_14),
.C1(n_64),
.C2(n_20),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_20),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_127),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_69),
.B1(n_18),
.B2(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_101),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_134),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_100),
.B1(n_117),
.B2(n_128),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_124),
.B1(n_120),
.B2(n_125),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_135),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_105),
.C(n_113),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_130),
.C(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_121),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_142),
.B(n_149),
.Y(n_152)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_136),
.C(n_118),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_138),
.B1(n_103),
.B2(n_106),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_157),
.B1(n_34),
.B2(n_19),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_133),
.B1(n_15),
.B2(n_13),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_13),
.C(n_34),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_1),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_7),
.Y(n_159)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_165),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_152),
.A2(n_147),
.A3(n_19),
.B1(n_11),
.B2(n_12),
.C1(n_34),
.C2(n_4),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_153),
.C(n_155),
.Y(n_167)
);

AO21x2_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_147),
.B(n_3),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_19),
.B(n_3),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_12),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_164),
.B1(n_163),
.B2(n_162),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_2),
.C(n_4),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_168),
.B1(n_5),
.B2(n_6),
.C(n_2),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.C(n_174),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_6),
.C(n_23),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_6),
.C(n_23),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_174),
.C(n_23),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_176),
.Y(n_179)
);


endmodule