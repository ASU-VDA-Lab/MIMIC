module fake_jpeg_19401_n_187 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_15),
.B(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_39),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_33),
.B1(n_30),
.B2(n_22),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_44),
.B1(n_47),
.B2(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_12),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_24),
.B1(n_15),
.B2(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_13),
.B1(n_14),
.B2(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_20),
.B1(n_23),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_57),
.B1(n_50),
.B2(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_56),
.B1(n_34),
.B2(n_43),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_61),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_15),
.B1(n_24),
.B2(n_16),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_25),
.B1(n_27),
.B2(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_13),
.Y(n_61)
);

FAx1_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_21),
.CI(n_20),
.CON(n_62),
.SN(n_62)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_13),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

FAx1_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_38),
.CI(n_36),
.CON(n_69),
.SN(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_45),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_37),
.B1(n_21),
.B2(n_25),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_54),
.C(n_59),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_14),
.C(n_27),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_56),
.B1(n_27),
.B2(n_25),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_51),
.B1(n_43),
.B2(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_87),
.B1(n_93),
.B2(n_80),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_78),
.B1(n_93),
.B2(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_34),
.B1(n_45),
.B2(n_61),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_90),
.B1(n_73),
.B2(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_58),
.B1(n_52),
.B2(n_34),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_14),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_80),
.B1(n_77),
.B2(n_79),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_97),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_64),
.C(n_21),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_75),
.B(n_70),
.Y(n_100)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_101),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_76),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_110),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_109),
.B1(n_89),
.B2(n_95),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_107),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_69),
.B1(n_67),
.B2(n_75),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_114),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_71),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_74),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_69),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_95),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_84),
.C(n_90),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_21),
.B1(n_18),
.B2(n_7),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_107),
.B1(n_6),
.B2(n_8),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_112),
.C(n_85),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_100),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_128),
.C(n_129),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_85),
.B1(n_94),
.B2(n_86),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_94),
.B1(n_97),
.B2(n_7),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_18),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_18),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_97),
.C(n_6),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_113),
.C(n_114),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_141),
.C(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_103),
.B1(n_101),
.B2(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_143),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_117),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_5),
.C(n_10),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_143)
);

XNOR2x2_ASAP7_75t_SL g144 ( 
.A(n_142),
.B(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_134),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_139),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_143),
.Y(n_162)
);

OA21x2_ASAP7_75t_SL g146 ( 
.A1(n_134),
.A2(n_125),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_131),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_129),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_152),
.A2(n_140),
.B1(n_127),
.B2(n_147),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_141),
.B(n_148),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_158),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_160),
.Y(n_165)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_149),
.C(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_156),
.B1(n_5),
.B2(n_8),
.C(n_11),
.Y(n_171)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_173),
.B(n_1),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_11),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_0),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_175),
.B(n_0),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_11),
.B(n_9),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_5),
.B(n_1),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_177),
.A2(n_171),
.B(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_0),
.C(n_2),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_3),
.B(n_4),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_3),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_184),
.Y(n_187)
);


endmodule