module real_jpeg_13334_n_7 (n_5, n_4, n_0, n_1, n_26, n_2, n_27, n_25, n_6, n_3, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_26;
input n_2;
input n_27;
input n_25;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_23;
wire n_11;
wire n_14;
wire n_22;
wire n_18;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

NAND3xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_4),
.C(n_10),
.Y(n_9)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_0),
.A2(n_4),
.B(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_2),
.A2(n_10),
.B(n_25),
.Y(n_15)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_10),
.C(n_27),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_21),
.B(n_22),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_21),
.C(n_22),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_13),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_11),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_20),
.B(n_23),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_16),
.B(n_19),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_26),
.Y(n_18)
);


endmodule