module real_aes_8823_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g161 ( .A1(n_0), .A2(n_162), .B(n_163), .C(n_167), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_1), .B(n_156), .Y(n_169) );
INVx1_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_3), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_4), .A2(n_150), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_5), .A2(n_130), .B(n_147), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_6), .A2(n_150), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_7), .B(n_156), .Y(n_475) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_8), .A2(n_122), .B(n_244), .Y(n_243) );
AND2x6_ASAP7_75t_L g147 ( .A(n_9), .B(n_148), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_10), .A2(n_130), .B(n_147), .C(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g566 ( .A(n_11), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_12), .B(n_39), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_13), .B(n_166), .Y(n_515) );
INVx1_ASAP7_75t_L g127 ( .A(n_14), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_15), .B(n_141), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_16), .A2(n_142), .B(n_524), .C(n_526), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_17), .B(n_156), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_18), .B(n_184), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_19), .A2(n_130), .B(n_176), .C(n_183), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_20), .A2(n_165), .B(n_218), .C(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_21), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_22), .B(n_166), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_23), .B(n_166), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_24), .Y(n_493) );
INVx1_ASAP7_75t_L g463 ( .A(n_25), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_26), .A2(n_130), .B(n_183), .C(n_247), .Y(n_246) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_27), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_28), .Y(n_511) );
INVx1_ASAP7_75t_L g487 ( .A(n_29), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_30), .A2(n_150), .B(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g132 ( .A(n_31), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_32), .A2(n_145), .B(n_199), .C(n_200), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_33), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_34), .A2(n_165), .B(n_472), .C(n_474), .Y(n_471) );
INVxp67_ASAP7_75t_L g488 ( .A(n_35), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_36), .B(n_249), .Y(n_248) );
CKINVDCx14_ASAP7_75t_R g470 ( .A(n_37), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_38), .A2(n_130), .B(n_183), .C(n_462), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_40), .A2(n_167), .B(n_564), .C(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_41), .B(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_42), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_43), .B(n_141), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_44), .B(n_150), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_45), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_46), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_47), .A2(n_145), .B(n_199), .C(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g164 ( .A(n_48), .Y(n_164) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_49), .A2(n_103), .B1(n_430), .B2(n_437), .C1(n_721), .C2(n_726), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g110 ( .A1(n_49), .A2(n_111), .B1(n_425), .B2(n_426), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_49), .Y(n_425) );
INVx1_ASAP7_75t_L g228 ( .A(n_50), .Y(n_228) );
INVx1_ASAP7_75t_L g531 ( .A(n_51), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_52), .B(n_150), .Y(n_225) );
OAI22xp5_ASAP7_75t_SL g112 ( .A1(n_53), .A2(n_71), .B1(n_113), .B2(n_114), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_53), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_54), .Y(n_188) );
AOI222xp33_ASAP7_75t_SL g438 ( .A1(n_55), .A2(n_439), .B1(n_445), .B2(n_715), .C1(n_716), .C2(n_717), .Y(n_438) );
CKINVDCx14_ASAP7_75t_R g562 ( .A(n_56), .Y(n_562) );
INVx1_ASAP7_75t_L g148 ( .A(n_57), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_58), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_59), .B(n_156), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_60), .A2(n_137), .B(n_182), .C(n_239), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_61), .A2(n_70), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_61), .Y(n_443) );
INVx1_ASAP7_75t_L g126 ( .A(n_62), .Y(n_126) );
INVx1_ASAP7_75t_SL g473 ( .A(n_63), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_64), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_65), .B(n_141), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_66), .B(n_156), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_67), .B(n_142), .Y(n_215) );
INVx1_ASAP7_75t_L g496 ( .A(n_68), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g159 ( .A(n_69), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_70), .Y(n_444) );
INVx1_ASAP7_75t_L g114 ( .A(n_71), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_72), .B(n_178), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_73), .A2(n_130), .B(n_135), .C(n_145), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_74), .Y(n_237) );
INVx1_ASAP7_75t_L g436 ( .A(n_75), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_76), .A2(n_150), .B(n_561), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_77), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_78), .A2(n_150), .B(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_79), .A2(n_174), .B(n_483), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_80), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_81), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_81), .Y(n_440) );
INVx1_ASAP7_75t_L g522 ( .A(n_82), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_83), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_84), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_85), .A2(n_150), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g525 ( .A(n_86), .Y(n_525) );
INVx2_ASAP7_75t_L g124 ( .A(n_87), .Y(n_124) );
INVx1_ASAP7_75t_L g514 ( .A(n_88), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_89), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_90), .B(n_166), .Y(n_216) );
OR2x2_ASAP7_75t_L g105 ( .A(n_91), .B(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g449 ( .A(n_91), .B(n_107), .Y(n_449) );
INVx2_ASAP7_75t_L g714 ( .A(n_91), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_92), .A2(n_130), .B(n_145), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_93), .B(n_150), .Y(n_197) );
INVx1_ASAP7_75t_L g201 ( .A(n_94), .Y(n_201) );
INVxp67_ASAP7_75t_L g240 ( .A(n_95), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_96), .B(n_122), .Y(n_567) );
INVx1_ASAP7_75t_L g136 ( .A(n_97), .Y(n_136) );
INVx1_ASAP7_75t_L g211 ( .A(n_98), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_99), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g534 ( .A(n_100), .Y(n_534) );
AND2x2_ASAP7_75t_L g230 ( .A(n_101), .B(n_186), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_110), .B(n_427), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_105), .Y(n_429) );
INVx1_ASAP7_75t_SL g725 ( .A(n_105), .Y(n_725) );
BUFx2_ASAP7_75t_L g728 ( .A(n_105), .Y(n_728) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_106), .B(n_714), .Y(n_715) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g713 ( .A(n_107), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g426 ( .A(n_111), .Y(n_426) );
XNOR2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_115), .Y(n_111) );
INVx1_ASAP7_75t_L g446 ( .A(n_115), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_115), .A2(n_451), .B1(n_718), .B2(n_719), .Y(n_717) );
OR3x1_ASAP7_75t_L g115 ( .A(n_116), .B(n_333), .C(n_382), .Y(n_115) );
NAND5xp2_ASAP7_75t_L g116 ( .A(n_117), .B(n_267), .C(n_296), .D(n_304), .E(n_319), .Y(n_116) );
O2A1O1Ixp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_190), .B(n_206), .C(n_251), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_170), .Y(n_118) );
AND2x2_ASAP7_75t_L g262 ( .A(n_119), .B(n_259), .Y(n_262) );
AND2x2_ASAP7_75t_L g295 ( .A(n_119), .B(n_171), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_119), .B(n_194), .Y(n_388) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_155), .Y(n_119) );
INVx2_ASAP7_75t_L g193 ( .A(n_120), .Y(n_193) );
BUFx2_ASAP7_75t_L g362 ( .A(n_120), .Y(n_362) );
AO21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_128), .B(n_153), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_121), .B(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g156 ( .A(n_121), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_121), .B(n_205), .Y(n_204) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_121), .A2(n_210), .B(n_220), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_121), .B(n_466), .Y(n_465) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_121), .A2(n_492), .B(n_499), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_121), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_122), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_122), .A2(n_245), .B(n_246), .Y(n_244) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g222 ( .A(n_123), .Y(n_222) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x2_ASAP7_75t_SL g186 ( .A(n_124), .B(n_125), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_149), .Y(n_128) );
INVx5_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
BUFx3_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g152 ( .A(n_132), .Y(n_152) );
INVx1_ASAP7_75t_L g219 ( .A(n_132), .Y(n_219) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_134), .Y(n_139) );
INVx3_ASAP7_75t_L g142 ( .A(n_134), .Y(n_142) );
AND2x2_ASAP7_75t_L g151 ( .A(n_134), .B(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_134), .Y(n_166) );
INVx1_ASAP7_75t_L g249 ( .A(n_134), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_140), .C(n_143), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_138), .A2(n_141), .B1(n_487), .B2(n_488), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_138), .B(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_138), .B(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
INVx2_ASAP7_75t_L g162 ( .A(n_141), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_141), .B(n_240), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_141), .A2(n_181), .B(n_463), .C(n_464), .Y(n_462) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_142), .B(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g474 ( .A(n_144), .Y(n_474) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_SL g158 ( .A1(n_146), .A2(n_159), .B(n_160), .C(n_161), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_146), .A2(n_160), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_146), .A2(n_160), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_146), .A2(n_160), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_146), .A2(n_160), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_146), .A2(n_160), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_SL g561 ( .A1(n_146), .A2(n_160), .B(n_562), .C(n_563), .Y(n_561) );
INVx4_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g150 ( .A(n_147), .B(n_151), .Y(n_150) );
BUFx3_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g212 ( .A(n_147), .B(n_151), .Y(n_212) );
BUFx2_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
INVx1_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
AND2x2_ASAP7_75t_L g170 ( .A(n_155), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g260 ( .A(n_155), .Y(n_260) );
AND2x2_ASAP7_75t_L g346 ( .A(n_155), .B(n_259), .Y(n_346) );
AND2x2_ASAP7_75t_L g401 ( .A(n_155), .B(n_193), .Y(n_401) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_169), .Y(n_155) );
INVx2_ASAP7_75t_L g199 ( .A(n_160), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_165), .B(n_473), .Y(n_472) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g564 ( .A(n_166), .Y(n_564) );
INVx2_ASAP7_75t_L g498 ( .A(n_167), .Y(n_498) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_168), .Y(n_203) );
INVx1_ASAP7_75t_L g526 ( .A(n_168), .Y(n_526) );
INVx1_ASAP7_75t_L g318 ( .A(n_170), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_170), .B(n_194), .Y(n_365) );
INVx5_ASAP7_75t_L g259 ( .A(n_171), .Y(n_259) );
AND2x4_ASAP7_75t_L g280 ( .A(n_171), .B(n_260), .Y(n_280) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_171), .Y(n_302) );
AND2x2_ASAP7_75t_L g377 ( .A(n_171), .B(n_362), .Y(n_377) );
AND2x2_ASAP7_75t_L g380 ( .A(n_171), .B(n_195), .Y(n_380) );
OR2x6_ASAP7_75t_L g171 ( .A(n_172), .B(n_187), .Y(n_171) );
AOI21xp5_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_175), .B(n_184), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B(n_181), .Y(n_176) );
INVx2_ASAP7_75t_L g180 ( .A(n_178), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_180), .A2(n_201), .B(n_202), .C(n_203), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_180), .A2(n_203), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_180), .A2(n_496), .B(n_497), .C(n_498), .Y(n_495) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_180), .A2(n_498), .B(n_514), .C(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_182), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_185), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g189 ( .A(n_186), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_186), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_186), .A2(n_225), .B(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_186), .A2(n_212), .B(n_460), .C(n_461), .Y(n_459) );
OA21x2_ASAP7_75t_L g559 ( .A1(n_186), .A2(n_560), .B(n_567), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_189), .A2(n_510), .B(n_516), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_190), .B(n_260), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_190), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_194), .Y(n_191) );
AND2x2_ASAP7_75t_L g285 ( .A(n_192), .B(n_260), .Y(n_285) );
AND2x2_ASAP7_75t_L g303 ( .A(n_192), .B(n_195), .Y(n_303) );
INVx1_ASAP7_75t_L g323 ( .A(n_192), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_192), .B(n_259), .Y(n_368) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_192), .Y(n_410) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_193), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_194), .B(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_194), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_194), .A2(n_255), .B(n_316), .C(n_318), .Y(n_315) );
AND2x2_ASAP7_75t_L g322 ( .A(n_194), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g331 ( .A(n_194), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g335 ( .A(n_194), .B(n_259), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_194), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g350 ( .A(n_194), .B(n_260), .Y(n_350) );
AND2x2_ASAP7_75t_L g400 ( .A(n_194), .B(n_401), .Y(n_400) );
INVx5_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
BUFx2_ASAP7_75t_L g264 ( .A(n_195), .Y(n_264) );
AND2x2_ASAP7_75t_L g305 ( .A(n_195), .B(n_258), .Y(n_305) );
AND2x2_ASAP7_75t_L g317 ( .A(n_195), .B(n_292), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_195), .B(n_346), .Y(n_364) );
OR2x6_ASAP7_75t_L g195 ( .A(n_196), .B(n_204), .Y(n_195) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_231), .Y(n_206) );
INVx1_ASAP7_75t_L g253 ( .A(n_207), .Y(n_253) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_223), .Y(n_207) );
OR2x2_ASAP7_75t_L g255 ( .A(n_208), .B(n_223), .Y(n_255) );
NAND3xp33_ASAP7_75t_L g261 ( .A(n_208), .B(n_262), .C(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_208), .B(n_233), .Y(n_272) );
OR2x2_ASAP7_75t_L g287 ( .A(n_208), .B(n_275), .Y(n_287) );
AND2x2_ASAP7_75t_L g293 ( .A(n_208), .B(n_242), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_208), .B(n_424), .Y(n_423) );
INVx5_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_209), .B(n_233), .Y(n_290) );
AND2x2_ASAP7_75t_L g329 ( .A(n_209), .B(n_243), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_209), .B(n_242), .Y(n_357) );
OR2x2_ASAP7_75t_L g360 ( .A(n_209), .B(n_242), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_212), .A2(n_493), .B(n_494), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_212), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_217), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_217), .A2(n_248), .B(n_250), .Y(n_247) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g481 ( .A(n_222), .Y(n_481) );
INVx5_ASAP7_75t_SL g275 ( .A(n_223), .Y(n_275) );
OR2x2_ASAP7_75t_L g281 ( .A(n_223), .B(n_232), .Y(n_281) );
AND2x2_ASAP7_75t_L g297 ( .A(n_223), .B(n_298), .Y(n_297) );
AOI321xp33_ASAP7_75t_L g304 ( .A1(n_223), .A2(n_305), .A3(n_306), .B1(n_307), .B2(n_313), .C(n_315), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_223), .B(n_231), .Y(n_314) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_223), .Y(n_327) );
OR2x2_ASAP7_75t_L g374 ( .A(n_223), .B(n_272), .Y(n_374) );
AND2x2_ASAP7_75t_L g396 ( .A(n_223), .B(n_293), .Y(n_396) );
AND2x2_ASAP7_75t_L g415 ( .A(n_223), .B(n_233), .Y(n_415) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_230), .Y(n_223) );
INVx1_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_242), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_233), .B(n_242), .Y(n_256) );
AND2x2_ASAP7_75t_L g265 ( .A(n_233), .B(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g292 ( .A(n_233), .Y(n_292) );
AND2x2_ASAP7_75t_L g298 ( .A(n_233), .B(n_293), .Y(n_298) );
INVxp67_ASAP7_75t_L g328 ( .A(n_233), .Y(n_328) );
OR2x2_ASAP7_75t_L g370 ( .A(n_233), .B(n_275), .Y(n_370) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_241), .Y(n_233) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_234), .A2(n_468), .B(n_475), .Y(n_467) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_234), .A2(n_520), .B(n_527), .Y(n_519) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_234), .A2(n_529), .B(n_535), .Y(n_528) );
OR2x2_ASAP7_75t_L g252 ( .A(n_242), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_SL g266 ( .A(n_242), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_242), .B(n_255), .Y(n_299) );
AND2x2_ASAP7_75t_L g348 ( .A(n_242), .B(n_292), .Y(n_348) );
AND2x2_ASAP7_75t_L g386 ( .A(n_242), .B(n_275), .Y(n_386) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_243), .B(n_275), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_254), .B(n_257), .C(n_261), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_252), .A2(n_254), .B1(n_379), .B2(n_381), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_254), .A2(n_277), .B1(n_332), .B2(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_SL g406 ( .A(n_255), .Y(n_406) );
INVx1_ASAP7_75t_SL g306 ( .A(n_256), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_258), .B(n_278), .Y(n_308) );
AOI222xp33_ASAP7_75t_L g319 ( .A1(n_258), .A2(n_299), .B1(n_306), .B2(n_320), .C1(n_324), .C2(n_330), .Y(n_319) );
AND2x2_ASAP7_75t_L g409 ( .A(n_258), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_259), .B(n_279), .Y(n_354) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_259), .Y(n_391) );
AND2x2_ASAP7_75t_L g394 ( .A(n_259), .B(n_303), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_259), .B(n_410), .Y(n_420) );
INVx1_ASAP7_75t_L g311 ( .A(n_260), .Y(n_311) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_260), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_262), .A2(n_403), .B(n_404), .C(n_407), .Y(n_402) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_264), .B(n_326), .C(n_329), .Y(n_325) );
OR2x2_ASAP7_75t_L g353 ( .A(n_264), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_264), .B(n_280), .Y(n_381) );
OR2x2_ASAP7_75t_L g286 ( .A(n_266), .B(n_287), .Y(n_286) );
AOI211xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_270), .B(n_276), .C(n_288), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_269), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g375 ( .A(n_270), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_271), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g289 ( .A(n_274), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_275), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g343 ( .A(n_275), .B(n_293), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_275), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_275), .B(n_292), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B1(n_282), .B2(n_286), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_278), .B(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_280), .B(n_322), .Y(n_321) );
OAI221xp5_ASAP7_75t_SL g344 ( .A1(n_281), .A2(n_345), .B1(n_347), .B2(n_349), .C(n_351), .Y(n_344) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g399 ( .A(n_284), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g412 ( .A(n_284), .B(n_401), .Y(n_412) );
INVx1_ASAP7_75t_L g332 ( .A(n_285), .Y(n_332) );
INVx1_ASAP7_75t_L g403 ( .A(n_286), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_287), .A2(n_370), .B(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B(n_294), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI21xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_299), .B(n_300), .Y(n_296) );
INVx1_ASAP7_75t_L g336 ( .A(n_297), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_298), .A2(n_384), .B1(n_387), .B2(n_389), .C(n_392), .Y(n_383) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_306), .A2(n_396), .B1(n_397), .B2(n_399), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g372 ( .A(n_308), .Y(n_372) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp67_ASAP7_75t_SL g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g376 ( .A(n_312), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g341 ( .A(n_317), .Y(n_341) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_322), .B(n_346), .Y(n_398) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_328), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g414 ( .A(n_329), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g421 ( .A(n_329), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI211xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_336), .B(n_337), .C(n_371), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI211xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B(n_344), .C(n_363), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g424 ( .A(n_348), .Y(n_424) );
AND2x2_ASAP7_75t_L g361 ( .A(n_350), .B(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B1(n_359), .B2(n_361), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OR2x2_ASAP7_75t_L g369 ( .A(n_357), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g422 ( .A(n_358), .Y(n_422) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI31xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .A3(n_366), .B(n_369), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI211xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B(n_375), .C(n_378), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g379 ( .A(n_380), .Y(n_379) );
NAND5xp2_ASAP7_75t_L g382 ( .A(n_383), .B(n_395), .C(n_402), .D(n_416), .E(n_419), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_394), .A2(n_420), .B1(n_421), .B2(n_423), .Y(n_419) );
INVx1_ASAP7_75t_SL g418 ( .A(n_396), .Y(n_418) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B(n_413), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_SL g723 ( .A(n_433), .B(n_435), .Y(n_723) );
OA21x2_ASAP7_75t_L g727 ( .A1(n_433), .A2(n_434), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g716 ( .A(n_439), .Y(n_716) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_447), .B1(n_450), .B2(n_713), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g718 ( .A(n_448), .Y(n_718) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR3x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_624), .C(n_671), .Y(n_451) );
NAND3xp33_ASAP7_75t_SL g452 ( .A(n_453), .B(n_570), .C(n_595), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_508), .B1(n_536), .B2(n_539), .C(n_547), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_476), .B(n_501), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_456), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_456), .B(n_552), .Y(n_668) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_467), .Y(n_456) );
AND2x2_ASAP7_75t_L g538 ( .A(n_457), .B(n_507), .Y(n_538) );
AND2x2_ASAP7_75t_L g588 ( .A(n_457), .B(n_506), .Y(n_588) );
AND2x2_ASAP7_75t_L g609 ( .A(n_457), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g614 ( .A(n_457), .B(n_581), .Y(n_614) );
OR2x2_ASAP7_75t_L g622 ( .A(n_457), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g694 ( .A(n_457), .B(n_490), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_457), .B(n_643), .Y(n_708) );
INVx3_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g553 ( .A(n_458), .B(n_467), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_458), .B(n_490), .Y(n_554) );
AND2x4_ASAP7_75t_L g576 ( .A(n_458), .B(n_507), .Y(n_576) );
AND2x2_ASAP7_75t_L g606 ( .A(n_458), .B(n_478), .Y(n_606) );
AND2x2_ASAP7_75t_L g615 ( .A(n_458), .B(n_605), .Y(n_615) );
AND2x2_ASAP7_75t_L g631 ( .A(n_458), .B(n_491), .Y(n_631) );
OR2x2_ASAP7_75t_L g640 ( .A(n_458), .B(n_623), .Y(n_640) );
AND2x2_ASAP7_75t_L g646 ( .A(n_458), .B(n_581), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_458), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g660 ( .A(n_458), .B(n_503), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_458), .B(n_549), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_458), .B(n_610), .Y(n_699) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_465), .Y(n_458) );
INVx2_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
AND2x2_ASAP7_75t_L g605 ( .A(n_467), .B(n_490), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_467), .B(n_491), .Y(n_610) );
INVx1_ASAP7_75t_L g666 ( .A(n_467), .Y(n_666) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g575 ( .A(n_477), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_490), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_478), .B(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
OR2x2_ASAP7_75t_L g623 ( .A(n_478), .B(n_490), .Y(n_623) );
OR2x2_ASAP7_75t_L g684 ( .A(n_478), .B(n_591), .Y(n_684) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_482), .B(n_489), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_480), .A2(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g504 ( .A(n_482), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_489), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_490), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g643 ( .A(n_490), .B(n_503), .Y(n_643) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g582 ( .A(n_491), .Y(n_582) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_502), .A2(n_688), .B1(n_692), .B2(n_695), .C(n_696), .Y(n_687) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .Y(n_502) );
INVx1_ASAP7_75t_SL g550 ( .A(n_503), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_503), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g682 ( .A(n_503), .B(n_538), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_506), .B(n_552), .Y(n_674) );
AND2x2_ASAP7_75t_L g581 ( .A(n_507), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g585 ( .A(n_508), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_508), .B(n_591), .Y(n_621) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
AND2x2_ASAP7_75t_L g546 ( .A(n_509), .B(n_519), .Y(n_546) );
INVx4_ASAP7_75t_L g558 ( .A(n_509), .Y(n_558) );
BUFx3_ASAP7_75t_L g601 ( .A(n_509), .Y(n_601) );
AND3x2_ASAP7_75t_L g616 ( .A(n_509), .B(n_617), .C(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g698 ( .A(n_518), .B(n_612), .Y(n_698) );
AND2x2_ASAP7_75t_L g706 ( .A(n_518), .B(n_591), .Y(n_706) );
INVx1_ASAP7_75t_SL g711 ( .A(n_518), .Y(n_711) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
INVx1_ASAP7_75t_SL g569 ( .A(n_519), .Y(n_569) );
AND2x2_ASAP7_75t_L g592 ( .A(n_519), .B(n_558), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_519), .B(n_542), .Y(n_594) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_519), .Y(n_634) );
OR2x2_ASAP7_75t_L g639 ( .A(n_519), .B(n_558), .Y(n_639) );
INVx2_ASAP7_75t_L g544 ( .A(n_528), .Y(n_544) );
AND2x2_ASAP7_75t_L g579 ( .A(n_528), .B(n_559), .Y(n_579) );
OR2x2_ASAP7_75t_L g599 ( .A(n_528), .B(n_559), .Y(n_599) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_528), .Y(n_619) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_537), .A2(n_578), .B(n_670), .Y(n_669) );
AOI322xp5_ASAP7_75t_L g705 ( .A1(n_539), .A2(n_549), .A3(n_576), .B1(n_706), .B2(n_707), .C1(n_709), .C2(n_712), .Y(n_705) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_541), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_542), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g568 ( .A(n_543), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g636 ( .A(n_544), .B(n_558), .Y(n_636) );
AND2x2_ASAP7_75t_L g703 ( .A(n_544), .B(n_559), .Y(n_703) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g644 ( .A(n_546), .B(n_598), .Y(n_644) );
AOI31xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_551), .A3(n_554), .B(n_555), .Y(n_547) );
AND2x2_ASAP7_75t_L g603 ( .A(n_549), .B(n_581), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_549), .B(n_573), .Y(n_685) );
AND2x2_ASAP7_75t_L g704 ( .A(n_549), .B(n_609), .Y(n_704) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_552), .B(n_581), .Y(n_593) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_552), .B(n_610), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_552), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_552), .B(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_553), .B(n_610), .Y(n_642) );
INVx1_ASAP7_75t_L g686 ( .A(n_553), .Y(n_686) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_568), .Y(n_556) );
INVxp67_ASAP7_75t_L g638 ( .A(n_557), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_558), .B(n_569), .Y(n_574) );
INVx1_ASAP7_75t_L g680 ( .A(n_558), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_558), .B(n_657), .Y(n_691) );
BUFx3_ASAP7_75t_L g591 ( .A(n_559), .Y(n_591) );
AND2x2_ASAP7_75t_L g617 ( .A(n_559), .B(n_569), .Y(n_617) );
INVx2_ASAP7_75t_L g657 ( .A(n_559), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_568), .B(n_690), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_575), .B(n_577), .C(n_586), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_572), .A2(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_573), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_573), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g653 ( .A(n_574), .B(n_599), .Y(n_653) );
INVx3_ASAP7_75t_L g584 ( .A(n_576), .Y(n_584) );
OAI22xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_580), .B1(n_583), .B2(n_585), .Y(n_577) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_579), .A2(n_603), .B(n_604), .Y(n_602) );
AND2x2_ASAP7_75t_L g628 ( .A(n_579), .B(n_592), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_579), .B(n_680), .Y(n_679) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g583 ( .A(n_582), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g652 ( .A(n_582), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_583), .A2(n_597), .B(n_602), .Y(n_596) );
OAI22xp33_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_589), .B1(n_593), .B2(n_594), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_588), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g612 ( .A(n_591), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_591), .B(n_634), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_607), .C(n_620), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g662 ( .A1(n_597), .A2(n_663), .B1(n_667), .B2(n_668), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g667 ( .A(n_599), .B(n_600), .Y(n_667) );
AND2x2_ASAP7_75t_L g675 ( .A(n_600), .B(n_656), .Y(n_675) );
CKINVDCx16_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_SL g683 ( .A1(n_601), .A2(n_684), .B(n_685), .C(n_686), .Y(n_683) );
OR2x2_ASAP7_75t_L g710 ( .A(n_601), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_611), .B(n_613), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_609), .A2(n_646), .B(n_647), .C(n_650), .Y(n_645) );
OAI21xp33_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_615), .B(n_616), .Y(n_613) );
AND2x2_ASAP7_75t_L g678 ( .A(n_617), .B(n_636), .Y(n_678) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g656 ( .A(n_619), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_621), .Y(n_661) );
NAND3xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_645), .C(n_658), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B(n_629), .C(n_637), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g695 ( .A(n_632), .Y(n_695) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_634), .B(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_640), .C(n_641), .Y(n_637) );
INVx2_ASAP7_75t_SL g649 ( .A(n_639), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_640), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_650) );
OAI21xp33_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_643), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_661), .B(n_662), .C(n_669), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVxp33_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g712 ( .A(n_666), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_672), .B(n_687), .C(n_700), .D(n_705), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B(n_676), .C(n_683), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B(n_681), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g696 ( .A1(n_677), .A2(n_697), .B(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_684), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_704), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g720 ( .A(n_713), .Y(n_720) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
NAND2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
endmodule