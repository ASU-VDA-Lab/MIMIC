module fake_jpeg_28232_n_205 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_12),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_29),
.B1(n_30),
.B2(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_53),
.Y(n_63)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_30),
.B1(n_24),
.B2(n_13),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_51),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_26),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_36),
.C(n_25),
.Y(n_68)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_29),
.B1(n_30),
.B2(n_13),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_31),
.B1(n_12),
.B2(n_28),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_26),
.B(n_25),
.C(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_25),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_84),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_49),
.B(n_43),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_54),
.B1(n_51),
.B2(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

XNOR2x1_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_54),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_62),
.B1(n_72),
.B2(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_53),
.B1(n_57),
.B2(n_50),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_62),
.B1(n_86),
.B2(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_32),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_97),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_99),
.B1(n_44),
.B2(n_58),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_62),
.B1(n_67),
.B2(n_65),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_88),
.B1(n_77),
.B2(n_75),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_62),
.B1(n_57),
.B2(n_50),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_69),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_108),
.B1(n_112),
.B2(n_114),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_76),
.B1(n_79),
.B2(n_83),
.C(n_80),
.Y(n_106)
);

OAI322xp33_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_21),
.A3(n_19),
.B1(n_14),
.B2(n_17),
.C1(n_23),
.C2(n_22),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_76),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_71),
.C(n_25),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_112),
.C(n_114),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_80),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_69),
.B1(n_58),
.B2(n_34),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_66),
.B(n_1),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_91),
.B(n_98),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_26),
.C(n_55),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_97),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_26),
.C(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_58),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_92),
.B(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_124),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_92),
.B(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_126),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_133),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_99),
.Y(n_128)
);

AOI31xp67_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_130),
.A3(n_21),
.B(n_19),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_28),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_58),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_15),
.B(n_17),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_131),
.B(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_142),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_69),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_15),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_23),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_122),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_22),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_146),
.C(n_150),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_23),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_149),
.B1(n_125),
.B2(n_136),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_52),
.B1(n_45),
.B2(n_48),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_23),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_122),
.C(n_127),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_161),
.C(n_163),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_19),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_14),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_133),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_123),
.B1(n_121),
.B2(n_31),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_162),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_32),
.C(n_45),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_32),
.C(n_19),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_5),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_138),
.B1(n_149),
.B2(n_9),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_167),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_8),
.B1(n_10),
.B2(n_9),
.Y(n_167)
);

AOI31xp33_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_7),
.A3(n_11),
.B(n_8),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_175),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_163),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_6),
.B(n_8),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_7),
.B(n_5),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_170),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_180),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_156),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_4),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_R g191 ( 
.A(n_183),
.B(n_4),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_156),
.B(n_7),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_184),
.A2(n_4),
.B(n_3),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_173),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_174),
.B1(n_169),
.B2(n_14),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_189),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_192),
.Y(n_195)
);

OA21x2_ASAP7_75t_SL g198 ( 
.A1(n_191),
.A2(n_0),
.B(n_21),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_3),
.B1(n_19),
.B2(n_2),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_185),
.A2(n_179),
.B(n_1),
.Y(n_194)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_0),
.B(n_38),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_198),
.A2(n_0),
.B1(n_197),
.B2(n_195),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_199),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_190),
.C(n_38),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_201),
.B(n_196),
.C(n_202),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_203),
.Y(n_205)
);


endmodule