module fake_jpeg_3673_n_170 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_25),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_66),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_63),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_89),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_66),
.B(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_53),
.B1(n_51),
.B2(n_57),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_96),
.B1(n_53),
.B2(n_60),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_88),
.Y(n_99)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_55),
.C(n_49),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_46),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_57),
.B1(n_56),
.B2(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_53),
.B1(n_52),
.B2(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_106),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_0),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_96),
.B1(n_91),
.B2(n_87),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_1),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_6),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_120),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_3),
.B(n_5),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_13),
.B(n_16),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_6),
.B(n_7),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_131),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_130),
.Y(n_133)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_11),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_12),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_110),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_13),
.B(n_15),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_110),
.C(n_102),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_146),
.C(n_116),
.Y(n_148)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_126),
.B1(n_119),
.B2(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_149),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_24),
.C(n_26),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_136),
.B1(n_133),
.B2(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_135),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_139),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_159),
.B(n_156),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_141),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_162),
.B1(n_150),
.B2(n_143),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_157),
.A2(n_139),
.B(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_160),
.A2(n_150),
.B1(n_146),
.B2(n_31),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_35),
.C(n_36),
.Y(n_167)
);

AOI221xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_44),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_43),
.Y(n_170)
);


endmodule