module fake_jpeg_2344_n_711 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_711);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_711;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_60),
.Y(n_151)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_63),
.B(n_70),
.Y(n_148)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_10),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_71),
.B(n_102),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_36),
.A2(n_9),
.B(n_17),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_72),
.A2(n_31),
.B(n_55),
.C(n_26),
.Y(n_194)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_78),
.Y(n_181)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_81),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_82),
.Y(n_212)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_84),
.Y(n_213)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_87),
.Y(n_184)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_88),
.Y(n_205)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_89),
.Y(n_186)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_92),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g221 ( 
.A(n_94),
.Y(n_221)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_97),
.Y(n_193)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_57),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_99),
.Y(n_224)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_27),
.B(n_18),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_41),
.B(n_17),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_120),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_111),
.Y(n_215)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_21),
.Y(n_112)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_113),
.Y(n_219)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_116),
.Y(n_229)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_39),
.B(n_17),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_122),
.Y(n_227)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_43),
.B(n_16),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_127),
.Y(n_179)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_41),
.B(n_16),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_131),
.Y(n_198)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_23),
.Y(n_132)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_48),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_140),
.B(n_206),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_40),
.B1(n_54),
.B2(n_25),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_141),
.A2(n_146),
.B1(n_200),
.B2(n_226),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_62),
.A2(n_40),
.B1(n_54),
.B2(n_25),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_73),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_149),
.B(n_161),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_157),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_92),
.B(n_53),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_74),
.A2(n_54),
.B1(n_45),
.B2(n_49),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_164),
.A2(n_178),
.B1(n_126),
.B2(n_122),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_90),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_172),
.B(n_177),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_99),
.B(n_53),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_65),
.A2(n_40),
.B1(n_52),
.B2(n_39),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_23),
.C(n_52),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_180),
.B(n_51),
.C(n_21),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_128),
.B(n_49),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_185),
.B(n_194),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_34),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_195),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_83),
.A2(n_44),
.B1(n_55),
.B2(n_24),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_191),
.A2(n_220),
.B1(n_20),
.B2(n_1),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_88),
.B(n_34),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_94),
.B(n_34),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_197),
.B(n_214),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_67),
.A2(n_44),
.B1(n_55),
.B2(n_24),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_115),
.B(n_44),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_112),
.B(n_31),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_208),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_80),
.B(n_31),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_117),
.A2(n_26),
.B(n_24),
.C(n_28),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_118),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_130),
.A2(n_44),
.B1(n_26),
.B2(n_58),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_82),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_84),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_91),
.Y(n_225)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_225),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_96),
.A2(n_58),
.B1(n_51),
.B2(n_28),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_103),
.Y(n_228)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_108),
.B(n_58),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_2),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_164),
.A2(n_28),
.B(n_51),
.C(n_21),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g349 ( 
.A1(n_232),
.A2(n_271),
.B(n_273),
.Y(n_349)
);

INVx11_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_233),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_234),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_235),
.B(n_288),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_236),
.A2(n_254),
.B1(n_301),
.B2(n_171),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_139),
.A2(n_116),
.B1(n_110),
.B2(n_109),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_237),
.A2(n_265),
.B1(n_297),
.B2(n_298),
.Y(n_322)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

INVx4_ASAP7_75t_SL g326 ( 
.A(n_240),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_68),
.B1(n_20),
.B2(n_16),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_241),
.A2(n_291),
.B1(n_190),
.B2(n_174),
.Y(n_328)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g341 ( 
.A(n_244),
.Y(n_341)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g372 ( 
.A(n_246),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_133),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_250),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_179),
.A2(n_20),
.B1(n_15),
.B2(n_14),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_251),
.A2(n_269),
.B1(n_284),
.B2(n_150),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_140),
.A2(n_209),
.B1(n_168),
.B2(n_148),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_253),
.A2(n_278),
.B1(n_248),
.B2(n_259),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_168),
.A2(n_20),
.B1(n_15),
.B2(n_14),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_133),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_255),
.Y(n_366)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_187),
.Y(n_256)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

INVx3_ASAP7_75t_SL g257 ( 
.A(n_151),
.Y(n_257)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_258),
.B(n_267),
.C(n_275),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_179),
.A2(n_20),
.B1(n_14),
.B2(n_13),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_260),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_189),
.B(n_0),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_274),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_136),
.Y(n_262)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_262),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_143),
.B(n_14),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_266),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_224),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_138),
.Y(n_268)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_268),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_148),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_269)
);

AO22x1_ASAP7_75t_SL g270 ( 
.A1(n_206),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_270)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_134),
.B(n_0),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_197),
.B(n_2),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_157),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_192),
.B(n_4),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_285),
.Y(n_330)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_153),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_289),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_226),
.A2(n_11),
.B1(n_12),
.B2(n_7),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_137),
.B(n_5),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_165),
.Y(n_286)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_217),
.Y(n_287)
);

BUFx24_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g288 ( 
.A1(n_220),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_167),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_144),
.Y(n_290)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_290),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_227),
.A2(n_12),
.B1(n_6),
.B2(n_8),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_183),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_293),
.Y(n_335)
);

INVx4_ASAP7_75t_SL g293 ( 
.A(n_218),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_294),
.Y(n_359)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_136),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_295),
.Y(n_327)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_162),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_299),
.Y(n_340)
);

INVx11_ASAP7_75t_L g297 ( 
.A(n_166),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_160),
.A2(n_12),
.B1(n_6),
.B2(n_8),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_181),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_191),
.A2(n_5),
.B(n_8),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_159),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_L g301 ( 
.A1(n_170),
.A2(n_5),
.B1(n_8),
.B2(n_230),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_202),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_302),
.B(n_303),
.Y(n_357)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_173),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_182),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_305),
.Y(n_361)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_145),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_156),
.A2(n_5),
.B1(n_8),
.B2(n_175),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_306),
.A2(n_314),
.B1(n_166),
.B2(n_152),
.Y(n_345)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_203),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_307),
.B(n_308),
.Y(n_363)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_184),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_158),
.B(n_135),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_309),
.B(n_311),
.Y(n_321)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_160),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_310),
.B(n_316),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_205),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_142),
.B(n_211),
.Y(n_312)
);

CKINVDCx12_ASAP7_75t_R g353 ( 
.A(n_312),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_151),
.B(n_176),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_313),
.B(n_315),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_154),
.A2(n_198),
.B1(n_147),
.B2(n_205),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_170),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_166),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_272),
.A2(n_230),
.B1(n_155),
.B2(n_229),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_318),
.A2(n_328),
.B1(n_334),
.B2(n_343),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_348),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_263),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_331),
.B(n_347),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_239),
.B(n_234),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_332),
.B(n_339),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_238),
.A2(n_229),
.B1(n_154),
.B2(n_212),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_333),
.A2(n_294),
.B1(n_297),
.B2(n_240),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_236),
.A2(n_249),
.B1(n_280),
.B2(n_241),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_261),
.B(n_186),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_249),
.A2(n_188),
.B1(n_213),
.B2(n_212),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_300),
.A2(n_171),
.B1(n_213),
.B2(n_188),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_344),
.A2(n_345),
.B1(n_362),
.B2(n_233),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_312),
.Y(n_347)
);

OR2x4_ASAP7_75t_L g354 ( 
.A(n_253),
.B(n_193),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_354),
.A2(n_369),
.B(n_325),
.C(n_319),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_279),
.B(n_199),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_355),
.B(n_365),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_288),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_247),
.A2(n_152),
.B1(n_163),
.B2(n_159),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_282),
.B(n_169),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_285),
.B(n_169),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_378),
.Y(n_381)
);

AOI32xp33_ASAP7_75t_L g369 ( 
.A1(n_274),
.A2(n_163),
.A3(n_216),
.B1(n_277),
.B2(n_260),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_235),
.B(n_271),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_379),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_271),
.A2(n_298),
.B1(n_232),
.B2(n_265),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_374),
.A2(n_322),
.B1(n_349),
.B2(n_346),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_312),
.B(n_243),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_380),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_374),
.A2(n_305),
.B1(n_290),
.B2(n_281),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_382),
.Y(n_447)
);

FAx1_ASAP7_75t_SL g383 ( 
.A(n_354),
.B(n_270),
.CI(n_265),
.CON(n_383),
.SN(n_383)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_383),
.B(n_419),
.Y(n_466)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_368),
.Y(n_384)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_330),
.B(n_319),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_385),
.B(n_398),
.Y(n_443)
);

AOI32xp33_ASAP7_75t_L g386 ( 
.A1(n_358),
.A2(n_303),
.A3(n_276),
.B1(n_270),
.B2(n_308),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_386),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_332),
.B(n_286),
.C(n_245),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_353),
.C(n_331),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_342),
.A2(n_265),
.B1(n_288),
.B2(n_302),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_389),
.A2(n_392),
.B1(n_393),
.B2(n_397),
.Y(n_432)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_368),
.Y(n_390)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_390),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_342),
.A2(n_346),
.B1(n_360),
.B2(n_348),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_394),
.B(n_399),
.Y(n_453)
);

AND2x2_ASAP7_75t_SL g396 ( 
.A(n_346),
.B(n_266),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_396),
.B(n_353),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_334),
.A2(n_288),
.B1(n_295),
.B2(n_301),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_330),
.B(n_242),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_310),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_328),
.A2(n_244),
.B1(n_246),
.B2(n_276),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_400),
.A2(n_403),
.B1(n_424),
.B2(n_414),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_321),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_401),
.B(n_412),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_337),
.Y(n_402)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_402),
.Y(n_445)
);

INVx3_ASAP7_75t_SL g404 ( 
.A(n_326),
.Y(n_404)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_404),
.Y(n_450)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_405),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_371),
.A2(n_262),
.B1(n_250),
.B2(n_255),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_406),
.A2(n_415),
.B1(n_417),
.B2(n_422),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_407),
.A2(n_416),
.B(n_418),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_409),
.A2(n_344),
.B1(n_415),
.B2(n_417),
.Y(n_434)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_411),
.Y(n_469)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_420),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_373),
.A2(n_256),
.B1(n_268),
.B2(n_293),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_369),
.B(n_292),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_367),
.A2(n_316),
.B1(n_257),
.B2(n_287),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_321),
.A2(n_266),
.B(n_252),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_329),
.B(n_252),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_378),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_423),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_371),
.A2(n_252),
.B1(n_355),
.B2(n_379),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_326),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_428),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_329),
.B(n_323),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_426),
.B(n_320),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_339),
.B(n_365),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_429),
.Y(n_463)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_433),
.B(n_468),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_434),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_440),
.C(n_452),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_416),
.A2(n_324),
.B1(n_318),
.B2(n_327),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_436),
.A2(n_438),
.B1(n_457),
.B2(n_387),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_416),
.A2(n_335),
.B(n_357),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_437),
.A2(n_462),
.B(n_386),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_424),
.A2(n_327),
.B1(n_343),
.B2(n_357),
.Y(n_438)
);

AO22x1_ASAP7_75t_L g439 ( 
.A1(n_392),
.A2(n_340),
.B1(n_335),
.B2(n_356),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_439),
.A2(n_408),
.B(n_418),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_385),
.B(n_317),
.C(n_340),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_393),
.A2(n_376),
.B(n_317),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_442),
.A2(n_418),
.B(n_407),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_397),
.A2(n_376),
.B1(n_375),
.B2(n_350),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_446),
.A2(n_449),
.B1(n_467),
.B2(n_429),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_387),
.A2(n_375),
.B1(n_364),
.B2(n_352),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_356),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_370),
.C(n_320),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_396),
.C(n_399),
.Y(n_482)
);

BUFx12_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_459),
.Y(n_478)
);

MAJx2_ASAP7_75t_L g461 ( 
.A(n_391),
.B(n_370),
.C(n_364),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_461),
.B(n_381),
.Y(n_494)
);

OAI22x1_ASAP7_75t_L g462 ( 
.A1(n_394),
.A2(n_352),
.B1(n_372),
.B2(n_341),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_391),
.B(n_338),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_465),
.B(n_419),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_387),
.A2(n_351),
.B1(n_366),
.B2(n_338),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_402),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_404),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_398),
.B(n_341),
.Y(n_471)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_471),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_473),
.A2(n_483),
.B1(n_486),
.B2(n_487),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_476),
.A2(n_481),
.B(n_485),
.Y(n_533)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_454),
.Y(n_477)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_477),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_479),
.B(n_492),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_426),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_480),
.B(n_498),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_482),
.B(n_435),
.C(n_433),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_432),
.A2(n_389),
.B1(n_394),
.B2(n_422),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_432),
.A2(n_427),
.B1(n_408),
.B2(n_395),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_436),
.A2(n_472),
.B1(n_438),
.B2(n_439),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_439),
.A2(n_395),
.B1(n_383),
.B2(n_410),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_488),
.A2(n_496),
.B1(n_502),
.B2(n_507),
.Y(n_535)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_454),
.Y(n_489)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_448),
.Y(n_490)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_463),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_493),
.A2(n_497),
.B1(n_499),
.B2(n_503),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_437),
.A2(n_399),
.B(n_383),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_495),
.B(n_505),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_460),
.A2(n_411),
.B1(n_420),
.B2(n_423),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_463),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_455),
.B(n_388),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_451),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_460),
.A2(n_425),
.B(n_396),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_500),
.A2(n_501),
.B(n_512),
.Y(n_523)
);

OAI32xp33_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_381),
.A3(n_405),
.B1(n_390),
.B2(n_428),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_446),
.A2(n_406),
.B1(n_396),
.B2(n_402),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_455),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_504),
.B(n_506),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_466),
.B(n_461),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_469),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_441),
.A2(n_384),
.B1(n_412),
.B2(n_380),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_508),
.A2(n_465),
.B1(n_449),
.B2(n_447),
.Y(n_526)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_469),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_444),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_441),
.A2(n_380),
.B1(n_351),
.B2(n_366),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_510),
.A2(n_507),
.B1(n_434),
.B2(n_478),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_464),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_511),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_453),
.A2(n_359),
.B(n_377),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_524),
.C(n_529),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_452),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_517),
.B(n_520),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_479),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_518),
.B(n_521),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_474),
.B(n_496),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_480),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_492),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_522),
.B(n_531),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_433),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_526),
.A2(n_483),
.B1(n_487),
.B2(n_475),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_484),
.A2(n_453),
.B1(n_443),
.B2(n_462),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_527),
.A2(n_532),
.B1(n_547),
.B2(n_476),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_482),
.B(n_458),
.C(n_440),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_512),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_484),
.A2(n_453),
.B1(n_443),
.B2(n_462),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_512),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_536),
.B(n_541),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_537),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_482),
.B(n_442),
.C(n_461),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_538),
.B(n_539),
.C(n_543),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_486),
.B(n_456),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_485),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_490),
.B(n_456),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_542),
.B(n_546),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_498),
.B(n_471),
.C(n_448),
.Y(n_543)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_544),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_485),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_545),
.B(n_491),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_494),
.B(n_464),
.C(n_430),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_473),
.A2(n_447),
.B1(n_467),
.B2(n_450),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_494),
.B(n_430),
.C(n_444),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_548),
.B(n_481),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_495),
.A2(n_450),
.B(n_470),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_551),
.A2(n_500),
.B(n_505),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_SL g552 ( 
.A(n_524),
.B(n_491),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g592 ( 
.A(n_552),
.B(n_515),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_553),
.A2(n_557),
.B1(n_584),
.B2(n_547),
.Y(n_601)
);

BUFx12_ASAP7_75t_L g556 ( 
.A(n_531),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_556),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_536),
.B(n_511),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_560),
.B(n_575),
.Y(n_612)
);

INVx13_ASAP7_75t_L g561 ( 
.A(n_551),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_533),
.A2(n_523),
.B(n_545),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_564),
.A2(n_580),
.B(n_550),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_565),
.B(n_566),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_534),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_535),
.A2(n_489),
.B1(n_477),
.B2(n_475),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_567),
.A2(n_569),
.B1(n_581),
.B2(n_582),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_535),
.A2(n_497),
.B1(n_493),
.B2(n_495),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_522),
.B(n_505),
.Y(n_570)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_570),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_514),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_572),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_514),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_521),
.B(n_488),
.Y(n_573)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_573),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_504),
.Y(n_574)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_574),
.Y(n_599)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_543),
.Y(n_576)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_576),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_523),
.Y(n_577)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_577),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_513),
.B(n_509),
.Y(n_578)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_578),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_549),
.A2(n_502),
.B1(n_510),
.B2(n_506),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_537),
.A2(n_513),
.B1(n_518),
.B2(n_541),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_527),
.A2(n_501),
.B1(n_508),
.B2(n_503),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_519),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_585),
.B(n_530),
.Y(n_588)
);

AOI22x1_ASAP7_75t_L g586 ( 
.A1(n_533),
.A2(n_499),
.B1(n_431),
.B2(n_478),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_SL g591 ( 
.A(n_586),
.B(n_560),
.C(n_582),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_583),
.B(n_520),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_587),
.B(n_594),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_588),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_554),
.A2(n_532),
.B1(n_519),
.B2(n_530),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_589),
.A2(n_600),
.B1(n_584),
.B2(n_581),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_579),
.B(n_529),
.C(n_517),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_590),
.B(n_605),
.Y(n_635)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_591),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_592),
.B(n_593),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_579),
.B(n_548),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_583),
.B(n_546),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_597),
.B(n_598),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_555),
.B(n_538),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_554),
.A2(n_516),
.B1(n_528),
.B2(n_526),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_601),
.A2(n_609),
.B1(n_569),
.B2(n_572),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_555),
.B(n_525),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_602),
.B(n_603),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_559),
.B(n_550),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_576),
.B(n_540),
.C(n_445),
.Y(n_605)
);

NOR3xp33_ASAP7_75t_SL g609 ( 
.A(n_562),
.B(n_540),
.C(n_445),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_608),
.B(n_566),
.Y(n_615)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_615),
.Y(n_646)
);

CKINVDCx16_ASAP7_75t_R g619 ( 
.A(n_604),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_619),
.A2(n_624),
.B1(n_632),
.B2(n_633),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_594),
.B(n_567),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_621),
.B(n_602),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_612),
.B(n_562),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_622),
.A2(n_628),
.B(n_630),
.Y(n_644)
);

BUFx24_ASAP7_75t_SL g623 ( 
.A(n_603),
.Y(n_623)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_623),
.Y(n_650)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_611),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_587),
.B(n_564),
.C(n_577),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_625),
.B(n_629),
.C(n_631),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_627),
.A2(n_554),
.B1(n_596),
.B2(n_570),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_612),
.B(n_578),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_598),
.B(n_568),
.C(n_552),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_614),
.B(n_571),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_590),
.B(n_568),
.C(n_560),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_609),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_593),
.B(n_586),
.C(n_563),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_634),
.B(n_607),
.C(n_610),
.Y(n_653)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_595),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_636),
.A2(n_637),
.B1(n_613),
.B2(n_558),
.Y(n_655)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_595),
.Y(n_637)
);

MAJx2_ASAP7_75t_L g639 ( 
.A(n_625),
.B(n_592),
.C(n_597),
.Y(n_639)
);

MAJx2_ASAP7_75t_L g668 ( 
.A(n_639),
.B(n_652),
.C(n_657),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_640),
.B(n_648),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_631),
.B(n_606),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_641),
.B(n_643),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_618),
.B(n_605),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_642),
.B(n_658),
.Y(n_669)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_638),
.B(n_601),
.Y(n_643)
);

NOR2x1_ASAP7_75t_L g647 ( 
.A(n_630),
.B(n_563),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_647),
.A2(n_556),
.B(n_561),
.Y(n_674)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_638),
.B(n_600),
.Y(n_648)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_618),
.B(n_634),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_649),
.B(n_654),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_SL g652 ( 
.A(n_621),
.B(n_580),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_653),
.B(n_626),
.Y(n_672)
);

XOR2xp5_ASAP7_75t_L g654 ( 
.A(n_629),
.B(n_589),
.Y(n_654)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_655),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_656),
.A2(n_627),
.B1(n_553),
.B2(n_599),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_620),
.A2(n_575),
.B(n_586),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_635),
.B(n_591),
.C(n_557),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_641),
.B(n_616),
.C(n_626),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_662),
.B(n_664),
.Y(n_677)
);

OAI321xp33_ASAP7_75t_L g663 ( 
.A1(n_644),
.A2(n_622),
.A3(n_628),
.B1(n_617),
.B2(n_585),
.C(n_558),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_663),
.A2(n_666),
.B1(n_675),
.B2(n_654),
.Y(n_679)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_646),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_647),
.A2(n_657),
.B(n_651),
.Y(n_667)
);

XNOR2xp5_ASAP7_75t_SL g685 ( 
.A(n_667),
.B(n_674),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_645),
.B(n_616),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_670),
.B(n_671),
.Y(n_684)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_653),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_672),
.B(n_341),
.Y(n_682)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_645),
.B(n_556),
.C(n_561),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_673),
.B(n_642),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_SL g675 ( 
.A1(n_658),
.A2(n_648),
.B1(n_643),
.B2(n_652),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_673),
.B(n_650),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_676),
.B(n_682),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_669),
.A2(n_649),
.B(n_639),
.Y(n_678)
);

AOI21x1_ASAP7_75t_SL g695 ( 
.A1(n_678),
.A2(n_681),
.B(n_687),
.Y(n_695)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_679),
.Y(n_688)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_680),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_SL g681 ( 
.A1(n_667),
.A2(n_556),
.B(n_640),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g683 ( 
.A(n_660),
.B(n_665),
.C(n_662),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_683),
.B(n_675),
.Y(n_691)
);

XOR2xp5_ASAP7_75t_L g686 ( 
.A(n_659),
.B(n_459),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_686),
.Y(n_696)
);

FAx1_ASAP7_75t_L g687 ( 
.A(n_668),
.B(n_459),
.CI(n_377),
.CON(n_687),
.SN(n_687)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_684),
.B(n_661),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_690),
.B(n_691),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_SL g692 ( 
.A1(n_677),
.A2(n_674),
.B(n_666),
.Y(n_692)
);

MAJx2_ASAP7_75t_L g699 ( 
.A(n_692),
.B(n_685),
.C(n_686),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_682),
.A2(n_660),
.B(n_665),
.Y(n_693)
);

OAI21x1_ASAP7_75t_SL g697 ( 
.A1(n_693),
.A2(n_687),
.B(n_668),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_697),
.B(n_700),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_694),
.B(n_659),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_698),
.B(n_699),
.Y(n_702)
);

MAJIxp5_ASAP7_75t_L g700 ( 
.A(n_688),
.B(n_685),
.C(n_459),
.Y(n_700)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_701),
.A2(n_689),
.B(n_695),
.C(n_696),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_704),
.A2(n_703),
.B(n_377),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_702),
.B(n_696),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_705),
.A2(n_706),
.B(n_336),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_707),
.A2(n_336),
.B(n_372),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_708),
.A2(n_336),
.B(n_341),
.Y(n_709)
);

MAJIxp5_ASAP7_75t_L g710 ( 
.A(n_709),
.B(n_336),
.C(n_372),
.Y(n_710)
);

XNOR2xp5_ASAP7_75t_L g711 ( 
.A(n_710),
.B(n_372),
.Y(n_711)
);


endmodule