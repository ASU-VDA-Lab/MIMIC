module fake_jpeg_26331_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_34),
.B1(n_19),
.B2(n_18),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_64),
.B1(n_41),
.B2(n_48),
.Y(n_98)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_68),
.Y(n_74)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_59),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_34),
.B1(n_19),
.B2(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_35),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_82),
.B(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_78),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_40),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_42),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_85),
.C(n_43),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_17),
.B(n_28),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_41),
.B1(n_38),
.B2(n_48),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_89),
.B1(n_93),
.B2(n_98),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_39),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_41),
.B1(n_34),
.B2(n_49),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_99),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_41),
.B1(n_19),
.B2(n_42),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_55),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_96),
.Y(n_129)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_106),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_63),
.B1(n_59),
.B2(n_54),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_97),
.B1(n_96),
.B2(n_90),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_118),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_23),
.B1(n_42),
.B2(n_45),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_93),
.B1(n_54),
.B2(n_51),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_120),
.Y(n_134)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_43),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_71),
.Y(n_121)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_43),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_85),
.B1(n_94),
.B2(n_99),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_132),
.B1(n_153),
.B2(n_101),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_38),
.C(n_92),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_44),
.Y(n_172)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_142),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_33),
.B(n_35),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_144),
.B(n_24),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_48),
.B1(n_45),
.B2(n_86),
.Y(n_171)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx5_ASAP7_75t_SL g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_155),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_33),
.B(n_69),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_69),
.B(n_47),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_150),
.B(n_154),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_89),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_158),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_100),
.B1(n_112),
.B2(n_128),
.Y(n_166)
);

AOI32xp33_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_45),
.A3(n_79),
.B1(n_72),
.B2(n_44),
.Y(n_150)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_59),
.B1(n_79),
.B2(n_100),
.Y(n_153)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_45),
.A3(n_44),
.B1(n_38),
.B2(n_43),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_156),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_49),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_113),
.B1(n_109),
.B2(n_101),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_166),
.B1(n_169),
.B2(n_171),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_161),
.A2(n_190),
.B1(n_31),
.B2(n_32),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_115),
.B1(n_122),
.B2(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_176),
.B1(n_187),
.B2(n_151),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_119),
.B(n_47),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_118),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_170),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_112),
.B1(n_100),
.B2(n_110),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_110),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_175),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_57),
.B1(n_116),
.B2(n_17),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_135),
.B(n_28),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_57),
.B1(n_86),
.B2(n_36),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_136),
.A2(n_20),
.B1(n_36),
.B2(n_27),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_86),
.B1(n_36),
.B2(n_27),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_36),
.B1(n_27),
.B2(n_20),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_133),
.A2(n_27),
.B1(n_20),
.B2(n_29),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_141),
.B1(n_152),
.B2(n_146),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_30),
.B(n_22),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_139),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_143),
.A2(n_30),
.B1(n_32),
.B2(n_2),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_145),
.B(n_32),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_32),
.Y(n_213)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_198),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_195),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_202),
.B1(n_166),
.B2(n_183),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_208),
.Y(n_226)
);

NOR4xp25_ASAP7_75t_SL g201 ( 
.A(n_186),
.B(n_150),
.C(n_137),
.D(n_145),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_214),
.B(n_220),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_155),
.B1(n_142),
.B2(n_148),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_138),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_146),
.C(n_156),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_191),
.C(n_172),
.Y(n_227)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_211),
.Y(n_240)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_218),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_161),
.A2(n_29),
.B1(n_25),
.B2(n_31),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_25),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_160),
.B(n_0),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_164),
.B(n_186),
.Y(n_239)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_16),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_223),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_209),
.C(n_202),
.Y(n_255)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_238),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_231),
.B1(n_242),
.B2(n_226),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_185),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_243),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_162),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

OA21x2_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_213),
.B(n_212),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_180),
.B1(n_177),
.B2(n_189),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_197),
.B1(n_196),
.B2(n_200),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_185),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_173),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_248),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_170),
.B(n_176),
.C(n_178),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_221),
.B(n_216),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_198),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_255),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_260),
.B1(n_264),
.B2(n_266),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_199),
.B1(n_192),
.B2(n_206),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_253),
.A2(n_257),
.B1(n_267),
.B2(n_248),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_216),
.C(n_196),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_268),
.C(n_270),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_197),
.B1(n_207),
.B2(n_208),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_231),
.A2(n_212),
.B1(n_187),
.B2(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_224),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_225),
.B1(n_238),
.B2(n_236),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_235),
.B(n_211),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_269),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_218),
.B1(n_210),
.B2(n_179),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_179),
.C(n_16),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_241),
.B(n_15),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_14),
.C(n_13),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_275),
.B1(n_276),
.B2(n_286),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_274),
.B(n_278),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_244),
.B1(n_228),
.B2(n_230),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_228),
.B1(n_232),
.B2(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_229),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_245),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_282),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_254),
.B1(n_259),
.B2(n_257),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_258),
.A2(n_233),
.B1(n_245),
.B2(n_239),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_246),
.C(n_240),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_284),
.C(n_11),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_14),
.C(n_13),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_254),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_13),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_3),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_3),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_253),
.B1(n_262),
.B2(n_269),
.Y(n_292)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_250),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_302),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_288),
.A2(n_265),
.B(n_250),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_295),
.A2(n_291),
.B(n_290),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_296)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_303),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_276),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_284),
.B1(n_273),
.B2(n_279),
.Y(n_306)
);

OA21x2_ASAP7_75t_SL g300 ( 
.A1(n_271),
.A2(n_10),
.B(n_4),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_300),
.A2(n_286),
.B(n_279),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_273),
.B(n_10),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_9),
.C(n_4),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_5),
.C(n_6),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_311),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_291),
.A2(n_3),
.B(n_4),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_308),
.B(n_309),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_315),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_298),
.A2(n_6),
.B(n_7),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_301),
.C(n_289),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_301),
.C(n_293),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_294),
.Y(n_322)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_302),
.Y(n_323)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_323),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_312),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_327),
.B(n_330),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_317),
.A2(n_297),
.B(n_314),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_328),
.A2(n_332),
.B(n_321),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_299),
.B1(n_306),
.B2(n_311),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_303),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_334),
.B(n_326),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_319),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_331),
.C(n_335),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_332),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_325),
.Y(n_339)
);

AOI321xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_295),
.A3(n_304),
.B1(n_309),
.B2(n_9),
.C(n_6),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_9),
.B(n_7),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_8),
.Y(n_342)
);


endmodule