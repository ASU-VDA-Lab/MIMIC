module fake_jpeg_19951_n_59 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_9),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_12),
.B1(n_23),
.B2(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_2),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.C(n_28),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_11),
.C(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_25),
.B1(n_27),
.B2(n_5),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_44),
.B(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_30),
.B1(n_7),
.B2(n_8),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_6),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_49),
.B1(n_51),
.B2(n_40),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_48),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_52),
.B1(n_46),
.B2(n_45),
.Y(n_56)
);

AOI21x1_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_13),
.B(n_14),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_15),
.C(n_17),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_19),
.B(n_24),
.Y(n_59)
);


endmodule