module fake_ibex_355_n_6427 (n_151, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_854, n_1008, n_458, n_244, n_73, n_343, n_310, n_714, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_1039, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_6427);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_1039;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_6427;

wire n_4557;
wire n_6210;
wire n_5285;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_5261;
wire n_5895;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_1078;
wire n_4422;
wire n_5743;
wire n_1865;
wire n_5033;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_1424;
wire n_2625;
wire n_2444;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_6114;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_3147;
wire n_3983;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6124;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_6136;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6128;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_6379;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_3796;
wire n_5719;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3477;
wire n_3070;
wire n_1575;
wire n_4416;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_3339;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_1517;
wire n_5973;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_5770;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2420;
wire n_2380;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_5566;
wire n_6185;
wire n_5342;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_1072;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_4919;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_4686;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_5384;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_6176;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_5097;
wire n_4688;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_2682;
wire n_1666;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4970;
wire n_4652;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_5983;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_6021;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_4610;
wire n_5854;
wire n_4067;
wire n_4997;
wire n_5906;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6117;
wire n_1312;
wire n_5844;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_6237;
wire n_4922;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_5488;
wire n_3107;
wire n_5465;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4965;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_3703;
wire n_5116;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_1775;
wire n_6361;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_5746;
wire n_5883;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_6062;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_1832;
wire n_3718;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_4878;
wire n_6252;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_1067;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_6398;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_5096;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5869;
wire n_5862;
wire n_1238;
wire n_3959;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_5277;
wire n_5900;
wire n_3647;
wire n_6240;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1669;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_1175;
wire n_4408;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_5645;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_2757;
wire n_1622;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_6380;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_5644;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_2168;
wire n_1442;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_5940;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_5324;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1780;
wire n_1091;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_6310;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_6249;
wire n_3559;
wire n_5184;
wire n_5747;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_5618;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_5464;
wire n_6420;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_2565;
wire n_4201;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4975;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_6025;
wire n_6168;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_1764;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_5123;
wire n_6160;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4126;
wire n_4103;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_2748;
wire n_5359;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_6140;
wire n_5903;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4681;
wire n_4253;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_5985;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_2300;
wire n_1120;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_4587;
wire n_6118;
wire n_6158;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1395;
wire n_1115;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_6049;
wire n_2419;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_5724;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_2458;
wire n_3401;
wire n_3032;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5595;
wire n_5334;
wire n_6260;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5725;
wire n_5034;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_2684;
wire n_2205;
wire n_1104;
wire n_3284;
wire n_2875;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_3960;
wire n_4007;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_1587;
wire n_2555;
wire n_6356;
wire n_5313;
wire n_2108;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_6225;
wire n_1642;
wire n_5744;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6364;
wire n_5715;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_2157;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_5853;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_1060;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_3989;
wire n_5565;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_1336;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6167;
wire n_6189;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5984;
wire n_6385;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_6015;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_2374;
wire n_1614;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6376;
wire n_2571;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_6132;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6089;
wire n_5211;
wire n_1668;
wire n_5861;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3896;
wire n_3533;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5430;
wire n_5182;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6175;
wire n_5279;
wire n_4650;
wire n_6415;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_6046;
wire n_1326;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_5720;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_5561;
wire n_4762;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_5682;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1566;
wire n_1464;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6214;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5855;
wire n_5819;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_3449;
wire n_2923;
wire n_2990;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_5992;
wire n_5105;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_6099;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_3747;
wire n_1323;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1458;
wire n_1694;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_5485;
wire n_5737;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_6250;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5349;
wire n_5054;
wire n_1167;
wire n_3231;
wire n_6423;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_1088;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_5298;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_4811;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_2870;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_2928;
wire n_3557;
wire n_1193;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_6261;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_5393;
wire n_4782;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

INVx1_ASAP7_75t_L g1043 ( 
.A(n_981),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_875),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_476),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_923),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_115),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_959),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_255),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_416),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_476),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_21),
.Y(n_1052)
);

INVx1_ASAP7_75t_SL g1053 ( 
.A(n_1007),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_201),
.Y(n_1054)
);

CKINVDCx14_ASAP7_75t_R g1055 ( 
.A(n_407),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_231),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_936),
.Y(n_1057)
);

INVxp33_ASAP7_75t_L g1058 ( 
.A(n_456),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_302),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_525),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_813),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_845),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_193),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_375),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_916),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_51),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_144),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_836),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_431),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_843),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_806),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_998),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_218),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_548),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_820),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_323),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_243),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_945),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_646),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_783),
.Y(n_1080)
);

CKINVDCx6p67_ASAP7_75t_R g1081 ( 
.A(n_50),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_940),
.Y(n_1082)
);

BUFx5_ASAP7_75t_L g1083 ( 
.A(n_29),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_44),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_787),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_3),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_29),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_398),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_304),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_119),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_973),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_382),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_417),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_629),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_849),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_986),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_634),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_892),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1033),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_827),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_848),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_982),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_122),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_947),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_238),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_23),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_546),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_703),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_271),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_73),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1008),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_427),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_45),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_655),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1003),
.Y(n_1115)
);

BUFx10_ASAP7_75t_L g1116 ( 
.A(n_1017),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_966),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_978),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_501),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1006),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_586),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_346),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_767),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_971),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_253),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1012),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_521),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_809),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_512),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_233),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_418),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_933),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_720),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_350),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_804),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_182),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1042),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_593),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_324),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_41),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_507),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_241),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_271),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_945),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1001),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1017),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_194),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_281),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_160),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_480),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_763),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_994),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_526),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_496),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_602),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_887),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_179),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_874),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_907),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_834),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_348),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_35),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_991),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_756),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_941),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_755),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_377),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_176),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_910),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_427),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_78),
.Y(n_1171)
);

BUFx10_ASAP7_75t_L g1172 ( 
.A(n_20),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_906),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_665),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_98),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_924),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1036),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_933),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_70),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_294),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_962),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_989),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_207),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_723),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_889),
.Y(n_1185)
);

CKINVDCx14_ASAP7_75t_R g1186 ( 
.A(n_125),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_317),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_718),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_414),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_69),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_13),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_729),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_605),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_388),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_917),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_918),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_913),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_900),
.Y(n_1198)
);

BUFx5_ASAP7_75t_L g1199 ( 
.A(n_989),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_707),
.Y(n_1200)
);

BUFx2_ASAP7_75t_SL g1201 ( 
.A(n_110),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_910),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_293),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_921),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_172),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_563),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_92),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_908),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_304),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_213),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_752),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_20),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_873),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_819),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1030),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_358),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_443),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1003),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_371),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_961),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_484),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_495),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_122),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1039),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_353),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_742),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_680),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_310),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_407),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_731),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_97),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_991),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_660),
.Y(n_1233)
);

BUFx10_ASAP7_75t_L g1234 ( 
.A(n_93),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_437),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_282),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_824),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_912),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_356),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_828),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1001),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_964),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_214),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_883),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_278),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_141),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_582),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_446),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_752),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_874),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_417),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_72),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_681),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_935),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_646),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_279),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_960),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_486),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_429),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_976),
.Y(n_1260)
);

CKINVDCx16_ASAP7_75t_R g1261 ( 
.A(n_935),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_308),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1035),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_161),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_735),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_376),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_938),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_836),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_291),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_705),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1013),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_69),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1002),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_3),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_223),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_621),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_415),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_154),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_237),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_135),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_564),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_658),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_732),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_808),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_18),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1010),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_673),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_548),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1023),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_681),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_167),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_789),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_665),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_942),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_712),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_675),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_856),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_81),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_61),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_719),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_251),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_970),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1019),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_397),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_723),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_598),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_905),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_436),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_291),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_920),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_388),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_803),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_326),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_921),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_643),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_930),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_972),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_993),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_619),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_67),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_986),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_995),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_141),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_841),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_929),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_224),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_678),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_355),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_229),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_728),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_123),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_51),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_958),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_915),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_955),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_831),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_950),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_901),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1029),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_845),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_949),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_339),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_466),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_953),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_954),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_2),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_434),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_411),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1028),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_614),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_677),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_64),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1034),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_888),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_53),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_48),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_330),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_907),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_380),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_440),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_467),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_258),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_810),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_977),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_893),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_952),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_266),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_889),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_504),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_703),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_992),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_951),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_866),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_763),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_467),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_523),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_914),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_396),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_250),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_807),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_811),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_965),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1018),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_801),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_693),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_380),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_919),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_928),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_996),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_963),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_854),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_920),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_265),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_438),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_257),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_349),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_990),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_283),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_674),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_774),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_402),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_73),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_602),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_42),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_324),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_367),
.Y(n_1406)
);

BUFx10_ASAP7_75t_L g1407 ( 
.A(n_442),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_769),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_207),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_157),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_642),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_233),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_164),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_50),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_119),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_956),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_526),
.Y(n_1417)
);

BUFx2_ASAP7_75t_SL g1418 ( 
.A(n_728),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_258),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_251),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_56),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1037),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_807),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_815),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_897),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_842),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_427),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_982),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_388),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_719),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_167),
.Y(n_1431)
);

BUFx5_ASAP7_75t_L g1432 ( 
.A(n_269),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_284),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_776),
.Y(n_1434)
);

CKINVDCx16_ASAP7_75t_R g1435 ( 
.A(n_447),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_58),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_722),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_211),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_398),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_65),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_983),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1006),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_225),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_422),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1020),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_737),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_974),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_776),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_967),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_815),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_392),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_292),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_700),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_458),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1009),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_664),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_955),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_19),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_82),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_395),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_351),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_847),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_689),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_898),
.Y(n_1464)
);

CKINVDCx14_ASAP7_75t_R g1465 ( 
.A(n_604),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1033),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_864),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_968),
.Y(n_1468)
);

BUFx10_ASAP7_75t_L g1469 ( 
.A(n_932),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_488),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_579),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_476),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_695),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_834),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_988),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1012),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_751),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_513),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_71),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_628),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_246),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_925),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_962),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_984),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_944),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_484),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_17),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1026),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_810),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_519),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_390),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1024),
.Y(n_1492)
);

BUFx10_ASAP7_75t_L g1493 ( 
.A(n_909),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1011),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_888),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_433),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_697),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_699),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1040),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_943),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_111),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_7),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_200),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_107),
.Y(n_1504)
);

INVxp33_ASAP7_75t_R g1505 ( 
.A(n_531),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_902),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_328),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_135),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_778),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_957),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_428),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_355),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_181),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_937),
.Y(n_1514)
);

BUFx10_ASAP7_75t_L g1515 ( 
.A(n_310),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_946),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_482),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_884),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_627),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_28),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_13),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_705),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1004),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_568),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_523),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_122),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_188),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_38),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_902),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_44),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_975),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1038),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_655),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_960),
.Y(n_1534)
);

INVxp67_ASAP7_75t_SL g1535 ( 
.A(n_346),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_997),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_987),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_563),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1031),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_438),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_393),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_731),
.Y(n_1542)
);

INVx1_ASAP7_75t_SL g1543 ( 
.A(n_201),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_667),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_568),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_894),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_677),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1020),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_899),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_906),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_244),
.Y(n_1551)
);

INVx2_ASAP7_75t_R g1552 ( 
.A(n_227),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_905),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_983),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_123),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_514),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_880),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_844),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_145),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_664),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_733),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_192),
.Y(n_1562)
);

CKINVDCx14_ASAP7_75t_R g1563 ( 
.A(n_490),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_118),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_609),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_679),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_153),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_629),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_148),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_189),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_85),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_787),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_505),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_97),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_436),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_161),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_290),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_495),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_531),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_908),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_850),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1022),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_553),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_904),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_957),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_773),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_828),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_980),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_943),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_629),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_191),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_28),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_5),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_436),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_171),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_818),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_969),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_106),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_406),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1000),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_784),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1013),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_746),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_231),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_456),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_810),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_420),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_926),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_452),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_511),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_621),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_90),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1041),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_896),
.Y(n_1615)
);

CKINVDCx14_ASAP7_75t_R g1616 ( 
.A(n_931),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_856),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_961),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_465),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_670),
.Y(n_1620)
);

CKINVDCx20_ASAP7_75t_R g1621 ( 
.A(n_948),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_927),
.Y(n_1622)
);

BUFx8_ASAP7_75t_SL g1623 ( 
.A(n_922),
.Y(n_1623)
);

BUFx8_ASAP7_75t_SL g1624 ( 
.A(n_1037),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_555),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_993),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_759),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_40),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_373),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_318),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_227),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1026),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_858),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_5),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_15),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_75),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_416),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1015),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_59),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1032),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_622),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_366),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_74),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_498),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1005),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_679),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_321),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1027),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_58),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_528),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_245),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_769),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_527),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_236),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_631),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_361),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_647),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_623),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_794),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_151),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_299),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_816),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_911),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_416),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_30),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_851),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_972),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_975),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_128),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_826),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_934),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_183),
.Y(n_1672)
);

CKINVDCx14_ASAP7_75t_R g1673 ( 
.A(n_247),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_344),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1014),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_745),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_296),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_939),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_979),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_166),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_812),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1004),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_903),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_804),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_203),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_282),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_110),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_229),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_191),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_761),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_610),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_275),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_313),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_431),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_895),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_533),
.Y(n_1696)
);

CKINVDCx14_ASAP7_75t_R g1697 ( 
.A(n_887),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_377),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_47),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_230),
.Y(n_1700)
);

BUFx10_ASAP7_75t_L g1701 ( 
.A(n_285),
.Y(n_1701)
);

CKINVDCx20_ASAP7_75t_R g1702 ( 
.A(n_781),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_516),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_633),
.Y(n_1704)
);

CKINVDCx20_ASAP7_75t_R g1705 ( 
.A(n_1016),
.Y(n_1705)
);

CKINVDCx20_ASAP7_75t_R g1706 ( 
.A(n_302),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_316),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_985),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_482),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_570),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_454),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_147),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_380),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_206),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_835),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_678),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_220),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_84),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_999),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_596),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1023),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_676),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_724),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_870),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1021),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1025),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_98),
.Y(n_1727)
);

INVxp67_ASAP7_75t_SL g1728 ( 
.A(n_1058),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1055),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1113),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1078),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1396),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1628),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1629),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1635),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1656),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1714),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1109),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1055),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1186),
.Y(n_1740)
);

INVxp33_ASAP7_75t_SL g1741 ( 
.A(n_1093),
.Y(n_1741)
);

INVxp33_ASAP7_75t_L g1742 ( 
.A(n_1342),
.Y(n_1742)
);

INVxp33_ASAP7_75t_SL g1743 ( 
.A(n_1463),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1058),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1331),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1366),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1717),
.Y(n_1747)
);

CKINVDCx16_ASAP7_75t_R g1748 ( 
.A(n_1183),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1186),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1363),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1473),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1555),
.Y(n_1752)
);

INVxp33_ASAP7_75t_SL g1753 ( 
.A(n_1566),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1599),
.Y(n_1754)
);

CKINVDCx20_ASAP7_75t_R g1755 ( 
.A(n_1465),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1654),
.Y(n_1756)
);

INVxp33_ASAP7_75t_L g1757 ( 
.A(n_1644),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1685),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1130),
.Y(n_1759)
);

CKINVDCx16_ASAP7_75t_R g1760 ( 
.A(n_1435),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1465),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_1563),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1130),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1563),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1151),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1673),
.Y(n_1766)
);

INVxp67_ASAP7_75t_SL g1767 ( 
.A(n_1151),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1050),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1054),
.Y(n_1769)
);

CKINVDCx20_ASAP7_75t_R g1770 ( 
.A(n_1673),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1060),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1063),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1064),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1069),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1074),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1085),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1086),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1088),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1090),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1103),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1081),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1105),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1112),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1616),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1122),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1123),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1129),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1131),
.Y(n_1788)
);

BUFx2_ASAP7_75t_SL g1789 ( 
.A(n_1172),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1133),
.Y(n_1790)
);

CKINVDCx14_ASAP7_75t_R g1791 ( 
.A(n_1616),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1697),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1140),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1147),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1157),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1172),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1161),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1089),
.Y(n_1798)
);

CKINVDCx20_ASAP7_75t_R g1799 ( 
.A(n_1079),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1697),
.Y(n_1800)
);

CKINVDCx16_ASAP7_75t_R g1801 ( 
.A(n_1172),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1162),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1199),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1079),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1168),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1170),
.Y(n_1806)
);

INVxp33_ASAP7_75t_L g1807 ( 
.A(n_1218),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1175),
.Y(n_1808)
);

CKINVDCx20_ASAP7_75t_R g1809 ( 
.A(n_1384),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1192),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1234),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1200),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1623),
.Y(n_1813)
);

CKINVDCx16_ASAP7_75t_R g1814 ( 
.A(n_1234),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1203),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1205),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1078),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1209),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1212),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1217),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1222),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_1623),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1199),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1226),
.Y(n_1824)
);

INVxp33_ASAP7_75t_L g1825 ( 
.A(n_1601),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1624),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1624),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1228),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1231),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1457),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1045),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1246),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1632),
.Y(n_1833)
);

CKINVDCx16_ASAP7_75t_R g1834 ( 
.A(n_1234),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1089),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1199),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1116),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1248),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1047),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1252),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1264),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1266),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1270),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1407),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1051),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1384),
.Y(n_1846)
);

INVxp33_ASAP7_75t_L g1847 ( 
.A(n_1043),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1272),
.Y(n_1848)
);

CKINVDCx20_ASAP7_75t_R g1849 ( 
.A(n_1413),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1199),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1283),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1121),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1052),
.Y(n_1853)
);

CKINVDCx16_ASAP7_75t_R g1854 ( 
.A(n_1407),
.Y(n_1854)
);

INVxp33_ASAP7_75t_L g1855 ( 
.A(n_1048),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1290),
.Y(n_1856)
);

BUFx3_ASAP7_75t_L g1857 ( 
.A(n_1366),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1407),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1299),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1078),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1304),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1308),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1351),
.Y(n_1863)
);

INVxp33_ASAP7_75t_L g1864 ( 
.A(n_1057),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_1413),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1357),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1515),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1600),
.Y(n_1868)
);

CKINVDCx14_ASAP7_75t_R g1869 ( 
.A(n_1515),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1360),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1370),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1378),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1379),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1515),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1491),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1380),
.Y(n_1876)
);

OA21x2_ASAP7_75t_L g1877 ( 
.A1(n_1803),
.A2(n_1219),
.B(n_1148),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1742),
.A2(n_1261),
.B1(n_1498),
.B2(n_1491),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1746),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1869),
.Y(n_1880)
);

OA21x2_ASAP7_75t_L g1881 ( 
.A1(n_1823),
.A2(n_1219),
.B(n_1148),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1801),
.Y(n_1882)
);

BUFx8_ASAP7_75t_L g1883 ( 
.A(n_1738),
.Y(n_1883)
);

INVx6_ASAP7_75t_L g1884 ( 
.A(n_1814),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1867),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1867),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1731),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1741),
.A2(n_1501),
.B1(n_1508),
.B2(n_1498),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1757),
.B(n_1701),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1728),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1744),
.A2(n_1056),
.B1(n_1061),
.B2(n_1059),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1765),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1767),
.B(n_1066),
.Y(n_1893)
);

OAI21x1_ASAP7_75t_L g1894 ( 
.A1(n_1836),
.A2(n_1280),
.B(n_1243),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1731),
.Y(n_1895)
);

XNOR2x2_ASAP7_75t_L g1896 ( 
.A(n_1796),
.B(n_1505),
.Y(n_1896)
);

NOR2x1_ASAP7_75t_L g1897 ( 
.A(n_1789),
.B(n_1745),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1834),
.B(n_1083),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1857),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1730),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1759),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1763),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1854),
.Y(n_1903)
);

INVx5_ASAP7_75t_L g1904 ( 
.A(n_1837),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1798),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1835),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1852),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1732),
.Y(n_1908)
);

OA21x2_ASAP7_75t_L g1909 ( 
.A1(n_1850),
.A2(n_1280),
.B(n_1243),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1731),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1817),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1817),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1733),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_L g1914 ( 
.A1(n_1743),
.A2(n_1508),
.B1(n_1509),
.B2(n_1501),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1796),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1734),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1748),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1831),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1858),
.B(n_1067),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1735),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1736),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1817),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1811),
.B(n_1071),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1747),
.B(n_1182),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1860),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1860),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1737),
.Y(n_1927)
);

INVx4_ASAP7_75t_L g1928 ( 
.A(n_1729),
.Y(n_1928)
);

INVx5_ASAP7_75t_L g1929 ( 
.A(n_1860),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1768),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1769),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1807),
.B(n_1825),
.Y(n_1932)
);

INVx5_ASAP7_75t_L g1933 ( 
.A(n_1760),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1839),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1799),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1771),
.Y(n_1936)
);

INVx4_ASAP7_75t_L g1937 ( 
.A(n_1739),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1772),
.Y(n_1938)
);

AOI22x1_ASAP7_75t_SL g1939 ( 
.A1(n_1804),
.A2(n_1567),
.B1(n_1593),
.B2(n_1509),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1750),
.B(n_1683),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1773),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1774),
.Y(n_1942)
);

OA21x2_ASAP7_75t_L g1943 ( 
.A1(n_1876),
.A2(n_1776),
.B(n_1775),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1777),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1844),
.B(n_1874),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1845),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1778),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1753),
.B(n_1073),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1751),
.B(n_1382),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1749),
.A2(n_1076),
.B1(n_1080),
.B2(n_1077),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1853),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1779),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1780),
.Y(n_1953)
);

BUFx2_ASAP7_75t_L g1954 ( 
.A(n_1740),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1782),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1868),
.B(n_1084),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1783),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1791),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_SL g1959 ( 
.A(n_1764),
.B(n_1701),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1785),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1786),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1766),
.B(n_1087),
.Y(n_1962)
);

OA21x2_ASAP7_75t_L g1963 ( 
.A1(n_1787),
.A2(n_1315),
.B(n_1312),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1788),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1752),
.B(n_1382),
.Y(n_1965)
);

AND2x6_ASAP7_75t_L g1966 ( 
.A(n_1754),
.B(n_1121),
.Y(n_1966)
);

XNOR2x2_ASAP7_75t_L g1967 ( 
.A(n_1756),
.B(n_1210),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1790),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1793),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1794),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1795),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1833),
.B(n_1094),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1797),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1802),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1758),
.B(n_1589),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1830),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1805),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1806),
.Y(n_1978)
);

AND2x6_ASAP7_75t_L g1979 ( 
.A(n_1808),
.B(n_1223),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1810),
.B(n_1097),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1812),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1815),
.Y(n_1982)
);

INVx6_ASAP7_75t_L g1983 ( 
.A(n_1847),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1816),
.B(n_1106),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1818),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_SL g1986 ( 
.A1(n_1809),
.A2(n_1849),
.B1(n_1865),
.B2(n_1846),
.Y(n_1986)
);

CKINVDCx16_ASAP7_75t_R g1987 ( 
.A(n_1755),
.Y(n_1987)
);

OAI21x1_ASAP7_75t_L g1988 ( 
.A1(n_1819),
.A2(n_1315),
.B(n_1312),
.Y(n_1988)
);

BUFx12f_ASAP7_75t_L g1989 ( 
.A(n_1781),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1820),
.B(n_1108),
.Y(n_1990)
);

CKINVDCx5p33_ASAP7_75t_R g1991 ( 
.A(n_1813),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1761),
.B(n_1589),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1855),
.B(n_1701),
.Y(n_1993)
);

OA21x2_ASAP7_75t_L g1994 ( 
.A1(n_1821),
.A2(n_1472),
.B(n_1423),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1824),
.Y(n_1995)
);

CKINVDCx8_ASAP7_75t_R g1996 ( 
.A(n_1822),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1828),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1762),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1864),
.B(n_1223),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1829),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1832),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1838),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1784),
.B(n_1277),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1840),
.Y(n_2004)
);

INVxp33_ASAP7_75t_SL g2005 ( 
.A(n_1792),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1841),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1842),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1800),
.B(n_1770),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1843),
.B(n_1110),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1848),
.B(n_1114),
.Y(n_2010)
);

OA21x2_ASAP7_75t_L g2011 ( 
.A1(n_1851),
.A2(n_1472),
.B(n_1423),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1856),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1859),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1861),
.B(n_1277),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1862),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1863),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1866),
.B(n_1348),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1870),
.B(n_1348),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1871),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1826),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1872),
.Y(n_2021)
);

BUFx3_ASAP7_75t_L g2022 ( 
.A(n_1873),
.Y(n_2022)
);

INVx3_ASAP7_75t_L g2023 ( 
.A(n_1827),
.Y(n_2023)
);

NAND2xp33_ASAP7_75t_L g2024 ( 
.A(n_1875),
.B(n_1083),
.Y(n_2024)
);

CKINVDCx8_ASAP7_75t_R g2025 ( 
.A(n_1801),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1742),
.B(n_1356),
.Y(n_2026)
);

AND2x6_ASAP7_75t_L g2027 ( 
.A(n_1796),
.B(n_1356),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1728),
.Y(n_2028)
);

OA21x2_ASAP7_75t_L g2029 ( 
.A1(n_1803),
.A2(n_1530),
.B(n_1522),
.Y(n_2029)
);

OA21x2_ASAP7_75t_L g2030 ( 
.A1(n_1803),
.A2(n_1530),
.B(n_1522),
.Y(n_2030)
);

OA21x2_ASAP7_75t_L g2031 ( 
.A1(n_1803),
.A2(n_1580),
.B(n_1551),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1731),
.Y(n_2032)
);

NAND2xp33_ASAP7_75t_L g2033 ( 
.A(n_1729),
.B(n_1083),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1728),
.Y(n_2034)
);

OAI22x1_ASAP7_75t_L g2035 ( 
.A1(n_1813),
.A2(n_1593),
.B1(n_1602),
.B2(n_1567),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1746),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1728),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1728),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1746),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1746),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1731),
.Y(n_2041)
);

INVx3_ASAP7_75t_L g2042 ( 
.A(n_1867),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1728),
.Y(n_2043)
);

BUFx2_ASAP7_75t_L g2044 ( 
.A(n_1869),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1746),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1728),
.B(n_1421),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1746),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1731),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1742),
.B(n_1421),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_1869),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1869),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1746),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1728),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1742),
.B(n_1569),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1728),
.A2(n_1127),
.B1(n_1128),
.B2(n_1125),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1746),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1867),
.B(n_1134),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1728),
.B(n_1135),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1728),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1731),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1731),
.Y(n_2061)
);

BUFx8_ASAP7_75t_L g2062 ( 
.A(n_1738),
.Y(n_2062)
);

INVx6_ASAP7_75t_L g2063 ( 
.A(n_1801),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1731),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1746),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1867),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1728),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1728),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1728),
.B(n_1136),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1746),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_SL g2071 ( 
.A1(n_1799),
.A2(n_1606),
.B1(n_1713),
.B2(n_1602),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1728),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_1867),
.B(n_1138),
.Y(n_2073)
);

INVx3_ASAP7_75t_L g2074 ( 
.A(n_1867),
.Y(n_2074)
);

INVx3_ASAP7_75t_L g2075 ( 
.A(n_1867),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1746),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1728),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1728),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_1869),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_L g2080 ( 
.A(n_1731),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1801),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_L g2082 ( 
.A1(n_1803),
.A2(n_1580),
.B(n_1551),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_1869),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_1741),
.A2(n_1713),
.B1(n_1606),
.B2(n_1143),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1728),
.B(n_1569),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_SL g2086 ( 
.A1(n_1799),
.A2(n_1092),
.B1(n_1107),
.B2(n_1049),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1728),
.B(n_1142),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1731),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_1869),
.Y(n_2089)
);

BUFx6f_ASAP7_75t_L g2090 ( 
.A(n_1731),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1746),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1746),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1731),
.Y(n_2093)
);

BUFx6f_ASAP7_75t_L g2094 ( 
.A(n_1731),
.Y(n_2094)
);

BUFx2_ASAP7_75t_L g2095 ( 
.A(n_1869),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1728),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_1869),
.Y(n_2097)
);

INVx3_ASAP7_75t_L g2098 ( 
.A(n_1867),
.Y(n_2098)
);

INVxp67_ASAP7_75t_L g2099 ( 
.A(n_1728),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1731),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1728),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1746),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1746),
.Y(n_2103)
);

AOI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1741),
.A2(n_1150),
.B1(n_1153),
.B2(n_1149),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1728),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1746),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1742),
.B(n_1630),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1728),
.B(n_1630),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1728),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1731),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_1728),
.A2(n_1164),
.B1(n_1167),
.B2(n_1155),
.Y(n_2111)
);

OA21x2_ASAP7_75t_L g2112 ( 
.A1(n_1803),
.A2(n_1660),
.B(n_1647),
.Y(n_2112)
);

OA21x2_ASAP7_75t_L g2113 ( 
.A1(n_1803),
.A2(n_1660),
.B(n_1647),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1746),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1920),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1983),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1988),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1921),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_1943),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1880),
.Y(n_2120)
);

CKINVDCx20_ASAP7_75t_R g2121 ( 
.A(n_1935),
.Y(n_2121)
);

CKINVDCx20_ASAP7_75t_R g2122 ( 
.A(n_1882),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1927),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_1932),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_2050),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_2051),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_2089),
.Y(n_2127)
);

BUFx2_ASAP7_75t_L g2128 ( 
.A(n_1915),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1999),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_2025),
.Y(n_2130)
);

CKINVDCx16_ASAP7_75t_R g2131 ( 
.A(n_2083),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1908),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_2044),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1988),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_2079),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_2095),
.Y(n_2136)
);

NOR2xp67_ASAP7_75t_L g2137 ( 
.A(n_1933),
.B(n_2081),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_R g2138 ( 
.A(n_1917),
.B(n_1119),
.Y(n_2138)
);

BUFx2_ASAP7_75t_L g2139 ( 
.A(n_1976),
.Y(n_2139)
);

CKINVDCx5p33_ASAP7_75t_R g2140 ( 
.A(n_1934),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1963),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1994),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2011),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_1946),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1894),
.Y(n_2145)
);

INVx1_ASAP7_75t_SL g2146 ( 
.A(n_2026),
.Y(n_2146)
);

BUFx2_ASAP7_75t_L g2147 ( 
.A(n_1903),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_1993),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_1951),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2049),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1885),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1877),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_1884),
.Y(n_2153)
);

BUFx8_ASAP7_75t_SL g2154 ( 
.A(n_1989),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_2063),
.Y(n_2155)
);

HB1xp67_ASAP7_75t_L g2156 ( 
.A(n_2054),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2107),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_2097),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_1991),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_1986),
.Y(n_2160)
);

NAND2xp33_ASAP7_75t_R g2161 ( 
.A(n_2005),
.B(n_1171),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1996),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1987),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1939),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_R g2165 ( 
.A(n_1959),
.B(n_1139),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_1933),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_R g2167 ( 
.A(n_2023),
.B(n_1141),
.Y(n_2167)
);

BUFx10_ASAP7_75t_L g2168 ( 
.A(n_2027),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1883),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_2062),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_2071),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_R g2172 ( 
.A(n_1954),
.B(n_1154),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_1888),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1913),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1881),
.Y(n_2175)
);

AOI21x1_ASAP7_75t_L g2176 ( 
.A1(n_2082),
.A2(n_1405),
.B(n_1395),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1916),
.Y(n_2177)
);

INVxp67_ASAP7_75t_SL g2178 ( 
.A(n_2022),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_1914),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_2084),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_1889),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_2086),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2018),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_1998),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1918),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1909),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1901),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_1897),
.B(n_1535),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2029),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1902),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_2020),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2030),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1931),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1950),
.Y(n_2194)
);

NAND2x1_ASAP7_75t_L g2195 ( 
.A(n_1979),
.B(n_1674),
.Y(n_2195)
);

CKINVDCx20_ASAP7_75t_R g2196 ( 
.A(n_2104),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1958),
.Y(n_2197)
);

CKINVDCx16_ASAP7_75t_R g2198 ( 
.A(n_2008),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1891),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_2055),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1931),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_2099),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2031),
.Y(n_2203)
);

CKINVDCx20_ASAP7_75t_R g2204 ( 
.A(n_1948),
.Y(n_2204)
);

INVx3_ASAP7_75t_L g2205 ( 
.A(n_1886),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1956),
.B(n_1116),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1938),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_2111),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1938),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1896),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_1928),
.Y(n_2211)
);

CKINVDCx20_ASAP7_75t_R g2212 ( 
.A(n_1923),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1937),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_L g2214 ( 
.A(n_1890),
.B(n_1174),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_2035),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_2027),
.Y(n_2216)
);

NOR2x1p5_ASAP7_75t_L g2217 ( 
.A(n_1992),
.B(n_1179),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2112),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1941),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_2027),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1966),
.Y(n_2221)
);

AO21x2_ASAP7_75t_L g2222 ( 
.A1(n_2082),
.A2(n_1410),
.B(n_1406),
.Y(n_2222)
);

INVx1_ASAP7_75t_SL g2223 ( 
.A(n_2058),
.Y(n_2223)
);

CKINVDCx20_ASAP7_75t_R g2224 ( 
.A(n_1945),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1966),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1941),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_R g2227 ( 
.A(n_2024),
.B(n_1194),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1966),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_1967),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2046),
.Y(n_2230)
);

CKINVDCx20_ASAP7_75t_R g2231 ( 
.A(n_1972),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_1919),
.Y(n_2232)
);

INVx1_ASAP7_75t_SL g2233 ( 
.A(n_2069),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2113),
.Y(n_2234)
);

BUFx10_ASAP7_75t_L g2235 ( 
.A(n_2057),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_R g2236 ( 
.A(n_1979),
.B(n_1245),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1904),
.Y(n_2237)
);

AOI21x1_ASAP7_75t_L g2238 ( 
.A1(n_1980),
.A2(n_1417),
.B(n_1411),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_1904),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1973),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_1962),
.Y(n_2241)
);

CKINVDCx16_ASAP7_75t_R g2242 ( 
.A(n_2003),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1900),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_2087),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1973),
.Y(n_2245)
);

INVxp67_ASAP7_75t_L g2246 ( 
.A(n_1893),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_2028),
.Y(n_2247)
);

BUFx2_ASAP7_75t_L g2248 ( 
.A(n_1979),
.Y(n_2248)
);

CKINVDCx20_ASAP7_75t_R g2249 ( 
.A(n_1984),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_2034),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_2037),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_2038),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1977),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1977),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_2043),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_1978),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1978),
.Y(n_2257)
);

INVx3_ASAP7_75t_L g2258 ( 
.A(n_2042),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_2053),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_2066),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_2059),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1981),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_2067),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_2074),
.Y(n_2264)
);

CKINVDCx5p33_ASAP7_75t_R g2265 ( 
.A(n_2068),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1981),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2072),
.B(n_1116),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_2077),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_2078),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1995),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1995),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2096),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_2101),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_2105),
.Y(n_2274)
);

NAND2x1_ASAP7_75t_L g2275 ( 
.A(n_1942),
.B(n_1674),
.Y(n_2275)
);

CKINVDCx20_ASAP7_75t_R g2276 ( 
.A(n_1990),
.Y(n_2276)
);

BUFx10_ASAP7_75t_L g2277 ( 
.A(n_2073),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_2109),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2085),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_1892),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_2000),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_1898),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2000),
.Y(n_2283)
);

CKINVDCx20_ASAP7_75t_R g2284 ( 
.A(n_1878),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_2108),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_2014),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_1905),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_1906),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_1907),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_R g2290 ( 
.A(n_2033),
.B(n_1247),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_2009),
.Y(n_2291)
);

BUFx6f_ASAP7_75t_L g2292 ( 
.A(n_2012),
.Y(n_2292)
);

BUFx2_ASAP7_75t_L g2293 ( 
.A(n_2017),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_2010),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_1924),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1940),
.Y(n_2296)
);

CKINVDCx20_ASAP7_75t_R g2297 ( 
.A(n_2012),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_1949),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_R g2299 ( 
.A(n_2075),
.B(n_1251),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_1965),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2013),
.Y(n_2301)
);

HB1xp67_ASAP7_75t_L g2302 ( 
.A(n_2013),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2098),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_1975),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1879),
.Y(n_2305)
);

AOI21x1_ASAP7_75t_L g2306 ( 
.A1(n_1947),
.A2(n_1420),
.B(n_1419),
.Y(n_2306)
);

CKINVDCx20_ASAP7_75t_R g2307 ( 
.A(n_1952),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1899),
.Y(n_2308)
);

OAI21x1_ASAP7_75t_L g2309 ( 
.A1(n_1953),
.A2(n_1712),
.B(n_1688),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_1930),
.B(n_1242),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_2036),
.Y(n_2311)
);

NAND2xp33_ASAP7_75t_R g2312 ( 
.A(n_2114),
.B(n_1180),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_R g2313 ( 
.A(n_1955),
.B(n_1276),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_2039),
.Y(n_2314)
);

BUFx10_ASAP7_75t_L g2315 ( 
.A(n_1957),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2040),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_2045),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1936),
.Y(n_2318)
);

CKINVDCx20_ASAP7_75t_R g2319 ( 
.A(n_1961),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1944),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_2047),
.Y(n_2321)
);

CKINVDCx16_ASAP7_75t_R g2322 ( 
.A(n_1964),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_2052),
.Y(n_2323)
);

BUFx2_ASAP7_75t_L g2324 ( 
.A(n_1960),
.Y(n_2324)
);

CKINVDCx20_ASAP7_75t_R g2325 ( 
.A(n_1969),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_1970),
.B(n_1083),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_1968),
.B(n_1242),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_2056),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_R g2329 ( 
.A(n_1997),
.B(n_1301),
.Y(n_2329)
);

CKINVDCx20_ASAP7_75t_R g2330 ( 
.A(n_2001),
.Y(n_2330)
);

CKINVDCx5p33_ASAP7_75t_R g2331 ( 
.A(n_2065),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1971),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2070),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_R g2334 ( 
.A(n_2002),
.B(n_1319),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2076),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_2091),
.Y(n_2336)
);

CKINVDCx20_ASAP7_75t_R g2337 ( 
.A(n_2006),
.Y(n_2337)
);

CKINVDCx5p33_ASAP7_75t_R g2338 ( 
.A(n_2092),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1974),
.Y(n_2339)
);

CKINVDCx20_ASAP7_75t_R g2340 ( 
.A(n_2007),
.Y(n_2340)
);

BUFx6f_ASAP7_75t_L g2341 ( 
.A(n_2102),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_2103),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_2106),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_1982),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_1985),
.Y(n_2345)
);

CKINVDCx20_ASAP7_75t_R g2346 ( 
.A(n_2015),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_2004),
.Y(n_2347)
);

CKINVDCx8_ASAP7_75t_R g2348 ( 
.A(n_1929),
.Y(n_2348)
);

CKINVDCx20_ASAP7_75t_R g2349 ( 
.A(n_2019),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_2016),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2021),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1929),
.Y(n_2352)
);

NOR2xp67_ASAP7_75t_L g2353 ( 
.A(n_1887),
.B(n_0),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_1887),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1895),
.Y(n_2355)
);

CKINVDCx20_ASAP7_75t_R g2356 ( 
.A(n_1895),
.Y(n_2356)
);

CKINVDCx20_ASAP7_75t_R g2357 ( 
.A(n_1910),
.Y(n_2357)
);

NOR2x1p5_ASAP7_75t_L g2358 ( 
.A(n_1910),
.B(n_1184),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1911),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1911),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_1912),
.Y(n_2361)
);

HB1xp67_ASAP7_75t_L g2362 ( 
.A(n_1912),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_1922),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_1922),
.Y(n_2364)
);

INVxp33_ASAP7_75t_L g2365 ( 
.A(n_2110),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_1925),
.Y(n_2366)
);

CKINVDCx20_ASAP7_75t_R g2367 ( 
.A(n_1925),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_1926),
.Y(n_2368)
);

NAND2xp33_ASAP7_75t_R g2369 ( 
.A(n_1926),
.B(n_1187),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_2032),
.B(n_1188),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2032),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2041),
.Y(n_2372)
);

BUFx10_ASAP7_75t_L g2373 ( 
.A(n_2041),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_2048),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_2048),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2060),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_2060),
.B(n_1688),
.Y(n_2377)
);

INVx3_ASAP7_75t_L g2378 ( 
.A(n_2061),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2061),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_2064),
.Y(n_2380)
);

HB1xp67_ASAP7_75t_L g2381 ( 
.A(n_2064),
.Y(n_2381)
);

BUFx6f_ASAP7_75t_L g2382 ( 
.A(n_2110),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_2080),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_2080),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_2088),
.Y(n_2385)
);

BUFx3_ASAP7_75t_L g2386 ( 
.A(n_2088),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_2090),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_2090),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2093),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2093),
.Y(n_2390)
);

INVxp67_ASAP7_75t_L g2391 ( 
.A(n_2094),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_2094),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_2100),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_2100),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_1983),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_1932),
.B(n_1242),
.Y(n_2396)
);

CKINVDCx5p33_ASAP7_75t_R g2397 ( 
.A(n_1983),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_1983),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_1983),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_1983),
.Y(n_2400)
);

BUFx10_ASAP7_75t_L g2401 ( 
.A(n_1983),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1920),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_1983),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_1988),
.Y(n_2404)
);

NOR2xp33_ASAP7_75t_R g2405 ( 
.A(n_1880),
.B(n_1352),
.Y(n_2405)
);

INVxp67_ASAP7_75t_R g2406 ( 
.A(n_1882),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_1983),
.Y(n_2407)
);

CKINVDCx5p33_ASAP7_75t_R g2408 ( 
.A(n_1983),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1920),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_1983),
.Y(n_2410)
);

INVx3_ASAP7_75t_L g2411 ( 
.A(n_1943),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_1983),
.Y(n_2412)
);

CKINVDCx5p33_ASAP7_75t_R g2413 ( 
.A(n_1983),
.Y(n_2413)
);

CKINVDCx5p33_ASAP7_75t_R g2414 ( 
.A(n_1983),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_1920),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1920),
.Y(n_2416)
);

HB1xp67_ASAP7_75t_L g2417 ( 
.A(n_1983),
.Y(n_2417)
);

CKINVDCx16_ASAP7_75t_R g2418 ( 
.A(n_1882),
.Y(n_2418)
);

BUFx3_ASAP7_75t_L g2419 ( 
.A(n_1983),
.Y(n_2419)
);

NAND2xp33_ASAP7_75t_R g2420 ( 
.A(n_1917),
.B(n_1189),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_1983),
.Y(n_2421)
);

CKINVDCx20_ASAP7_75t_R g2422 ( 
.A(n_1935),
.Y(n_2422)
);

INVx3_ASAP7_75t_L g2423 ( 
.A(n_1943),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_R g2424 ( 
.A(n_1880),
.B(n_1676),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_R g2425 ( 
.A(n_1880),
.B(n_1702),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_1983),
.Y(n_2426)
);

CKINVDCx20_ASAP7_75t_R g2427 ( 
.A(n_1935),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_1983),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1999),
.B(n_1083),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_2401),
.Y(n_2430)
);

HB1xp67_ASAP7_75t_L g2431 ( 
.A(n_2139),
.Y(n_2431)
);

BUFx6f_ASAP7_75t_SL g2432 ( 
.A(n_2401),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2223),
.B(n_1190),
.Y(n_2433)
);

CKINVDCx20_ASAP7_75t_R g2434 ( 
.A(n_2122),
.Y(n_2434)
);

INVxp67_ASAP7_75t_SL g2435 ( 
.A(n_2297),
.Y(n_2435)
);

AND2x4_ASAP7_75t_L g2436 ( 
.A(n_2419),
.B(n_1389),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2315),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2233),
.B(n_1191),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2315),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2324),
.Y(n_2440)
);

NOR2xp33_ASAP7_75t_L g2441 ( 
.A(n_2244),
.B(n_1706),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2246),
.B(n_1193),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2202),
.B(n_1206),
.Y(n_2443)
);

NOR2x1_ASAP7_75t_L g2444 ( 
.A(n_2217),
.B(n_1389),
.Y(n_2444)
);

AND2x4_ASAP7_75t_SL g2445 ( 
.A(n_2417),
.B(n_1469),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2132),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_2348),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2232),
.B(n_1207),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2174),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2256),
.Y(n_2450)
);

BUFx3_ASAP7_75t_L g2451 ( 
.A(n_2356),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2178),
.B(n_1211),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2146),
.B(n_1495),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2309),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2177),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2241),
.B(n_1216),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2150),
.B(n_1495),
.Y(n_2457)
);

AOI22xp33_ASAP7_75t_L g2458 ( 
.A1(n_2188),
.A2(n_1552),
.B1(n_1664),
.B2(n_1651),
.Y(n_2458)
);

XNOR2xp5_ASAP7_75t_L g2459 ( 
.A(n_2121),
.B(n_1536),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2183),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2243),
.B(n_1221),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2344),
.B(n_1227),
.Y(n_2462)
);

INVx2_ASAP7_75t_SL g2463 ( 
.A(n_2399),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2115),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_SL g2465 ( 
.A(n_2140),
.B(n_1536),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_L g2466 ( 
.A(n_2181),
.B(n_2295),
.Y(n_2466)
);

BUFx4f_ASAP7_75t_L g2467 ( 
.A(n_2147),
.Y(n_2467)
);

BUFx10_ASAP7_75t_L g2468 ( 
.A(n_2169),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2118),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_2116),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2322),
.B(n_1229),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2156),
.B(n_1550),
.Y(n_2472)
);

AOI22xp33_ASAP7_75t_L g2473 ( 
.A1(n_2188),
.A2(n_1552),
.B1(n_1664),
.B2(n_1651),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2123),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2157),
.B(n_2124),
.Y(n_2475)
);

NOR2xp33_ASAP7_75t_L g2476 ( 
.A(n_2296),
.B(n_1233),
.Y(n_2476)
);

INVx5_ASAP7_75t_L g2477 ( 
.A(n_2154),
.Y(n_2477)
);

INVx3_ASAP7_75t_L g2478 ( 
.A(n_2395),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2141),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2402),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_SL g2481 ( 
.A(n_2170),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_SL g2482 ( 
.A(n_2247),
.B(n_1235),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2409),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2142),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2415),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2416),
.Y(n_2486)
);

NOR2x1p5_ASAP7_75t_L g2487 ( 
.A(n_2162),
.B(n_1236),
.Y(n_2487)
);

NOR2xp33_ASAP7_75t_L g2488 ( 
.A(n_2148),
.B(n_1239),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2313),
.B(n_1550),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_L g2490 ( 
.A(n_2291),
.B(n_2294),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2345),
.B(n_2347),
.Y(n_2491)
);

NOR2x1p5_ASAP7_75t_L g2492 ( 
.A(n_2144),
.B(n_1249),
.Y(n_2492)
);

BUFx2_ASAP7_75t_L g2493 ( 
.A(n_2329),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2334),
.B(n_1621),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_L g2495 ( 
.A(n_2285),
.B(n_1253),
.Y(n_2495)
);

OR2x6_ASAP7_75t_L g2496 ( 
.A(n_2137),
.B(n_1201),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2129),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2350),
.B(n_1255),
.Y(n_2498)
);

OR2x6_ASAP7_75t_L g2499 ( 
.A(n_2128),
.B(n_1418),
.Y(n_2499)
);

AND2x4_ASAP7_75t_L g2500 ( 
.A(n_2397),
.B(n_1621),
.Y(n_2500)
);

NAND3xp33_ASAP7_75t_L g2501 ( 
.A(n_2161),
.B(n_1259),
.C(n_1256),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2318),
.Y(n_2502)
);

INVx4_ASAP7_75t_L g2503 ( 
.A(n_2398),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2214),
.B(n_2206),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2143),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2320),
.Y(n_2506)
);

OR2x6_ASAP7_75t_L g2507 ( 
.A(n_2358),
.B(n_1062),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2250),
.B(n_1262),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2332),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2339),
.Y(n_2510)
);

NAND2xp33_ASAP7_75t_L g2511 ( 
.A(n_2117),
.B(n_1083),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2251),
.B(n_1265),
.Y(n_2512)
);

INVxp67_ASAP7_75t_SL g2513 ( 
.A(n_2307),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2252),
.B(n_1269),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2351),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2187),
.Y(n_2516)
);

INVx4_ASAP7_75t_L g2517 ( 
.A(n_2400),
.Y(n_2517)
);

AND2x4_ASAP7_75t_L g2518 ( 
.A(n_2403),
.B(n_1101),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2190),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2117),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2117),
.Y(n_2521)
);

AOI22xp33_ASAP7_75t_L g2522 ( 
.A1(n_2255),
.A2(n_1432),
.B1(n_1083),
.B2(n_1275),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2267),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_2407),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2326),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2408),
.Y(n_2526)
);

BUFx6f_ASAP7_75t_L g2527 ( 
.A(n_2256),
.Y(n_2527)
);

NAND3xp33_ASAP7_75t_L g2528 ( 
.A(n_2420),
.B(n_1278),
.C(n_1274),
.Y(n_2528)
);

OR2x2_ASAP7_75t_L g2529 ( 
.A(n_2418),
.B(n_1258),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2396),
.B(n_1469),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2256),
.Y(n_2531)
);

INVx3_ASAP7_75t_L g2532 ( 
.A(n_2410),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2259),
.B(n_1279),
.Y(n_2533)
);

INVx2_ASAP7_75t_SL g2534 ( 
.A(n_2412),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2249),
.B(n_1281),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_2165),
.Y(n_2536)
);

BUFx6f_ASAP7_75t_L g2537 ( 
.A(n_2281),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2429),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2413),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2238),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_SL g2541 ( 
.A(n_2261),
.B(n_1282),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_2281),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2414),
.B(n_2421),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2263),
.B(n_2265),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2426),
.B(n_1144),
.Y(n_2545)
);

INVx3_ASAP7_75t_L g2546 ( 
.A(n_2428),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_SL g2547 ( 
.A(n_2268),
.B(n_1284),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_L g2548 ( 
.A(n_2276),
.B(n_1285),
.Y(n_2548)
);

BUFx6f_ASAP7_75t_L g2549 ( 
.A(n_2281),
.Y(n_2549)
);

BUFx6f_ASAP7_75t_L g2550 ( 
.A(n_2292),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2292),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2172),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_L g2553 ( 
.A(n_2280),
.B(n_1287),
.Y(n_2553)
);

HB1xp67_ASAP7_75t_L g2554 ( 
.A(n_2319),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2269),
.B(n_1288),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2292),
.Y(n_2556)
);

OAI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2272),
.A2(n_2274),
.B1(n_2278),
.B2(n_2273),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2310),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2406),
.B(n_1469),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2327),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2275),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2303),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2287),
.B(n_1291),
.Y(n_2563)
);

BUFx4f_ASAP7_75t_L g2564 ( 
.A(n_2293),
.Y(n_2564)
);

INVx2_ASAP7_75t_SL g2565 ( 
.A(n_2131),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2236),
.Y(n_2566)
);

AO22x2_ASAP7_75t_L g2567 ( 
.A1(n_2284),
.A2(n_1344),
.B1(n_1373),
.B2(n_1159),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_L g2568 ( 
.A(n_2288),
.B(n_1292),
.Y(n_2568)
);

BUFx6f_ASAP7_75t_L g2569 ( 
.A(n_2373),
.Y(n_2569)
);

AO22x2_ASAP7_75t_L g2570 ( 
.A1(n_2138),
.A2(n_1705),
.B1(n_1367),
.B2(n_1369),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2316),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2333),
.Y(n_2572)
);

INVx2_ASAP7_75t_SL g2573 ( 
.A(n_2158),
.Y(n_2573)
);

INVx3_ASAP7_75t_L g2574 ( 
.A(n_2211),
.Y(n_2574)
);

NOR2xp33_ASAP7_75t_L g2575 ( 
.A(n_2289),
.B(n_1293),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2151),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2242),
.B(n_1493),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_L g2578 ( 
.A(n_2231),
.B(n_1295),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2235),
.B(n_1296),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2298),
.B(n_1298),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2151),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2185),
.B(n_1493),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2152),
.Y(n_2583)
);

OAI21xp33_ASAP7_75t_SL g2584 ( 
.A1(n_2134),
.A2(n_1459),
.B(n_1313),
.Y(n_2584)
);

NOR2xp33_ASAP7_75t_SL g2585 ( 
.A(n_2149),
.B(n_1300),
.Y(n_2585)
);

AND2x2_ASAP7_75t_L g2586 ( 
.A(n_2325),
.B(n_1493),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_2153),
.B(n_1053),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2175),
.Y(n_2588)
);

NOR2x1p5_ASAP7_75t_L g2589 ( 
.A(n_2130),
.B(n_1305),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2205),
.Y(n_2590)
);

OR2x6_ASAP7_75t_L g2591 ( 
.A(n_2230),
.B(n_1062),
.Y(n_2591)
);

INVx5_ASAP7_75t_L g2592 ( 
.A(n_2205),
.Y(n_2592)
);

AND2x2_ASAP7_75t_SL g2593 ( 
.A(n_2198),
.B(n_1712),
.Y(n_2593)
);

INVx8_ASAP7_75t_L g2594 ( 
.A(n_2155),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2405),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2186),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2235),
.B(n_1306),
.Y(n_2597)
);

INVx2_ASAP7_75t_SL g2598 ( 
.A(n_2133),
.Y(n_2598)
);

AND2x6_ASAP7_75t_L g2599 ( 
.A(n_2404),
.B(n_1166),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2277),
.B(n_1309),
.Y(n_2600)
);

BUFx4f_ASAP7_75t_L g2601 ( 
.A(n_2258),
.Y(n_2601)
);

INVx3_ASAP7_75t_L g2602 ( 
.A(n_2213),
.Y(n_2602)
);

INVx4_ASAP7_75t_SL g2603 ( 
.A(n_2341),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2258),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2300),
.B(n_1311),
.Y(n_2605)
);

INVx5_ASAP7_75t_L g2606 ( 
.A(n_2260),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2330),
.A2(n_2337),
.B1(n_2346),
.B2(n_2340),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2189),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2277),
.B(n_1320),
.Y(n_2609)
);

NAND2xp33_ASAP7_75t_L g2610 ( 
.A(n_2221),
.B(n_1432),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2349),
.B(n_1323),
.Y(n_2611)
);

INVx2_ASAP7_75t_SL g2612 ( 
.A(n_2135),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2304),
.B(n_1326),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2167),
.B(n_1327),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2192),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2203),
.Y(n_2616)
);

CKINVDCx5p33_ASAP7_75t_R g2617 ( 
.A(n_2424),
.Y(n_2617)
);

AOI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2212),
.A2(n_1329),
.B1(n_1330),
.B2(n_1328),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2279),
.B(n_1332),
.Y(n_2619)
);

OR2x6_ASAP7_75t_L g2620 ( 
.A(n_2286),
.B(n_1068),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_2199),
.B(n_1343),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2218),
.Y(n_2622)
);

NAND3xp33_ASAP7_75t_L g2623 ( 
.A(n_2312),
.B(n_1347),
.C(n_1346),
.Y(n_2623)
);

HB1xp67_ASAP7_75t_L g2624 ( 
.A(n_2299),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2260),
.B(n_1350),
.Y(n_2625)
);

BUFx6f_ASAP7_75t_L g2626 ( 
.A(n_2373),
.Y(n_2626)
);

HB1xp67_ASAP7_75t_L g2627 ( 
.A(n_2369),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_L g2628 ( 
.A(n_2200),
.B(n_1359),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2264),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_2425),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2264),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2302),
.Y(n_2632)
);

INVx3_ASAP7_75t_L g2633 ( 
.A(n_2166),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2305),
.B(n_1361),
.Y(n_2634)
);

INVx3_ASAP7_75t_L g2635 ( 
.A(n_2341),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2234),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2308),
.B(n_1362),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2119),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_L g2639 ( 
.A(n_2168),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2311),
.B(n_1374),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2314),
.B(n_1375),
.Y(n_2641)
);

BUFx6f_ASAP7_75t_L g2642 ( 
.A(n_2168),
.Y(n_2642)
);

INVx6_ASAP7_75t_L g2643 ( 
.A(n_2341),
.Y(n_2643)
);

INVx2_ASAP7_75t_SL g2644 ( 
.A(n_2136),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2306),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_L g2646 ( 
.A(n_2208),
.B(n_1376),
.Y(n_2646)
);

AND2x4_ASAP7_75t_L g2647 ( 
.A(n_2120),
.B(n_1072),
.Y(n_2647)
);

AND2x4_ASAP7_75t_L g2648 ( 
.A(n_2125),
.B(n_1102),
.Y(n_2648)
);

BUFx3_ASAP7_75t_L g2649 ( 
.A(n_2357),
.Y(n_2649)
);

INVx2_ASAP7_75t_SL g2650 ( 
.A(n_2191),
.Y(n_2650)
);

NAND3xp33_ASAP7_75t_SL g2651 ( 
.A(n_2215),
.B(n_1385),
.C(n_1381),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2119),
.Y(n_2652)
);

BUFx6f_ASAP7_75t_L g2653 ( 
.A(n_2361),
.Y(n_2653)
);

AND2x6_ASAP7_75t_L g2654 ( 
.A(n_2411),
.B(n_1166),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2194),
.B(n_2180),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2411),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2126),
.B(n_1117),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2423),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2204),
.B(n_1393),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2423),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2370),
.Y(n_2661)
);

OR2x2_ASAP7_75t_L g2662 ( 
.A(n_2173),
.B(n_1511),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2317),
.B(n_1394),
.Y(n_2663)
);

AND2x4_ASAP7_75t_L g2664 ( 
.A(n_2127),
.B(n_1176),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2321),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2145),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2323),
.B(n_1398),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2328),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2331),
.Y(n_2669)
);

OR2x6_ASAP7_75t_L g2670 ( 
.A(n_2195),
.B(n_1068),
.Y(n_2670)
);

BUFx3_ASAP7_75t_L g2671 ( 
.A(n_2367),
.Y(n_2671)
);

OR2x2_ASAP7_75t_L g2672 ( 
.A(n_2179),
.B(n_1533),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2176),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2224),
.B(n_2335),
.Y(n_2674)
);

INVx2_ASAP7_75t_SL g2675 ( 
.A(n_2197),
.Y(n_2675)
);

INVx3_ASAP7_75t_L g2676 ( 
.A(n_2237),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2222),
.Y(n_2677)
);

BUFx3_ASAP7_75t_L g2678 ( 
.A(n_2159),
.Y(n_2678)
);

AND3x4_ASAP7_75t_L g2679 ( 
.A(n_2422),
.B(n_1126),
.C(n_1111),
.Y(n_2679)
);

INVx3_ASAP7_75t_L g2680 ( 
.A(n_2239),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2336),
.Y(n_2681)
);

INVxp67_ASAP7_75t_SL g2682 ( 
.A(n_2248),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2338),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2342),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2343),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2184),
.B(n_1399),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2163),
.B(n_1254),
.Y(n_2687)
);

INVx4_ASAP7_75t_L g2688 ( 
.A(n_2363),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2282),
.B(n_1400),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2193),
.Y(n_2690)
);

BUFx10_ASAP7_75t_L g2691 ( 
.A(n_2352),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_2427),
.B(n_1263),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2222),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2201),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2225),
.B(n_1401),
.Y(n_2695)
);

BUFx4f_ASAP7_75t_L g2696 ( 
.A(n_2207),
.Y(n_2696)
);

INVx3_ASAP7_75t_L g2697 ( 
.A(n_2366),
.Y(n_2697)
);

BUFx6f_ASAP7_75t_L g2698 ( 
.A(n_2368),
.Y(n_2698)
);

BUFx3_ASAP7_75t_L g2699 ( 
.A(n_2371),
.Y(n_2699)
);

INVx6_ASAP7_75t_L g2700 ( 
.A(n_2386),
.Y(n_2700)
);

INVx3_ASAP7_75t_L g2701 ( 
.A(n_2374),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2228),
.B(n_1402),
.Y(n_2702)
);

OR2x2_ASAP7_75t_L g2703 ( 
.A(n_2171),
.B(n_1543),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2209),
.Y(n_2704)
);

INVx1_ASAP7_75t_SL g2705 ( 
.A(n_2375),
.Y(n_2705)
);

AOI22xp5_ASAP7_75t_L g2706 ( 
.A1(n_2229),
.A2(n_1404),
.B1(n_1408),
.B2(n_1403),
.Y(n_2706)
);

INVx2_ASAP7_75t_SL g2707 ( 
.A(n_2227),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2219),
.B(n_1409),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2226),
.Y(n_2709)
);

BUFx2_ASAP7_75t_L g2710 ( 
.A(n_2290),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2240),
.B(n_1412),
.Y(n_2711)
);

INVx3_ASAP7_75t_L g2712 ( 
.A(n_2379),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_SL g2713 ( 
.A(n_2216),
.B(n_1414),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2245),
.Y(n_2714)
);

BUFx4f_ASAP7_75t_L g2715 ( 
.A(n_2253),
.Y(n_2715)
);

BUFx3_ASAP7_75t_L g2716 ( 
.A(n_2380),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2257),
.B(n_1415),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2266),
.Y(n_2718)
);

BUFx6f_ASAP7_75t_L g2719 ( 
.A(n_2383),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2196),
.B(n_1427),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2254),
.Y(n_2721)
);

AND2x6_ASAP7_75t_L g2722 ( 
.A(n_2270),
.B(n_1166),
.Y(n_2722)
);

INVx3_ASAP7_75t_L g2723 ( 
.A(n_2384),
.Y(n_2723)
);

INVxp67_ASAP7_75t_SL g2724 ( 
.A(n_2365),
.Y(n_2724)
);

AND2x4_ASAP7_75t_L g2725 ( 
.A(n_2160),
.B(n_1466),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2182),
.B(n_1430),
.Y(n_2726)
);

BUFx6f_ASAP7_75t_L g2727 ( 
.A(n_2385),
.Y(n_2727)
);

BUFx6f_ASAP7_75t_L g2728 ( 
.A(n_2387),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2271),
.Y(n_2729)
);

NOR2x1p5_ASAP7_75t_L g2730 ( 
.A(n_2164),
.B(n_1431),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2283),
.B(n_1434),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_2220),
.A2(n_1432),
.B1(n_1437),
.B2(n_1436),
.Y(n_2732)
);

BUFx4f_ASAP7_75t_L g2733 ( 
.A(n_2301),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2353),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_SL g2735 ( 
.A(n_2262),
.B(n_1439),
.Y(n_2735)
);

BUFx3_ASAP7_75t_L g2736 ( 
.A(n_2388),
.Y(n_2736)
);

INVx4_ASAP7_75t_L g2737 ( 
.A(n_2392),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2210),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2377),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2362),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2393),
.B(n_1440),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_SL g2742 ( 
.A(n_2394),
.B(n_1444),
.Y(n_2742)
);

OAI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2381),
.A2(n_1448),
.B1(n_1452),
.B2(n_1446),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2364),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2391),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2364),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2376),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2376),
.Y(n_2748)
);

AOI22xp5_ASAP7_75t_SL g2749 ( 
.A1(n_2378),
.A2(n_1460),
.B1(n_1461),
.B2(n_1454),
.Y(n_2749)
);

BUFx6f_ASAP7_75t_L g2750 ( 
.A(n_2382),
.Y(n_2750)
);

CKINVDCx5p33_ASAP7_75t_R g2751 ( 
.A(n_2378),
.Y(n_2751)
);

AO22x2_ASAP7_75t_L g2752 ( 
.A1(n_2354),
.A2(n_1672),
.B1(n_1698),
.B2(n_1516),
.Y(n_2752)
);

AND2x2_ASAP7_75t_SL g2753 ( 
.A(n_2382),
.B(n_1429),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2382),
.B(n_1471),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2355),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2359),
.B(n_1478),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2360),
.B(n_1481),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_2390),
.B(n_1065),
.Y(n_2758)
);

INVx4_ASAP7_75t_L g2759 ( 
.A(n_2372),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2389),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2309),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2139),
.B(n_1487),
.Y(n_2762)
);

INVx3_ASAP7_75t_L g2763 ( 
.A(n_2401),
.Y(n_2763)
);

BUFx10_ASAP7_75t_L g2764 ( 
.A(n_2169),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2139),
.B(n_1490),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2315),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2154),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2401),
.Y(n_2768)
);

NOR2xp33_ASAP7_75t_L g2769 ( 
.A(n_2244),
.B(n_1496),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_SL g2770 ( 
.A(n_2315),
.B(n_1497),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2315),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2315),
.Y(n_2772)
);

NAND2xp33_ASAP7_75t_L g2773 ( 
.A(n_2117),
.B(n_1432),
.Y(n_2773)
);

AND2x6_ASAP7_75t_L g2774 ( 
.A(n_2223),
.B(n_1166),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2223),
.B(n_1502),
.Y(n_2775)
);

OR2x6_ASAP7_75t_L g2776 ( 
.A(n_2399),
.B(n_1111),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2315),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2315),
.Y(n_2778)
);

OR2x6_ASAP7_75t_L g2779 ( 
.A(n_2399),
.B(n_1126),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2315),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2223),
.B(n_1503),
.Y(n_2781)
);

INVx3_ASAP7_75t_L g2782 ( 
.A(n_2401),
.Y(n_2782)
);

BUFx4_ASAP7_75t_L g2783 ( 
.A(n_2154),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2309),
.Y(n_2784)
);

NAND2xp33_ASAP7_75t_L g2785 ( 
.A(n_2117),
.B(n_1432),
.Y(n_2785)
);

AOI22xp33_ASAP7_75t_L g2786 ( 
.A1(n_2188),
.A2(n_1432),
.B1(n_1519),
.B2(n_1507),
.Y(n_2786)
);

INVx3_ASAP7_75t_L g2787 ( 
.A(n_2401),
.Y(n_2787)
);

AOI22xp33_ASAP7_75t_L g2788 ( 
.A1(n_2188),
.A2(n_1432),
.B1(n_1527),
.B2(n_1520),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2244),
.B(n_1528),
.Y(n_2789)
);

BUFx10_ASAP7_75t_L g2790 ( 
.A(n_2169),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2315),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2315),
.B(n_1542),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_L g2793 ( 
.A(n_2244),
.B(n_1544),
.Y(n_2793)
);

NAND3xp33_ASAP7_75t_L g2794 ( 
.A(n_2244),
.B(n_1561),
.C(n_1560),
.Y(n_2794)
);

INVx4_ASAP7_75t_SL g2795 ( 
.A(n_2139),
.Y(n_2795)
);

NOR2xp33_ASAP7_75t_L g2796 ( 
.A(n_2244),
.B(n_1568),
.Y(n_2796)
);

INVx3_ASAP7_75t_L g2797 ( 
.A(n_2401),
.Y(n_2797)
);

OR2x6_ASAP7_75t_L g2798 ( 
.A(n_2399),
.B(n_1273),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2309),
.Y(n_2799)
);

BUFx3_ASAP7_75t_L g2800 ( 
.A(n_2356),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2223),
.B(n_1570),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2309),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2419),
.B(n_1075),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2309),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2154),
.Y(n_2805)
);

AND2x2_ASAP7_75t_SL g2806 ( 
.A(n_2322),
.B(n_1433),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2315),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2309),
.Y(n_2808)
);

INVx2_ASAP7_75t_SL g2809 ( 
.A(n_2401),
.Y(n_2809)
);

BUFx6f_ASAP7_75t_L g2810 ( 
.A(n_2401),
.Y(n_2810)
);

INVxp33_ASAP7_75t_L g2811 ( 
.A(n_2313),
.Y(n_2811)
);

OR2x2_ASAP7_75t_L g2812 ( 
.A(n_2322),
.B(n_1571),
.Y(n_2812)
);

AO22x2_ASAP7_75t_L g2813 ( 
.A1(n_2146),
.A2(n_1100),
.B1(n_1115),
.B2(n_1098),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2315),
.Y(n_2814)
);

INVx5_ASAP7_75t_L g2815 ( 
.A(n_2401),
.Y(n_2815)
);

BUFx6f_ASAP7_75t_L g2816 ( 
.A(n_2401),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2315),
.Y(n_2817)
);

OR2x2_ASAP7_75t_L g2818 ( 
.A(n_2322),
.B(n_1572),
.Y(n_2818)
);

AO22x2_ASAP7_75t_L g2819 ( 
.A1(n_2146),
.A2(n_1137),
.B1(n_1146),
.B2(n_1124),
.Y(n_2819)
);

OR2x2_ASAP7_75t_L g2820 ( 
.A(n_2322),
.B(n_1573),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2139),
.B(n_1574),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2223),
.B(n_1575),
.Y(n_2822)
);

INVx1_ASAP7_75t_SL g2823 ( 
.A(n_2139),
.Y(n_2823)
);

AND2x6_ASAP7_75t_L g2824 ( 
.A(n_2223),
.B(n_1225),
.Y(n_2824)
);

AOI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2244),
.A2(n_1578),
.B1(n_1579),
.B2(n_1576),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_L g2826 ( 
.A(n_2823),
.B(n_1584),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2544),
.B(n_1591),
.Y(n_2827)
);

AO22x2_ASAP7_75t_L g2828 ( 
.A1(n_2679),
.A2(n_1443),
.B1(n_1451),
.B2(n_1438),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2431),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2441),
.B(n_1596),
.Y(n_2830)
);

NAND2x1p5_ASAP7_75t_L g2831 ( 
.A(n_2815),
.B(n_1225),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2446),
.Y(n_2832)
);

AO22x2_ASAP7_75t_L g2833 ( 
.A1(n_2557),
.A2(n_1456),
.B1(n_1458),
.B2(n_1453),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2449),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2455),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2437),
.B(n_1156),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2460),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2497),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2479),
.Y(n_2839)
);

OR2x2_ASAP7_75t_SL g2840 ( 
.A(n_2783),
.B(n_1165),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2439),
.B(n_1605),
.Y(n_2841)
);

NAND3x1_ASAP7_75t_L g2842 ( 
.A(n_2607),
.B(n_1177),
.C(n_1173),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2766),
.B(n_1607),
.Y(n_2843)
);

AND2x4_ASAP7_75t_L g2844 ( 
.A(n_2771),
.B(n_1178),
.Y(n_2844)
);

AOI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2806),
.A2(n_1611),
.B1(n_1612),
.B2(n_1608),
.Y(n_2845)
);

INVxp67_ASAP7_75t_L g2846 ( 
.A(n_2465),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2535),
.A2(n_1619),
.B1(n_1625),
.B2(n_1613),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2772),
.B(n_1631),
.Y(n_2848)
);

BUFx8_ASAP7_75t_L g2849 ( 
.A(n_2481),
.Y(n_2849)
);

AO22x2_ASAP7_75t_L g2850 ( 
.A1(n_2795),
.A2(n_1477),
.B1(n_1479),
.B2(n_1470),
.Y(n_2850)
);

BUFx3_ASAP7_75t_L g2851 ( 
.A(n_2430),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2440),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2464),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2469),
.Y(n_2854)
);

AND2x4_ASAP7_75t_L g2855 ( 
.A(n_2777),
.B(n_1181),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2474),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2480),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2484),
.Y(n_2858)
);

BUFx2_ASAP7_75t_L g2859 ( 
.A(n_2434),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2505),
.Y(n_2860)
);

AND2x4_ASAP7_75t_L g2861 ( 
.A(n_2778),
.B(n_2780),
.Y(n_2861)
);

OAI221xp5_ASAP7_75t_L g2862 ( 
.A1(n_2504),
.A2(n_1637),
.B1(n_1641),
.B2(n_1636),
.C(n_1634),
.Y(n_2862)
);

AND2x4_ASAP7_75t_L g2863 ( 
.A(n_2791),
.B(n_1196),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2583),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2807),
.B(n_1643),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2483),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2485),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2762),
.B(n_1646),
.Y(n_2868)
);

OR2x2_ASAP7_75t_SL g2869 ( 
.A(n_2624),
.B(n_1197),
.Y(n_2869)
);

OR2x2_ASAP7_75t_SL g2870 ( 
.A(n_2554),
.B(n_1198),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_SL g2871 ( 
.A(n_2767),
.B(n_1650),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2486),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2814),
.B(n_1652),
.Y(n_2873)
);

AO22x2_ASAP7_75t_L g2874 ( 
.A1(n_2795),
.A2(n_1486),
.B1(n_1489),
.B2(n_1480),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2817),
.B(n_1653),
.Y(n_2875)
);

A2O1A1Ixp33_ASAP7_75t_L g2876 ( 
.A1(n_2525),
.A2(n_1512),
.B(n_1513),
.C(n_1504),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2588),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2765),
.B(n_1655),
.Y(n_2878)
);

CKINVDCx20_ASAP7_75t_R g2879 ( 
.A(n_2594),
.Y(n_2879)
);

BUFx2_ASAP7_75t_L g2880 ( 
.A(n_2513),
.Y(n_2880)
);

AND2x4_ASAP7_75t_L g2881 ( 
.A(n_2523),
.B(n_1208),
.Y(n_2881)
);

INVxp67_ASAP7_75t_L g2882 ( 
.A(n_2529),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2596),
.Y(n_2883)
);

AOI22xp33_ASAP7_75t_L g2884 ( 
.A1(n_2593),
.A2(n_1659),
.B1(n_1665),
.B2(n_1658),
.Y(n_2884)
);

NAND2x1p5_ASAP7_75t_L g2885 ( 
.A(n_2815),
.B(n_2430),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2770),
.B(n_1213),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_SL g2887 ( 
.A(n_2585),
.B(n_1669),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2821),
.B(n_1677),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2502),
.Y(n_2889)
);

AO22x2_ASAP7_75t_L g2890 ( 
.A1(n_2489),
.A2(n_1521),
.B1(n_1524),
.B2(n_1517),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2506),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2608),
.Y(n_2892)
);

CKINVDCx5p33_ASAP7_75t_R g2893 ( 
.A(n_2805),
.Y(n_2893)
);

AO22x2_ASAP7_75t_L g2894 ( 
.A1(n_2494),
.A2(n_2813),
.B1(n_2819),
.B2(n_2540),
.Y(n_2894)
);

INVxp67_ASAP7_75t_L g2895 ( 
.A(n_2611),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2453),
.B(n_2457),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2615),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2509),
.Y(n_2898)
);

AO22x2_ASAP7_75t_L g2899 ( 
.A1(n_2813),
.A2(n_1526),
.B1(n_1538),
.B2(n_1525),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_SL g2900 ( 
.A(n_2753),
.B(n_2749),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2510),
.Y(n_2901)
);

AO22x2_ASAP7_75t_L g2902 ( 
.A1(n_2819),
.A2(n_1541),
.B1(n_1545),
.B2(n_1540),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2558),
.B(n_1681),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2516),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2560),
.B(n_2433),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2519),
.Y(n_2906)
);

INVx1_ASAP7_75t_SL g2907 ( 
.A(n_2451),
.Y(n_2907)
);

NAND2xp33_ASAP7_75t_L g2908 ( 
.A(n_2750),
.B(n_1690),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2515),
.Y(n_2909)
);

NAND2x1p5_ASAP7_75t_L g2910 ( 
.A(n_2768),
.B(n_1225),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2438),
.B(n_1687),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2475),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2571),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2720),
.B(n_2769),
.Y(n_2914)
);

INVx3_ASAP7_75t_L g2915 ( 
.A(n_2569),
.Y(n_2915)
);

OAI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2458),
.A2(n_1692),
.B1(n_1694),
.B2(n_1689),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2616),
.Y(n_2917)
);

INVxp67_ASAP7_75t_L g2918 ( 
.A(n_2491),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2572),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2621),
.B(n_1696),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_L g2921 ( 
.A(n_2628),
.B(n_1703),
.Y(n_2921)
);

HB1xp67_ASAP7_75t_L g2922 ( 
.A(n_2649),
.Y(n_2922)
);

AO22x2_ASAP7_75t_L g2923 ( 
.A1(n_2677),
.A2(n_1556),
.B1(n_1559),
.B2(n_1547),
.Y(n_2923)
);

AO22x2_ASAP7_75t_L g2924 ( 
.A1(n_2693),
.A2(n_1564),
.B1(n_1565),
.B2(n_1562),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2622),
.Y(n_2925)
);

INVx2_ASAP7_75t_SL g2926 ( 
.A(n_2594),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2632),
.Y(n_2927)
);

OA22x2_ASAP7_75t_L g2928 ( 
.A1(n_2459),
.A2(n_1707),
.B1(n_1709),
.B2(n_1704),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2562),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2758),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2740),
.Y(n_2931)
);

O2A1O1Ixp33_ASAP7_75t_L g2932 ( 
.A1(n_2584),
.A2(n_1587),
.B(n_1592),
.C(n_1577),
.Y(n_2932)
);

INVxp67_ASAP7_75t_L g2933 ( 
.A(n_2686),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2625),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2636),
.Y(n_2935)
);

INVxp67_ASAP7_75t_L g2936 ( 
.A(n_2812),
.Y(n_2936)
);

A2O1A1Ixp33_ASAP7_75t_L g2937 ( 
.A1(n_2538),
.A2(n_1595),
.B(n_1610),
.C(n_1594),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2754),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2775),
.B(n_1710),
.Y(n_2939)
);

AOI22xp33_ASAP7_75t_L g2940 ( 
.A1(n_2662),
.A2(n_1716),
.B1(n_1718),
.B2(n_1711),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2756),
.Y(n_2941)
);

NAND2x1p5_ASAP7_75t_L g2942 ( 
.A(n_2768),
.B(n_1225),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2708),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2711),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2717),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2781),
.B(n_1722),
.Y(n_2946)
);

NAND2x1p5_ASAP7_75t_L g2947 ( 
.A(n_2810),
.B(n_1230),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2731),
.Y(n_2948)
);

AND2x4_ASAP7_75t_L g2949 ( 
.A(n_2792),
.B(n_1220),
.Y(n_2949)
);

INVxp67_ASAP7_75t_L g2950 ( 
.A(n_2818),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2530),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2660),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2452),
.Y(n_2953)
);

HB1xp67_ASAP7_75t_L g2954 ( 
.A(n_2671),
.Y(n_2954)
);

AND2x4_ASAP7_75t_L g2955 ( 
.A(n_2574),
.B(n_1238),
.Y(n_2955)
);

AND2x4_ASAP7_75t_L g2956 ( 
.A(n_2602),
.B(n_1241),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2690),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2666),
.Y(n_2958)
);

INVxp67_ASAP7_75t_L g2959 ( 
.A(n_2820),
.Y(n_2959)
);

CKINVDCx14_ASAP7_75t_R g2960 ( 
.A(n_2477),
.Y(n_2960)
);

AO22x2_ASAP7_75t_L g2961 ( 
.A1(n_2707),
.A2(n_1627),
.B1(n_1639),
.B2(n_1620),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2694),
.Y(n_2962)
);

A2O1A1Ixp33_ASAP7_75t_L g2963 ( 
.A1(n_2473),
.A2(n_2661),
.B(n_2645),
.C(n_2488),
.Y(n_2963)
);

AO22x2_ASAP7_75t_L g2964 ( 
.A1(n_2672),
.A2(n_1649),
.B1(n_1657),
.B2(n_1642),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2704),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2709),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2638),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2718),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2652),
.Y(n_2969)
);

A2O1A1Ixp33_ASAP7_75t_L g2970 ( 
.A1(n_2522),
.A2(n_1680),
.B(n_1691),
.C(n_1661),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2729),
.Y(n_2971)
);

BUFx2_ASAP7_75t_L g2972 ( 
.A(n_2800),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2801),
.B(n_1723),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2822),
.B(n_1727),
.Y(n_2974)
);

CKINVDCx5p33_ASAP7_75t_R g2975 ( 
.A(n_2432),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2789),
.B(n_1044),
.Y(n_2976)
);

BUFx2_ASAP7_75t_L g2977 ( 
.A(n_2435),
.Y(n_2977)
);

INVx2_ASAP7_75t_SL g2978 ( 
.A(n_2810),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2745),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2442),
.B(n_1693),
.Y(n_2980)
);

AND2x4_ASAP7_75t_L g2981 ( 
.A(n_2592),
.B(n_1257),
.Y(n_2981)
);

BUFx8_ASAP7_75t_L g2982 ( 
.A(n_2526),
.Y(n_2982)
);

O2A1O1Ixp33_ASAP7_75t_L g2983 ( 
.A1(n_2462),
.A2(n_1700),
.B(n_1720),
.C(n_1699),
.Y(n_2983)
);

BUFx2_ASAP7_75t_L g2984 ( 
.A(n_2776),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2576),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2656),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2793),
.B(n_1046),
.Y(n_2987)
);

CKINVDCx20_ASAP7_75t_R g2988 ( 
.A(n_2477),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2658),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2581),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2590),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2604),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2629),
.Y(n_2993)
);

BUFx2_ASAP7_75t_L g2994 ( 
.A(n_2776),
.Y(n_2994)
);

AO22x2_ASAP7_75t_L g2995 ( 
.A1(n_2650),
.A2(n_1294),
.B1(n_1297),
.B2(n_1260),
.Y(n_2995)
);

BUFx6f_ASAP7_75t_L g2996 ( 
.A(n_2750),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2631),
.Y(n_2997)
);

OR2x2_ASAP7_75t_L g2998 ( 
.A(n_2472),
.B(n_1070),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2796),
.B(n_1082),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2454),
.Y(n_3000)
);

AOI211xp5_ASAP7_75t_L g3001 ( 
.A1(n_2811),
.A2(n_1314),
.B(n_1317),
.C(n_1302),
.Y(n_3001)
);

OAI22xp5_ASAP7_75t_L g3002 ( 
.A1(n_2490),
.A2(n_1091),
.B1(n_1096),
.B2(n_1095),
.Y(n_3002)
);

OR2x2_ASAP7_75t_SL g3003 ( 
.A(n_2627),
.B(n_1318),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2761),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2784),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2443),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2739),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2799),
.Y(n_3008)
);

INVx2_ASAP7_75t_SL g3009 ( 
.A(n_2816),
.Y(n_3009)
);

AND3x4_ASAP7_75t_L g3010 ( 
.A(n_2444),
.B(n_1340),
.C(n_1273),
.Y(n_3010)
);

OAI221xp5_ASAP7_75t_L g3011 ( 
.A1(n_2703),
.A2(n_1104),
.B1(n_1132),
.B2(n_1118),
.C(n_1099),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2646),
.B(n_1145),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2448),
.B(n_2659),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2802),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2735),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2561),
.Y(n_3016)
);

AOI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_2548),
.A2(n_1158),
.B1(n_1160),
.B2(n_1152),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2786),
.B(n_1163),
.Y(n_3018)
);

A2O1A1Ixp33_ASAP7_75t_L g3019 ( 
.A1(n_2757),
.A2(n_1324),
.B(n_1337),
.C(n_1335),
.Y(n_3019)
);

INVxp67_ASAP7_75t_L g3020 ( 
.A(n_2493),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2752),
.Y(n_3021)
);

AND2x4_ASAP7_75t_L g3022 ( 
.A(n_2592),
.B(n_2606),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2788),
.B(n_1169),
.Y(n_3023)
);

AO22x2_ASAP7_75t_L g3024 ( 
.A1(n_2570),
.A2(n_1354),
.B1(n_1358),
.B2(n_1339),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2825),
.B(n_2456),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2553),
.B(n_1185),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2734),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2555),
.B(n_1195),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2724),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2804),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2808),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2450),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2691),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2450),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2665),
.Y(n_3035)
);

AOI22xp33_ASAP7_75t_L g3036 ( 
.A1(n_2655),
.A2(n_1202),
.B1(n_1214),
.B2(n_1204),
.Y(n_3036)
);

INVx1_ASAP7_75t_SL g3037 ( 
.A(n_2705),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2668),
.Y(n_3038)
);

AND2x4_ASAP7_75t_L g3039 ( 
.A(n_2606),
.B(n_1372),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2669),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_SL g3041 ( 
.A(n_2569),
.B(n_1695),
.Y(n_3041)
);

AO22x2_ASAP7_75t_L g3042 ( 
.A1(n_2500),
.A2(n_1397),
.B1(n_1416),
.B2(n_1387),
.Y(n_3042)
);

AND2x2_ASAP7_75t_L g3043 ( 
.A(n_2568),
.B(n_1215),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_2468),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2575),
.B(n_1224),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2681),
.Y(n_3046)
);

INVx2_ASAP7_75t_SL g3047 ( 
.A(n_2816),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_2578),
.B(n_2577),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2683),
.Y(n_3049)
);

NOR2xp67_ASAP7_75t_L g3050 ( 
.A(n_2503),
.B(n_0),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2684),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2527),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2685),
.Y(n_3053)
);

NAND2x1p5_ASAP7_75t_L g3054 ( 
.A(n_2626),
.B(n_1230),
.Y(n_3054)
);

NAND2x1p5_ASAP7_75t_L g3055 ( 
.A(n_2626),
.B(n_1230),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2614),
.B(n_1232),
.Y(n_3056)
);

AND2x4_ASAP7_75t_L g3057 ( 
.A(n_2699),
.B(n_1428),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2591),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2591),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2586),
.B(n_1237),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2620),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2620),
.Y(n_3062)
);

AND2x4_ASAP7_75t_L g3063 ( 
.A(n_2716),
.B(n_1445),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2670),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_SL g3065 ( 
.A(n_2467),
.B(n_2743),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2670),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2498),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2527),
.Y(n_3068)
);

INVxp67_ASAP7_75t_L g3069 ( 
.A(n_2741),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2537),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2537),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_2471),
.B(n_1240),
.Y(n_3072)
);

BUFx6f_ASAP7_75t_L g3073 ( 
.A(n_2542),
.Y(n_3073)
);

NAND2x1p5_ASAP7_75t_L g3074 ( 
.A(n_2517),
.B(n_1230),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2573),
.B(n_2675),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2508),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2512),
.Y(n_3077)
);

OR2x2_ASAP7_75t_SL g3078 ( 
.A(n_2651),
.B(n_1678),
.Y(n_3078)
);

AND2x4_ASAP7_75t_L g3079 ( 
.A(n_2736),
.B(n_1447),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2514),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2618),
.B(n_1244),
.Y(n_3081)
);

BUFx3_ASAP7_75t_L g3082 ( 
.A(n_2653),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2542),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2533),
.Y(n_3084)
);

BUFx3_ASAP7_75t_L g3085 ( 
.A(n_2653),
.Y(n_3085)
);

AO22x2_ASAP7_75t_L g3086 ( 
.A1(n_2692),
.A2(n_1474),
.B1(n_1483),
.B2(n_1464),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2563),
.Y(n_3087)
);

NAND2xp33_ASAP7_75t_L g3088 ( 
.A(n_2654),
.B(n_1199),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2803),
.Y(n_3089)
);

CKINVDCx5p33_ASAP7_75t_R g3090 ( 
.A(n_2764),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2549),
.Y(n_3091)
);

NAND2x1p5_ASAP7_75t_L g3092 ( 
.A(n_2698),
.B(n_1355),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2755),
.Y(n_3093)
);

BUFx8_ASAP7_75t_L g3094 ( 
.A(n_2543),
.Y(n_3094)
);

NAND2x1p5_ASAP7_75t_L g3095 ( 
.A(n_2698),
.B(n_1355),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2760),
.Y(n_3096)
);

NAND3x1_ASAP7_75t_L g3097 ( 
.A(n_2674),
.B(n_1715),
.C(n_1488),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2482),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2541),
.Y(n_3099)
);

AO22x2_ASAP7_75t_L g3100 ( 
.A1(n_2566),
.A2(n_2565),
.B1(n_2518),
.B2(n_2545),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2476),
.B(n_1250),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2466),
.B(n_1267),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2634),
.B(n_1268),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2547),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2637),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2640),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2641),
.B(n_1271),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2663),
.Y(n_3108)
);

CKINVDCx5p33_ASAP7_75t_R g3109 ( 
.A(n_2790),
.Y(n_3109)
);

BUFx2_ASAP7_75t_L g3110 ( 
.A(n_2779),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2667),
.Y(n_3111)
);

AOI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_2726),
.A2(n_1286),
.B1(n_1303),
.B2(n_1289),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2579),
.B(n_1307),
.Y(n_3113)
);

NAND2x1p5_ASAP7_75t_L g3114 ( 
.A(n_2719),
.B(n_1355),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2597),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2549),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2550),
.Y(n_3117)
);

AO22x2_ASAP7_75t_L g3118 ( 
.A1(n_2598),
.A2(n_1499),
.B1(n_1506),
.B2(n_1485),
.Y(n_3118)
);

INVxp67_ASAP7_75t_L g3119 ( 
.A(n_2779),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2550),
.Y(n_3120)
);

AND2x4_ASAP7_75t_L g3121 ( 
.A(n_2688),
.B(n_1510),
.Y(n_3121)
);

OAI22xp5_ASAP7_75t_SL g3122 ( 
.A1(n_2738),
.A2(n_1721),
.B1(n_1725),
.B2(n_1708),
.Y(n_3122)
);

AO22x2_ASAP7_75t_L g3123 ( 
.A1(n_2612),
.A2(n_1529),
.B1(n_1532),
.B2(n_1514),
.Y(n_3123)
);

CKINVDCx5p33_ASAP7_75t_R g3124 ( 
.A(n_2595),
.Y(n_3124)
);

CKINVDCx5p33_ASAP7_75t_R g3125 ( 
.A(n_2617),
.Y(n_3125)
);

NAND2x1p5_ASAP7_75t_L g3126 ( 
.A(n_2719),
.B(n_1355),
.Y(n_3126)
);

AOI22xp5_ASAP7_75t_L g3127 ( 
.A1(n_2580),
.A2(n_1310),
.B1(n_1321),
.B2(n_1316),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_2706),
.B(n_1322),
.Y(n_3128)
);

A2O1A1Ixp33_ASAP7_75t_L g3129 ( 
.A1(n_2619),
.A2(n_1557),
.B(n_1581),
.C(n_1554),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_2582),
.B(n_1325),
.Y(n_3130)
);

A2O1A1Ixp33_ASAP7_75t_L g3131 ( 
.A1(n_2794),
.A2(n_1597),
.B(n_1603),
.C(n_1582),
.Y(n_3131)
);

BUFx8_ASAP7_75t_L g3132 ( 
.A(n_2534),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2600),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2609),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2751),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2499),
.Y(n_3136)
);

AO22x2_ASAP7_75t_L g3137 ( 
.A1(n_2644),
.A2(n_1668),
.B1(n_1670),
.B2(n_1662),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_SL g3138 ( 
.A(n_2678),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2499),
.Y(n_3139)
);

INVx3_ASAP7_75t_L g3140 ( 
.A(n_2727),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2689),
.B(n_1333),
.Y(n_3141)
);

INVxp67_ASAP7_75t_L g3142 ( 
.A(n_2798),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2507),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2507),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2682),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2559),
.B(n_1334),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2747),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2531),
.Y(n_3148)
);

CKINVDCx5p33_ASAP7_75t_R g3149 ( 
.A(n_2630),
.Y(n_3149)
);

NOR2xp33_ASAP7_75t_L g3150 ( 
.A(n_2495),
.B(n_1336),
.Y(n_3150)
);

AND2x4_ASAP7_75t_L g3151 ( 
.A(n_2737),
.B(n_2496),
.Y(n_3151)
);

HB1xp67_ASAP7_75t_L g3152 ( 
.A(n_2463),
.Y(n_3152)
);

NOR3xp33_ASAP7_75t_L g3153 ( 
.A(n_2501),
.B(n_1675),
.C(n_1345),
.Y(n_3153)
);

AOI22xp33_ASAP7_75t_L g3154 ( 
.A1(n_2725),
.A2(n_1338),
.B1(n_1364),
.B2(n_1353),
.Y(n_3154)
);

CKINVDCx20_ASAP7_75t_R g3155 ( 
.A(n_2552),
.Y(n_3155)
);

AO22x2_ASAP7_75t_L g3156 ( 
.A1(n_2436),
.A2(n_1341),
.B1(n_1349),
.B2(n_1340),
.Y(n_3156)
);

BUFx6f_ASAP7_75t_L g3157 ( 
.A(n_2654),
.Y(n_3157)
);

BUFx8_ASAP7_75t_L g3158 ( 
.A(n_2727),
.Y(n_3158)
);

NOR2xp33_ASAP7_75t_L g3159 ( 
.A(n_2605),
.B(n_2613),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2732),
.B(n_1365),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2551),
.Y(n_3161)
);

AND2x4_ASAP7_75t_L g3162 ( 
.A(n_2496),
.B(n_1341),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2567),
.B(n_1368),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2714),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2623),
.B(n_2774),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_SL g3166 ( 
.A(n_2536),
.B(n_1371),
.Y(n_3166)
);

INVxp67_ASAP7_75t_L g3167 ( 
.A(n_2798),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2721),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2556),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2696),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2715),
.Y(n_3171)
);

OR2x2_ASAP7_75t_L g3172 ( 
.A(n_2710),
.B(n_1377),
.Y(n_3172)
);

NAND2x1p5_ASAP7_75t_L g3173 ( 
.A(n_2728),
.B(n_2470),
.Y(n_3173)
);

NOR2xp33_ASAP7_75t_L g3174 ( 
.A(n_2461),
.B(n_1383),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2733),
.Y(n_3175)
);

AOI22x1_ASAP7_75t_L g3176 ( 
.A1(n_2673),
.A2(n_1386),
.B1(n_1684),
.B2(n_1604),
.Y(n_3176)
);

BUFx8_ASAP7_75t_L g3177 ( 
.A(n_2728),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2492),
.B(n_1388),
.Y(n_3178)
);

AO22x2_ASAP7_75t_L g3179 ( 
.A1(n_2647),
.A2(n_1583),
.B1(n_1609),
.B2(n_1349),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2639),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2643),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2639),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2642),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2642),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2759),
.Y(n_3185)
);

AOI22x1_ASAP7_75t_L g3186 ( 
.A1(n_2520),
.A2(n_2521),
.B1(n_2635),
.B2(n_2744),
.Y(n_3186)
);

AND2x4_ASAP7_75t_L g3187 ( 
.A(n_2676),
.B(n_1583),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2774),
.B(n_1390),
.Y(n_3188)
);

NOR2x1p5_ASAP7_75t_L g3189 ( 
.A(n_2478),
.B(n_1391),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2603),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2746),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2748),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2824),
.B(n_2774),
.Y(n_3193)
);

NOR2xp33_ASAP7_75t_L g3194 ( 
.A(n_2564),
.B(n_1392),
.Y(n_3194)
);

OR2x2_ASAP7_75t_SL g3195 ( 
.A(n_2539),
.B(n_2528),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2742),
.Y(n_3196)
);

INVxp67_ASAP7_75t_L g3197 ( 
.A(n_2587),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2713),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2695),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2702),
.Y(n_3200)
);

AND2x2_ASAP7_75t_SL g3201 ( 
.A(n_2445),
.B(n_1684),
.Y(n_3201)
);

NAND2x1p5_ASAP7_75t_L g3202 ( 
.A(n_2524),
.B(n_2532),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2603),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2700),
.Y(n_3204)
);

INVx2_ASAP7_75t_SL g3205 ( 
.A(n_2601),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2633),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_2654),
.Y(n_3207)
);

AOI22xp5_ASAP7_75t_L g3208 ( 
.A1(n_2687),
.A2(n_2648),
.B1(n_2664),
.B2(n_2657),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_SL g3209 ( 
.A(n_2697),
.B(n_1640),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2824),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_2701),
.B(n_1645),
.Y(n_3211)
);

OAI22xp33_ASAP7_75t_L g3212 ( 
.A1(n_2546),
.A2(n_1424),
.B1(n_1426),
.B2(n_1425),
.Y(n_3212)
);

INVxp67_ASAP7_75t_L g3213 ( 
.A(n_2809),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2824),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2722),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2680),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2712),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_2487),
.B(n_1441),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2723),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2589),
.B(n_1442),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2763),
.B(n_1449),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2782),
.B(n_1450),
.Y(n_3222)
);

INVx3_ASAP7_75t_L g3223 ( 
.A(n_2599),
.Y(n_3223)
);

NAND2x1p5_ASAP7_75t_L g3224 ( 
.A(n_2787),
.B(n_2797),
.Y(n_3224)
);

A2O1A1Ixp33_ASAP7_75t_L g3225 ( 
.A1(n_2610),
.A2(n_1617),
.B(n_1719),
.C(n_1609),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_2447),
.B(n_1455),
.Y(n_3226)
);

NAND2x1p5_ASAP7_75t_L g3227 ( 
.A(n_2730),
.B(n_1386),
.Y(n_3227)
);

AOI22xp5_ASAP7_75t_SL g3228 ( 
.A1(n_2599),
.A2(n_1462),
.B1(n_1468),
.B2(n_1467),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2722),
.Y(n_3229)
);

NAND2x1p5_ASAP7_75t_L g3230 ( 
.A(n_2599),
.B(n_1386),
.Y(n_3230)
);

AOI22xp33_ASAP7_75t_L g3231 ( 
.A1(n_2511),
.A2(n_1476),
.B1(n_1482),
.B2(n_1475),
.Y(n_3231)
);

CKINVDCx5p33_ASAP7_75t_R g3232 ( 
.A(n_2722),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2773),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2785),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_L g3235 ( 
.A(n_2823),
.B(n_1484),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2446),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_2430),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2446),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2479),
.Y(n_3239)
);

OAI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_2753),
.A2(n_1492),
.B1(n_1500),
.B2(n_1494),
.Y(n_3240)
);

AOI22xp5_ASAP7_75t_L g3241 ( 
.A1(n_2441),
.A2(n_1518),
.B1(n_1531),
.B2(n_1523),
.Y(n_3241)
);

INVx3_ASAP7_75t_L g3242 ( 
.A(n_2569),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_2823),
.B(n_1534),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2446),
.Y(n_3244)
);

NAND3xp33_ASAP7_75t_L g3245 ( 
.A(n_2553),
.B(n_1604),
.C(n_1386),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2437),
.B(n_1537),
.Y(n_3246)
);

INVxp67_ASAP7_75t_L g3247 ( 
.A(n_2431),
.Y(n_3247)
);

OAI22xp5_ASAP7_75t_L g3248 ( 
.A1(n_2753),
.A2(n_1546),
.B1(n_1548),
.B2(n_1539),
.Y(n_3248)
);

AND2x4_ASAP7_75t_L g3249 ( 
.A(n_2437),
.B(n_1617),
.Y(n_3249)
);

AND2x4_ASAP7_75t_L g3250 ( 
.A(n_2437),
.B(n_1719),
.Y(n_3250)
);

INVx2_ASAP7_75t_SL g3251 ( 
.A(n_2815),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_2446),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2823),
.B(n_1549),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2446),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2446),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_2446),
.Y(n_3256)
);

INVx3_ASAP7_75t_L g3257 ( 
.A(n_2569),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2446),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2437),
.B(n_1553),
.Y(n_3259)
);

A2O1A1Ixp33_ASAP7_75t_L g3260 ( 
.A1(n_2525),
.A2(n_1724),
.B(n_1604),
.C(n_1686),
.Y(n_3260)
);

INVx3_ASAP7_75t_L g3261 ( 
.A(n_2569),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2446),
.Y(n_3262)
);

CKINVDCx5p33_ASAP7_75t_R g3263 ( 
.A(n_2434),
.Y(n_3263)
);

OAI22xp5_ASAP7_75t_SL g3264 ( 
.A1(n_2434),
.A2(n_1648),
.B1(n_1663),
.B2(n_1638),
.Y(n_3264)
);

HB1xp67_ASAP7_75t_L g3265 ( 
.A(n_2823),
.Y(n_3265)
);

INVx2_ASAP7_75t_SL g3266 ( 
.A(n_2815),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2446),
.Y(n_3267)
);

AOI22x1_ASAP7_75t_L g3268 ( 
.A1(n_2540),
.A2(n_1684),
.B1(n_1686),
.B2(n_1604),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2446),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2446),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_2479),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2446),
.Y(n_3272)
);

AND2x4_ASAP7_75t_L g3273 ( 
.A(n_2437),
.B(n_1724),
.Y(n_3273)
);

BUFx6f_ASAP7_75t_L g3274 ( 
.A(n_2750),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2446),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_2823),
.B(n_1558),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_2437),
.B(n_1585),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_2446),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2446),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2446),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2446),
.Y(n_3281)
);

INVx2_ASAP7_75t_L g3282 ( 
.A(n_2479),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2479),
.Y(n_3283)
);

NOR2xp33_ASAP7_75t_L g3284 ( 
.A(n_2823),
.B(n_1586),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2446),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2446),
.Y(n_3286)
);

AND2x6_ASAP7_75t_L g3287 ( 
.A(n_2437),
.B(n_1684),
.Y(n_3287)
);

AO22x2_ASAP7_75t_L g3288 ( 
.A1(n_2679),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2446),
.Y(n_3289)
);

INVxp67_ASAP7_75t_L g3290 ( 
.A(n_2431),
.Y(n_3290)
);

INVxp67_ASAP7_75t_L g3291 ( 
.A(n_2431),
.Y(n_3291)
);

BUFx8_ASAP7_75t_L g3292 ( 
.A(n_2481),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2446),
.Y(n_3293)
);

AO22x2_ASAP7_75t_L g3294 ( 
.A1(n_2679),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2446),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2446),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2446),
.Y(n_3297)
);

AND2x4_ASAP7_75t_L g3298 ( 
.A(n_2437),
.B(n_4),
.Y(n_3298)
);

AO22x2_ASAP7_75t_L g3299 ( 
.A1(n_2679),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2446),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2446),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_2446),
.Y(n_3302)
);

A2O1A1Ixp33_ASAP7_75t_L g3303 ( 
.A1(n_2525),
.A2(n_1686),
.B(n_1120),
.C(n_1422),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_2437),
.B(n_1588),
.Y(n_3304)
);

AND2x4_ASAP7_75t_L g3305 ( 
.A(n_2437),
.B(n_4),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2446),
.Y(n_3306)
);

AO22x2_ASAP7_75t_L g3307 ( 
.A1(n_2679),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_3307)
);

AOI22xp33_ASAP7_75t_L g3308 ( 
.A1(n_2806),
.A2(n_1590),
.B1(n_1614),
.B2(n_1598),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_SL g3309 ( 
.A(n_2557),
.B(n_1626),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_2446),
.Y(n_3310)
);

AOI22xp5_ASAP7_75t_L g3311 ( 
.A1(n_2441),
.A2(n_1615),
.B1(n_1622),
.B2(n_1618),
.Y(n_3311)
);

BUFx8_ASAP7_75t_L g3312 ( 
.A(n_2481),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_2479),
.Y(n_3313)
);

NAND2x1p5_ASAP7_75t_L g3314 ( 
.A(n_2815),
.B(n_1686),
.Y(n_3314)
);

INVx3_ASAP7_75t_L g3315 ( 
.A(n_2569),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2446),
.Y(n_3316)
);

INVx2_ASAP7_75t_SL g3317 ( 
.A(n_2815),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2446),
.Y(n_3318)
);

INVx3_ASAP7_75t_L g3319 ( 
.A(n_2569),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2446),
.Y(n_3320)
);

CKINVDCx5p33_ASAP7_75t_R g3321 ( 
.A(n_2434),
.Y(n_3321)
);

CKINVDCx5p33_ASAP7_75t_R g3322 ( 
.A(n_2434),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2446),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_2823),
.B(n_1633),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2446),
.Y(n_3325)
);

BUFx3_ASAP7_75t_L g3326 ( 
.A(n_2430),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_2479),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2479),
.Y(n_3328)
);

CKINVDCx20_ASAP7_75t_R g3329 ( 
.A(n_2434),
.Y(n_3329)
);

AO22x2_ASAP7_75t_L g3330 ( 
.A1(n_2679),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_2806),
.A2(n_1666),
.B1(n_1671),
.B2(n_1667),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2437),
.B(n_1679),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_2446),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_2441),
.A2(n_1682),
.B1(n_1726),
.B2(n_1199),
.Y(n_3334)
);

AO22x2_ASAP7_75t_L g3335 ( 
.A1(n_2679),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_3335)
);

INVxp67_ASAP7_75t_L g3336 ( 
.A(n_2431),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_2446),
.Y(n_3337)
);

BUFx2_ASAP7_75t_L g3338 ( 
.A(n_2434),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_SL g3339 ( 
.A(n_2557),
.B(n_1199),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_L g3340 ( 
.A1(n_2806),
.A2(n_1120),
.B1(n_1422),
.B2(n_1078),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2479),
.Y(n_3341)
);

BUFx6f_ASAP7_75t_L g3342 ( 
.A(n_2750),
.Y(n_3342)
);

INVx2_ASAP7_75t_SL g3343 ( 
.A(n_2815),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2446),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2446),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_2823),
.B(n_9),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_2437),
.B(n_9),
.Y(n_3347)
);

INVxp67_ASAP7_75t_L g3348 ( 
.A(n_2431),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_2479),
.Y(n_3349)
);

AND2x4_ASAP7_75t_L g3350 ( 
.A(n_2437),
.B(n_10),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_2446),
.Y(n_3351)
);

INVxp67_ASAP7_75t_L g3352 ( 
.A(n_2431),
.Y(n_3352)
);

NAND2x1p5_ASAP7_75t_L g3353 ( 
.A(n_2815),
.B(n_1120),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_2437),
.B(n_10),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2446),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2446),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2446),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_2479),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2479),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_2437),
.B(n_11),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_2823),
.B(n_11),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_2823),
.B(n_11),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2446),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2446),
.Y(n_3364)
);

AND2x2_ASAP7_75t_L g3365 ( 
.A(n_2823),
.B(n_12),
.Y(n_3365)
);

NOR2xp33_ASAP7_75t_L g3366 ( 
.A(n_2823),
.B(n_12),
.Y(n_3366)
);

AND2x4_ASAP7_75t_L g3367 ( 
.A(n_2437),
.B(n_12),
.Y(n_3367)
);

INVx3_ASAP7_75t_L g3368 ( 
.A(n_2569),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2437),
.B(n_13),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_2479),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2479),
.Y(n_3371)
);

NAND2x1p5_ASAP7_75t_L g3372 ( 
.A(n_2815),
.B(n_1120),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_2437),
.B(n_14),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2446),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_2479),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2446),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2446),
.Y(n_3377)
);

BUFx2_ASAP7_75t_L g3378 ( 
.A(n_2434),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_2446),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2446),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_2437),
.B(n_14),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_2823),
.B(n_14),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2446),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_2823),
.B(n_15),
.Y(n_3384)
);

HB1xp67_ASAP7_75t_L g3385 ( 
.A(n_2823),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2446),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2446),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_2479),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_2437),
.B(n_15),
.Y(n_3389)
);

BUFx2_ASAP7_75t_L g3390 ( 
.A(n_2434),
.Y(n_3390)
);

AOI22xp33_ASAP7_75t_L g3391 ( 
.A1(n_2806),
.A2(n_1422),
.B1(n_18),
.B2(n_16),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_2446),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2446),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_L g3394 ( 
.A(n_2823),
.B(n_16),
.Y(n_3394)
);

OAI221xp5_ASAP7_75t_L g3395 ( 
.A1(n_2504),
.A2(n_1422),
.B1(n_18),
.B2(n_16),
.C(n_17),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_2823),
.B(n_17),
.Y(n_3396)
);

NAND2x1p5_ASAP7_75t_L g3397 ( 
.A(n_2815),
.B(n_19),
.Y(n_3397)
);

AND2x6_ASAP7_75t_L g3398 ( 
.A(n_2437),
.B(n_19),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_2437),
.B(n_20),
.Y(n_3399)
);

INVxp67_ASAP7_75t_L g3400 ( 
.A(n_2431),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2437),
.B(n_21),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2479),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2437),
.B(n_21),
.Y(n_3403)
);

AND2x6_ASAP7_75t_L g3404 ( 
.A(n_2437),
.B(n_22),
.Y(n_3404)
);

NAND2xp33_ASAP7_75t_L g3405 ( 
.A(n_2750),
.B(n_23),
.Y(n_3405)
);

NAND2x1p5_ASAP7_75t_L g3406 ( 
.A(n_2815),
.B(n_22),
.Y(n_3406)
);

NOR2xp33_ASAP7_75t_L g3407 ( 
.A(n_2823),
.B(n_22),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_2479),
.Y(n_3408)
);

NOR2xp33_ASAP7_75t_L g3409 ( 
.A(n_2823),
.B(n_23),
.Y(n_3409)
);

OAI22xp5_ASAP7_75t_L g3410 ( 
.A1(n_2753),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_3410)
);

AND2x4_ASAP7_75t_L g3411 ( 
.A(n_2437),
.B(n_24),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2479),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2446),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_2446),
.Y(n_3414)
);

NAND2x1p5_ASAP7_75t_L g3415 ( 
.A(n_2815),
.B(n_24),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2446),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_2479),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2446),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_2479),
.Y(n_3419)
);

INVx4_ASAP7_75t_L g3420 ( 
.A(n_2569),
.Y(n_3420)
);

NOR3xp33_ASAP7_75t_L g3421 ( 
.A(n_2557),
.B(n_27),
.C(n_26),
.Y(n_3421)
);

BUFx3_ASAP7_75t_L g3422 ( 
.A(n_2430),
.Y(n_3422)
);

AOI22x1_ASAP7_75t_L g3423 ( 
.A1(n_2540),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_2446),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2437),
.B(n_25),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_2479),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2446),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_2479),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_SL g3429 ( 
.A(n_2557),
.B(n_28),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_2446),
.Y(n_3430)
);

A2O1A1Ixp33_ASAP7_75t_L g3431 ( 
.A1(n_2525),
.A2(n_30),
.B(n_27),
.C(n_29),
.Y(n_3431)
);

INVxp67_ASAP7_75t_SL g3432 ( 
.A(n_2431),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_SL g3433 ( 
.A(n_2557),
.B(n_31),
.Y(n_3433)
);

NAND2xp33_ASAP7_75t_L g3434 ( 
.A(n_2750),
.B(n_31),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2446),
.Y(n_3435)
);

AND2x4_ASAP7_75t_L g3436 ( 
.A(n_2437),
.B(n_30),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2446),
.Y(n_3437)
);

NAND3xp33_ASAP7_75t_L g3438 ( 
.A(n_2553),
.B(n_31),
.C(n_32),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_L g3439 ( 
.A1(n_2806),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_3439)
);

INVxp67_ASAP7_75t_L g3440 ( 
.A(n_2431),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_2437),
.B(n_32),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_2437),
.B(n_33),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_2823),
.B(n_33),
.Y(n_3443)
);

INVxp67_ASAP7_75t_L g3444 ( 
.A(n_2431),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_2823),
.B(n_34),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_2437),
.B(n_34),
.Y(n_3446)
);

INVx3_ASAP7_75t_L g3447 ( 
.A(n_2569),
.Y(n_3447)
);

AO22x2_ASAP7_75t_L g3448 ( 
.A1(n_2679),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_2557),
.B(n_36),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_2446),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_2446),
.Y(n_3451)
);

AO22x2_ASAP7_75t_L g3452 ( 
.A1(n_2679),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_2557),
.B(n_38),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_2446),
.Y(n_3454)
);

NOR3xp33_ASAP7_75t_L g3455 ( 
.A(n_2557),
.B(n_39),
.C(n_38),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_2446),
.Y(n_3456)
);

NAND2x1p5_ASAP7_75t_L g3457 ( 
.A(n_2815),
.B(n_37),
.Y(n_3457)
);

AND2x4_ASAP7_75t_L g3458 ( 
.A(n_2437),
.B(n_39),
.Y(n_3458)
);

CKINVDCx5p33_ASAP7_75t_R g3459 ( 
.A(n_2434),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_2446),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_2446),
.Y(n_3461)
);

AND2x4_ASAP7_75t_L g3462 ( 
.A(n_2437),
.B(n_39),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_2823),
.B(n_40),
.Y(n_3463)
);

INVx2_ASAP7_75t_SL g3464 ( 
.A(n_2815),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2446),
.Y(n_3465)
);

INVx3_ASAP7_75t_L g3466 ( 
.A(n_2569),
.Y(n_3466)
);

BUFx6f_ASAP7_75t_L g3467 ( 
.A(n_2750),
.Y(n_3467)
);

NOR2xp33_ASAP7_75t_L g3468 ( 
.A(n_2823),
.B(n_40),
.Y(n_3468)
);

AOI22xp5_ASAP7_75t_L g3469 ( 
.A1(n_2441),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_3469)
);

AO22x2_ASAP7_75t_L g3470 ( 
.A1(n_2679),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_3470)
);

CKINVDCx16_ASAP7_75t_R g3471 ( 
.A(n_2434),
.Y(n_3471)
);

NOR2xp33_ASAP7_75t_L g3472 ( 
.A(n_2823),
.B(n_43),
.Y(n_3472)
);

A2O1A1Ixp33_ASAP7_75t_L g3473 ( 
.A1(n_2525),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_2479),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_2479),
.Y(n_3475)
);

INVxp67_ASAP7_75t_L g3476 ( 
.A(n_2431),
.Y(n_3476)
);

AOI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_2441),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_2446),
.Y(n_3478)
);

AND2x4_ASAP7_75t_L g3479 ( 
.A(n_2437),
.B(n_46),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_2430),
.Y(n_3480)
);

BUFx8_ASAP7_75t_L g3481 ( 
.A(n_2481),
.Y(n_3481)
);

INVx2_ASAP7_75t_SL g3482 ( 
.A(n_2815),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_2479),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_2446),
.Y(n_3484)
);

NAND3x1_ASAP7_75t_L g3485 ( 
.A(n_2607),
.B(n_47),
.C(n_48),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_2479),
.Y(n_3486)
);

HB1xp67_ASAP7_75t_L g3487 ( 
.A(n_3265),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_2963),
.A2(n_48),
.B(n_49),
.Y(n_3488)
);

NOR3xp33_ASAP7_75t_L g3489 ( 
.A(n_3159),
.B(n_49),
.C(n_50),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2896),
.B(n_49),
.Y(n_3490)
);

INVx11_ASAP7_75t_L g3491 ( 
.A(n_2849),
.Y(n_3491)
);

OAI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_2970),
.A2(n_51),
.B(n_52),
.Y(n_3492)
);

OAI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_2937),
.A2(n_52),
.B(n_53),
.Y(n_3493)
);

O2A1O1Ixp33_ASAP7_75t_L g3494 ( 
.A1(n_3021),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_3494)
);

A2O1A1Ixp33_ASAP7_75t_L g3495 ( 
.A1(n_2983),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3000),
.A2(n_54),
.B(n_55),
.Y(n_3496)
);

CKINVDCx10_ASAP7_75t_R g3497 ( 
.A(n_3471),
.Y(n_3497)
);

AO21x2_ASAP7_75t_L g3498 ( 
.A1(n_3004),
.A2(n_55),
.B(n_56),
.Y(n_3498)
);

BUFx6f_ASAP7_75t_L g3499 ( 
.A(n_2996),
.Y(n_3499)
);

INVx8_ASAP7_75t_L g3500 ( 
.A(n_2879),
.Y(n_3500)
);

BUFx6f_ASAP7_75t_L g3501 ( 
.A(n_2996),
.Y(n_3501)
);

O2A1O1Ixp33_ASAP7_75t_SL g3502 ( 
.A1(n_3193),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3005),
.A2(n_3014),
.B(n_3008),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_SL g3504 ( 
.A(n_3201),
.B(n_814),
.Y(n_3504)
);

BUFx12f_ASAP7_75t_L g3505 ( 
.A(n_2849),
.Y(n_3505)
);

OAI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3006),
.A2(n_57),
.B(n_59),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_2839),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_2912),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3076),
.B(n_3077),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3080),
.B(n_57),
.Y(n_3510)
);

BUFx6f_ASAP7_75t_L g3511 ( 
.A(n_2996),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3030),
.A2(n_60),
.B(n_61),
.Y(n_3512)
);

AOI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_3031),
.A2(n_60),
.B(n_61),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3084),
.B(n_60),
.Y(n_3514)
);

AO21x1_ASAP7_75t_L g3515 ( 
.A1(n_3210),
.A2(n_3214),
.B(n_3165),
.Y(n_3515)
);

O2A1O1Ixp33_ASAP7_75t_L g3516 ( 
.A1(n_3129),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3087),
.B(n_62),
.Y(n_3517)
);

BUFx2_ASAP7_75t_L g3518 ( 
.A(n_3329),
.Y(n_3518)
);

AND2x6_ASAP7_75t_L g3519 ( 
.A(n_3157),
.B(n_62),
.Y(n_3519)
);

AND2x4_ASAP7_75t_L g3520 ( 
.A(n_2861),
.B(n_63),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3067),
.B(n_63),
.Y(n_3521)
);

OAI22xp5_ASAP7_75t_L g3522 ( 
.A1(n_2894),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_2852),
.Y(n_3523)
);

AOI21x1_ASAP7_75t_L g3524 ( 
.A1(n_2923),
.A2(n_65),
.B(n_66),
.Y(n_3524)
);

A2O1A1Ixp33_ASAP7_75t_L g3525 ( 
.A1(n_2953),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3105),
.B(n_67),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_3176),
.A2(n_68),
.B(n_69),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3106),
.B(n_68),
.Y(n_3528)
);

OAI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_2894),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3108),
.B(n_70),
.Y(n_3530)
);

NOR2xp33_ASAP7_75t_L g3531 ( 
.A(n_3025),
.B(n_71),
.Y(n_3531)
);

AOI21x1_ASAP7_75t_L g3532 ( 
.A1(n_2923),
.A2(n_72),
.B(n_73),
.Y(n_3532)
);

BUFx6f_ASAP7_75t_L g3533 ( 
.A(n_3073),
.Y(n_3533)
);

BUFx6f_ASAP7_75t_L g3534 ( 
.A(n_3073),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_2927),
.Y(n_3535)
);

BUFx4f_ASAP7_75t_L g3536 ( 
.A(n_3398),
.Y(n_3536)
);

INVx2_ASAP7_75t_L g3537 ( 
.A(n_2858),
.Y(n_3537)
);

AOI21xp5_ASAP7_75t_L g3538 ( 
.A1(n_3233),
.A2(n_74),
.B(n_75),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3111),
.B(n_74),
.Y(n_3539)
);

AOI21xp5_ASAP7_75t_L g3540 ( 
.A1(n_3234),
.A2(n_75),
.B(n_76),
.Y(n_3540)
);

O2A1O1Ixp33_ASAP7_75t_L g3541 ( 
.A1(n_3429),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_2951),
.B(n_76),
.Y(n_3542)
);

OAI21xp5_ASAP7_75t_L g3543 ( 
.A1(n_2876),
.A2(n_2943),
.B(n_2941),
.Y(n_3543)
);

O2A1O1Ixp33_ASAP7_75t_L g3544 ( 
.A1(n_3433),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_3544)
);

A2O1A1Ixp33_ASAP7_75t_L g3545 ( 
.A1(n_2944),
.A2(n_2948),
.B(n_2945),
.C(n_2934),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_2860),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3268),
.A2(n_77),
.B(n_79),
.Y(n_3547)
);

AND2x6_ASAP7_75t_L g3548 ( 
.A(n_3157),
.B(n_79),
.Y(n_3548)
);

NOR2xp67_ASAP7_75t_L g3549 ( 
.A(n_3420),
.B(n_80),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2931),
.Y(n_3550)
);

BUFx2_ASAP7_75t_L g3551 ( 
.A(n_2982),
.Y(n_3551)
);

OA22x2_ASAP7_75t_L g3552 ( 
.A1(n_2900),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_3552)
);

AOI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_2980),
.A2(n_80),
.B(n_81),
.Y(n_3553)
);

OAI22xp5_ASAP7_75t_L g3554 ( 
.A1(n_2899),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_3554)
);

OAI321xp33_ASAP7_75t_L g3555 ( 
.A1(n_3395),
.A2(n_85),
.A3(n_87),
.B1(n_83),
.B2(n_84),
.C(n_86),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_2905),
.B(n_83),
.Y(n_3556)
);

AOI21xp5_ASAP7_75t_L g3557 ( 
.A1(n_3088),
.A2(n_85),
.B(n_86),
.Y(n_3557)
);

AOI21xp5_ASAP7_75t_L g3558 ( 
.A1(n_3339),
.A2(n_86),
.B(n_87),
.Y(n_3558)
);

OR2x2_ASAP7_75t_L g3559 ( 
.A(n_3385),
.B(n_87),
.Y(n_3559)
);

AOI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_2958),
.A2(n_88),
.B(n_89),
.Y(n_3560)
);

AOI21x1_ASAP7_75t_L g3561 ( 
.A1(n_2924),
.A2(n_3207),
.B(n_3229),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_2864),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_2877),
.Y(n_3563)
);

A2O1A1Ixp33_ASAP7_75t_L g3564 ( 
.A1(n_2932),
.A2(n_3115),
.B(n_3134),
.C(n_3133),
.Y(n_3564)
);

O2A1O1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_3449),
.A2(n_90),
.B(n_88),
.C(n_89),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_2837),
.B(n_88),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_3483),
.A2(n_89),
.B(n_90),
.Y(n_3567)
);

A2O1A1Ixp33_ASAP7_75t_L g3568 ( 
.A1(n_3438),
.A2(n_93),
.B(n_91),
.C(n_92),
.Y(n_3568)
);

AOI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3486),
.A2(n_91),
.B(n_92),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_2883),
.A2(n_91),
.B(n_93),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_2892),
.A2(n_94),
.B(n_95),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_2838),
.B(n_2832),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_2924),
.Y(n_3573)
);

AOI22xp5_ASAP7_75t_L g3574 ( 
.A1(n_2828),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_SL g3575 ( 
.A(n_3228),
.B(n_3208),
.Y(n_3575)
);

A2O1A1Ixp33_ASAP7_75t_L g3576 ( 
.A1(n_2938),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_2834),
.B(n_96),
.Y(n_3577)
);

AOI21xp5_ASAP7_75t_L g3578 ( 
.A1(n_2897),
.A2(n_97),
.B(n_98),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_2835),
.B(n_99),
.Y(n_3579)
);

OAI21x1_ASAP7_75t_L g3580 ( 
.A1(n_3186),
.A2(n_99),
.B(n_100),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_2917),
.A2(n_99),
.B(n_100),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3236),
.B(n_100),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_2925),
.A2(n_101),
.B(n_102),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3238),
.Y(n_3584)
);

O2A1O1Ixp33_ASAP7_75t_L g3585 ( 
.A1(n_3453),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3244),
.B(n_101),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3252),
.B(n_102),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3254),
.B(n_103),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3255),
.B(n_103),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3474),
.A2(n_104),
.B(n_105),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_3475),
.A2(n_104),
.B(n_105),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_2935),
.A2(n_104),
.B(n_105),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3256),
.B(n_106),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3239),
.A2(n_106),
.B(n_107),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3271),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3258),
.B(n_107),
.Y(n_3596)
);

OA21x2_ASAP7_75t_L g3597 ( 
.A1(n_3303),
.A2(n_108),
.B(n_109),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_SL g3598 ( 
.A(n_2846),
.B(n_814),
.Y(n_3598)
);

AO22x1_ASAP7_75t_L g3599 ( 
.A1(n_3398),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_3599)
);

AND2x6_ASAP7_75t_L g3600 ( 
.A(n_3157),
.B(n_108),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3262),
.B(n_3267),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3269),
.B(n_109),
.Y(n_3602)
);

HB1xp67_ASAP7_75t_L g3603 ( 
.A(n_2829),
.Y(n_3603)
);

INVxp67_ASAP7_75t_L g3604 ( 
.A(n_3432),
.Y(n_3604)
);

NOR3xp33_ASAP7_75t_L g3605 ( 
.A(n_3048),
.B(n_111),
.C(n_112),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3270),
.B(n_111),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3272),
.B(n_112),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3282),
.A2(n_112),
.B(n_113),
.Y(n_3608)
);

AOI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3283),
.A2(n_113),
.B(n_114),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3275),
.B(n_113),
.Y(n_3610)
);

NOR2xp33_ASAP7_75t_SL g3611 ( 
.A(n_3263),
.B(n_114),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3313),
.A2(n_114),
.B(n_115),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3278),
.B(n_115),
.Y(n_3613)
);

BUFx3_ASAP7_75t_L g3614 ( 
.A(n_3158),
.Y(n_3614)
);

O2A1O1Ixp33_ASAP7_75t_L g3615 ( 
.A1(n_3019),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_L g3616 ( 
.A(n_2933),
.B(n_116),
.Y(n_3616)
);

INVx4_ASAP7_75t_L g3617 ( 
.A(n_2885),
.Y(n_3617)
);

HB1xp67_ASAP7_75t_L g3618 ( 
.A(n_3321),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_SL g3619 ( 
.A(n_2984),
.B(n_816),
.Y(n_3619)
);

AOI22xp5_ASAP7_75t_L g3620 ( 
.A1(n_2828),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_3620)
);

OAI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_2911),
.A2(n_117),
.B(n_119),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3327),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_SL g3623 ( 
.A(n_2994),
.B(n_817),
.Y(n_3623)
);

A2O1A1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_3421),
.A2(n_123),
.B(n_120),
.C(n_121),
.Y(n_3624)
);

AOI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_3328),
.A2(n_120),
.B(n_121),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3279),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_3341),
.A2(n_120),
.B(n_121),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3349),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3280),
.B(n_124),
.Y(n_3629)
);

NAND3xp33_ASAP7_75t_L g3630 ( 
.A(n_3001),
.B(n_124),
.C(n_125),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_3358),
.A2(n_3370),
.B(n_3359),
.Y(n_3631)
);

AND2x4_ASAP7_75t_L g3632 ( 
.A(n_2861),
.B(n_124),
.Y(n_3632)
);

NOR2xp33_ASAP7_75t_L g3633 ( 
.A(n_2936),
.B(n_125),
.Y(n_3633)
);

BUFx3_ASAP7_75t_L g3634 ( 
.A(n_3158),
.Y(n_3634)
);

A2O1A1Ixp33_ASAP7_75t_L g3635 ( 
.A1(n_3455),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_3635)
);

BUFx8_ASAP7_75t_L g3636 ( 
.A(n_3138),
.Y(n_3636)
);

NOR2xp33_ASAP7_75t_L g3637 ( 
.A(n_2950),
.B(n_126),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_SL g3638 ( 
.A(n_3110),
.B(n_817),
.Y(n_3638)
);

AND2x4_ASAP7_75t_L g3639 ( 
.A(n_3420),
.B(n_126),
.Y(n_3639)
);

AOI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_3371),
.A2(n_127),
.B(n_128),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3281),
.B(n_127),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3285),
.B(n_129),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_3375),
.A2(n_129),
.B(n_130),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_3388),
.A2(n_3408),
.B(n_3402),
.Y(n_3644)
);

INVx2_ASAP7_75t_SL g3645 ( 
.A(n_3177),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3286),
.B(n_3289),
.Y(n_3646)
);

OAI22xp5_ASAP7_75t_L g3647 ( 
.A1(n_2899),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3293),
.B(n_130),
.Y(n_3648)
);

INVxp67_ASAP7_75t_L g3649 ( 
.A(n_3243),
.Y(n_3649)
);

OAI22xp5_ASAP7_75t_L g3650 ( 
.A1(n_2902),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_3650)
);

NOR2x1p5_ASAP7_75t_L g3651 ( 
.A(n_3322),
.B(n_3459),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3412),
.Y(n_3652)
);

BUFx12f_ASAP7_75t_L g3653 ( 
.A(n_3292),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3295),
.B(n_131),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3296),
.B(n_132),
.Y(n_3655)
);

AND2x4_ASAP7_75t_L g3656 ( 
.A(n_2915),
.B(n_132),
.Y(n_3656)
);

AOI22xp33_ASAP7_75t_L g3657 ( 
.A1(n_2914),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3297),
.B(n_133),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3417),
.A2(n_134),
.B(n_136),
.Y(n_3659)
);

AOI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_3419),
.A2(n_134),
.B(n_136),
.Y(n_3660)
);

O2A1O1Ixp33_ASAP7_75t_L g3661 ( 
.A1(n_3131),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3426),
.A2(n_137),
.B(n_138),
.Y(n_3662)
);

NOR2xp33_ASAP7_75t_L g3663 ( 
.A(n_2959),
.B(n_137),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3300),
.B(n_138),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3428),
.Y(n_3665)
);

OAI21xp33_ASAP7_75t_SL g3666 ( 
.A1(n_3050),
.A2(n_139),
.B(n_140),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3301),
.B(n_139),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3302),
.B(n_139),
.Y(n_3668)
);

INVx4_ASAP7_75t_L g3669 ( 
.A(n_2851),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3306),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3310),
.B(n_3316),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3260),
.A2(n_140),
.B(n_141),
.Y(n_3672)
);

AO21x1_ASAP7_75t_L g3673 ( 
.A1(n_3410),
.A2(n_819),
.B(n_818),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_2895),
.B(n_3069),
.Y(n_3674)
);

AOI22xp5_ASAP7_75t_L g3675 ( 
.A1(n_2902),
.A2(n_143),
.B1(n_140),
.B2(n_142),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3318),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3320),
.Y(n_3677)
);

AOI21xp5_ASAP7_75t_L g3678 ( 
.A1(n_2967),
.A2(n_142),
.B(n_143),
.Y(n_3678)
);

AOI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_2969),
.A2(n_142),
.B(n_143),
.Y(n_3679)
);

AOI21xp5_ASAP7_75t_L g3680 ( 
.A1(n_2986),
.A2(n_144),
.B(n_145),
.Y(n_3680)
);

AO21x1_ASAP7_75t_L g3681 ( 
.A1(n_3405),
.A2(n_821),
.B(n_820),
.Y(n_3681)
);

A2O1A1Ixp33_ASAP7_75t_L g3682 ( 
.A1(n_3431),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3323),
.B(n_146),
.Y(n_3683)
);

INVx1_ASAP7_75t_SL g3684 ( 
.A(n_3037),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_3325),
.Y(n_3685)
);

AO32x2_ASAP7_75t_L g3686 ( 
.A1(n_2916),
.A2(n_148),
.A3(n_146),
.B1(n_147),
.B2(n_149),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_SL g3687 ( 
.A(n_3298),
.B(n_3305),
.Y(n_3687)
);

AOI22xp33_ASAP7_75t_L g3688 ( 
.A1(n_3013),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_3688)
);

OR2x2_ASAP7_75t_L g3689 ( 
.A(n_2882),
.B(n_149),
.Y(n_3689)
);

OAI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_2964),
.A2(n_3391),
.B1(n_3305),
.B2(n_3350),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3333),
.B(n_150),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_2989),
.A2(n_150),
.B(n_151),
.Y(n_3692)
);

BUFx12f_ASAP7_75t_L g3693 ( 
.A(n_3292),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_2952),
.A2(n_150),
.B(n_151),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3337),
.B(n_152),
.Y(n_3695)
);

OAI21xp5_ASAP7_75t_L g3696 ( 
.A1(n_2939),
.A2(n_152),
.B(n_153),
.Y(n_3696)
);

AOI21x1_ASAP7_75t_L g3697 ( 
.A1(n_3188),
.A2(n_152),
.B(n_153),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3344),
.Y(n_3698)
);

NOR3xp33_ASAP7_75t_L g3699 ( 
.A(n_3065),
.B(n_154),
.C(n_155),
.Y(n_3699)
);

OAI22xp5_ASAP7_75t_L g3700 ( 
.A1(n_2964),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3345),
.B(n_155),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_SL g3702 ( 
.A(n_3298),
.B(n_821),
.Y(n_3702)
);

AND2x2_ASAP7_75t_SL g3703 ( 
.A(n_3350),
.B(n_156),
.Y(n_3703)
);

AOI22x1_ASAP7_75t_L g3704 ( 
.A1(n_3074),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_3704)
);

BUFx6f_ASAP7_75t_L g3705 ( 
.A(n_3073),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3288),
.B(n_157),
.Y(n_3706)
);

OAI22xp5_ASAP7_75t_L g3707 ( 
.A1(n_3367),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_3434),
.A2(n_158),
.B(n_159),
.Y(n_3708)
);

HB1xp67_ASAP7_75t_L g3709 ( 
.A(n_3247),
.Y(n_3709)
);

O2A1O1Ixp33_ASAP7_75t_L g3710 ( 
.A1(n_2862),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_3710)
);

O2A1O1Ixp5_ASAP7_75t_SL g3711 ( 
.A1(n_3016),
.A2(n_823),
.B(n_824),
.C(n_822),
.Y(n_3711)
);

CKINVDCx5p33_ASAP7_75t_R g3712 ( 
.A(n_3312),
.Y(n_3712)
);

OAI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3367),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_SL g3714 ( 
.A(n_3411),
.B(n_822),
.Y(n_3714)
);

A2O1A1Ixp33_ASAP7_75t_L g3715 ( 
.A1(n_3473),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3288),
.B(n_162),
.Y(n_3716)
);

OAI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_2946),
.A2(n_163),
.B(n_165),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_3148),
.A2(n_165),
.B(n_166),
.Y(n_3718)
);

AND2x6_ASAP7_75t_L g3719 ( 
.A(n_3411),
.B(n_3436),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3161),
.A2(n_165),
.B(n_166),
.Y(n_3720)
);

INVxp67_ASAP7_75t_L g3721 ( 
.A(n_3253),
.Y(n_3721)
);

INVx8_ASAP7_75t_L g3722 ( 
.A(n_2988),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_3169),
.A2(n_167),
.B(n_168),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3351),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3164),
.A2(n_168),
.B(n_169),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3294),
.B(n_168),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3355),
.Y(n_3727)
);

OAI21xp33_ASAP7_75t_L g3728 ( 
.A1(n_2920),
.A2(n_169),
.B(n_170),
.Y(n_3728)
);

O2A1O1Ixp33_ASAP7_75t_L g3729 ( 
.A1(n_3056),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_3729)
);

NAND2x1p5_ASAP7_75t_L g3730 ( 
.A(n_3237),
.B(n_170),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3356),
.B(n_171),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3357),
.Y(n_3732)
);

NOR2xp33_ASAP7_75t_L g3733 ( 
.A(n_2918),
.B(n_172),
.Y(n_3733)
);

INVx3_ASAP7_75t_L g3734 ( 
.A(n_3274),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3363),
.B(n_172),
.Y(n_3735)
);

AOI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_3168),
.A2(n_173),
.B(n_174),
.Y(n_3736)
);

OAI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_2973),
.A2(n_173),
.B(n_174),
.Y(n_3737)
);

BUFx2_ASAP7_75t_L g3738 ( 
.A(n_2982),
.Y(n_3738)
);

AOI21x1_ASAP7_75t_L g3739 ( 
.A1(n_3245),
.A2(n_173),
.B(n_174),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_SL g3740 ( 
.A(n_3436),
.B(n_823),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3364),
.Y(n_3741)
);

O2A1O1Ixp33_ASAP7_75t_SL g3742 ( 
.A1(n_3223),
.A2(n_177),
.B(n_175),
.C(n_176),
.Y(n_3742)
);

OAI22xp5_ASAP7_75t_L g3743 ( 
.A1(n_3458),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3374),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3376),
.B(n_175),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_2974),
.A2(n_177),
.B(n_178),
.Y(n_3746)
);

INVx4_ASAP7_75t_L g3747 ( 
.A(n_3326),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_3377),
.B(n_178),
.Y(n_3748)
);

AND2x4_ASAP7_75t_L g3749 ( 
.A(n_2915),
.B(n_178),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3294),
.B(n_179),
.Y(n_3750)
);

NOR2xp33_ASAP7_75t_L g3751 ( 
.A(n_3197),
.B(n_179),
.Y(n_3751)
);

INVxp67_ASAP7_75t_L g3752 ( 
.A(n_3276),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_SL g3753 ( 
.A(n_3458),
.B(n_825),
.Y(n_3753)
);

BUFx2_ASAP7_75t_L g3754 ( 
.A(n_3132),
.Y(n_3754)
);

NOR2xp33_ASAP7_75t_L g3755 ( 
.A(n_2830),
.B(n_180),
.Y(n_3755)
);

AOI21x1_ASAP7_75t_L g3756 ( 
.A1(n_3347),
.A2(n_180),
.B(n_181),
.Y(n_3756)
);

AOI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_2826),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_3757)
);

AOI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_2921),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3225),
.A2(n_183),
.B(n_184),
.Y(n_3759)
);

NOR2xp33_ASAP7_75t_L g3760 ( 
.A(n_3119),
.B(n_184),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3379),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_SL g3762 ( 
.A(n_3462),
.B(n_3479),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3380),
.B(n_185),
.Y(n_3763)
);

INVx3_ASAP7_75t_L g3764 ( 
.A(n_3274),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3007),
.A2(n_185),
.B(n_186),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3383),
.Y(n_3766)
);

AOI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_2957),
.A2(n_185),
.B(n_186),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_2962),
.A2(n_186),
.B(n_187),
.Y(n_3768)
);

NAND3xp33_ASAP7_75t_L g3769 ( 
.A(n_3340),
.B(n_187),
.C(n_188),
.Y(n_3769)
);

INVx1_ASAP7_75t_SL g3770 ( 
.A(n_3422),
.Y(n_3770)
);

NAND3xp33_ASAP7_75t_SL g3771 ( 
.A(n_2871),
.B(n_187),
.C(n_188),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3386),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_2965),
.A2(n_189),
.B(n_190),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3387),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3392),
.B(n_189),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3393),
.B(n_190),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3299),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3413),
.B(n_192),
.Y(n_3778)
);

AOI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_2966),
.A2(n_193),
.B(n_194),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_3299),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_3780)
);

AOI21xp5_ASAP7_75t_L g3781 ( 
.A1(n_2968),
.A2(n_195),
.B(n_196),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_SL g3782 ( 
.A(n_3462),
.B(n_825),
.Y(n_3782)
);

OAI22xp5_ASAP7_75t_L g3783 ( 
.A1(n_3479),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_3783)
);

OAI21x1_ASAP7_75t_L g3784 ( 
.A1(n_3223),
.A2(n_196),
.B(n_197),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3142),
.B(n_197),
.Y(n_3785)
);

OAI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_3354),
.A2(n_198),
.B(n_199),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3414),
.Y(n_3787)
);

A2O1A1Ixp33_ASAP7_75t_L g3788 ( 
.A1(n_3469),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_3788)
);

OAI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_2995),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3416),
.B(n_201),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3418),
.B(n_202),
.Y(n_3791)
);

OAI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3360),
.A2(n_202),
.B(n_203),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_2971),
.A2(n_202),
.B(n_203),
.Y(n_3793)
);

NAND3xp33_ASAP7_75t_L g3794 ( 
.A(n_3423),
.B(n_204),
.C(n_205),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_2909),
.A2(n_204),
.B(n_205),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_2913),
.A2(n_204),
.B(n_205),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3424),
.B(n_206),
.Y(n_3797)
);

A2O1A1Ixp33_ASAP7_75t_L g3798 ( 
.A1(n_3477),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3427),
.B(n_208),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_SL g3800 ( 
.A(n_3212),
.B(n_826),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3430),
.B(n_208),
.Y(n_3801)
);

O2A1O1Ixp33_ASAP7_75t_L g3802 ( 
.A1(n_3011),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_3802)
);

OAI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3369),
.A2(n_209),
.B(n_210),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_SL g3804 ( 
.A(n_3151),
.B(n_827),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_2919),
.A2(n_209),
.B(n_210),
.Y(n_3805)
);

O2A1O1Ixp33_ASAP7_75t_L g3806 ( 
.A1(n_3362),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3435),
.B(n_212),
.Y(n_3807)
);

AND2x4_ASAP7_75t_L g3808 ( 
.A(n_3242),
.B(n_212),
.Y(n_3808)
);

AO21x1_ASAP7_75t_L g3809 ( 
.A1(n_3230),
.A2(n_830),
.B(n_829),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_3093),
.A2(n_213),
.B(n_214),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3096),
.A2(n_2854),
.B(n_2853),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3437),
.B(n_214),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3450),
.Y(n_3813)
);

AOI21x1_ASAP7_75t_L g3814 ( 
.A1(n_3373),
.A2(n_215),
.B(n_216),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_2856),
.A2(n_215),
.B(n_216),
.Y(n_3815)
);

AND2x4_ASAP7_75t_L g3816 ( 
.A(n_3242),
.B(n_3315),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_3451),
.B(n_215),
.Y(n_3817)
);

O2A1O1Ixp33_ASAP7_75t_L g3818 ( 
.A1(n_3366),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_SL g3819 ( 
.A(n_3151),
.B(n_2880),
.Y(n_3819)
);

NOR2xp33_ASAP7_75t_L g3820 ( 
.A(n_3167),
.B(n_3060),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3454),
.B(n_3456),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_L g3822 ( 
.A(n_3460),
.B(n_217),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3461),
.B(n_217),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3465),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_2857),
.A2(n_218),
.B(n_219),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3478),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3484),
.B(n_219),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_L g3828 ( 
.A(n_3290),
.B(n_219),
.Y(n_3828)
);

BUFx2_ASAP7_75t_L g3829 ( 
.A(n_3132),
.Y(n_3829)
);

AOI21xp5_ASAP7_75t_L g3830 ( 
.A1(n_2866),
.A2(n_220),
.B(n_221),
.Y(n_3830)
);

AOI21x1_ASAP7_75t_L g3831 ( 
.A1(n_3381),
.A2(n_220),
.B(n_221),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_2868),
.B(n_221),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_2867),
.A2(n_222),
.B(n_223),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_2872),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_2889),
.Y(n_3835)
);

BUFx6f_ASAP7_75t_L g3836 ( 
.A(n_3274),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_2891),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_2878),
.B(n_222),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_2888),
.B(n_222),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_2831),
.B(n_829),
.Y(n_3840)
);

AOI21xp5_ASAP7_75t_L g3841 ( 
.A1(n_2898),
.A2(n_223),
.B(n_224),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_2901),
.Y(n_3842)
);

HB1xp67_ASAP7_75t_L g3843 ( 
.A(n_3291),
.Y(n_3843)
);

AOI21x1_ASAP7_75t_L g3844 ( 
.A1(n_3389),
.A2(n_224),
.B(n_225),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_2904),
.A2(n_225),
.B(n_226),
.Y(n_3845)
);

AOI21xp5_ASAP7_75t_L g3846 ( 
.A1(n_2906),
.A2(n_226),
.B(n_227),
.Y(n_3846)
);

BUFx4f_ASAP7_75t_L g3847 ( 
.A(n_3398),
.Y(n_3847)
);

AOI21xp5_ASAP7_75t_L g3848 ( 
.A1(n_3399),
.A2(n_226),
.B(n_228),
.Y(n_3848)
);

A2O1A1Ixp33_ASAP7_75t_L g3849 ( 
.A1(n_3401),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_3849)
);

AOI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3403),
.A2(n_228),
.B(n_230),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3307),
.B(n_231),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3035),
.B(n_232),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_2929),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3425),
.A2(n_232),
.B(n_233),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_3314),
.B(n_830),
.Y(n_3855)
);

AOI21xp5_ASAP7_75t_L g3856 ( 
.A1(n_3441),
.A2(n_232),
.B(n_234),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3038),
.B(n_234),
.Y(n_3857)
);

OAI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_2995),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_2985),
.Y(n_3859)
);

CKINVDCx10_ASAP7_75t_R g3860 ( 
.A(n_3312),
.Y(n_3860)
);

AOI21xp5_ASAP7_75t_L g3861 ( 
.A1(n_3442),
.A2(n_235),
.B(n_236),
.Y(n_3861)
);

HB1xp67_ASAP7_75t_L g3862 ( 
.A(n_3336),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_2979),
.Y(n_3863)
);

AOI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_3446),
.A2(n_235),
.B(n_237),
.Y(n_3864)
);

AOI22xp5_ASAP7_75t_L g3865 ( 
.A1(n_2827),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_3865)
);

O2A1O1Ixp5_ASAP7_75t_SL g3866 ( 
.A1(n_3064),
.A2(n_832),
.B(n_833),
.C(n_831),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_2990),
.Y(n_3867)
);

AOI21x1_ASAP7_75t_L g3868 ( 
.A1(n_3215),
.A2(n_238),
.B(n_239),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_2991),
.Y(n_3869)
);

OAI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_2903),
.A2(n_239),
.B(n_240),
.Y(n_3870)
);

AO22x1_ASAP7_75t_L g3871 ( 
.A1(n_3398),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3040),
.B(n_240),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3046),
.B(n_241),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_SL g3874 ( 
.A(n_3342),
.B(n_832),
.Y(n_3874)
);

AOI22xp33_ASAP7_75t_L g3875 ( 
.A1(n_3307),
.A2(n_3335),
.B1(n_3448),
.B2(n_3330),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3049),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3051),
.B(n_242),
.Y(n_3877)
);

AND2x2_ASAP7_75t_L g3878 ( 
.A(n_3330),
.B(n_242),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3053),
.B(n_243),
.Y(n_3879)
);

AOI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3235),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_3880)
);

A2O1A1Ixp33_ASAP7_75t_L g3881 ( 
.A1(n_3012),
.A2(n_246),
.B(n_244),
.C(n_245),
.Y(n_3881)
);

INVx3_ASAP7_75t_L g3882 ( 
.A(n_3342),
.Y(n_3882)
);

O2A1O1Ixp33_ASAP7_75t_SL g3883 ( 
.A1(n_2887),
.A2(n_248),
.B(n_246),
.C(n_247),
.Y(n_3883)
);

AO21x1_ASAP7_75t_L g3884 ( 
.A1(n_3353),
.A2(n_835),
.B(n_833),
.Y(n_3884)
);

A2O1A1Ixp33_ASAP7_75t_L g3885 ( 
.A1(n_3394),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_L g3886 ( 
.A(n_2881),
.B(n_2890),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_2881),
.B(n_248),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_SL g3888 ( 
.A(n_3342),
.B(n_837),
.Y(n_3888)
);

NOR3xp33_ASAP7_75t_L g3889 ( 
.A(n_3045),
.B(n_249),
.C(n_250),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3118),
.A2(n_251),
.B1(n_249),
.B2(n_250),
.Y(n_3890)
);

AOI22xp5_ASAP7_75t_L g3891 ( 
.A1(n_3284),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_3891)
);

OAI21xp5_ASAP7_75t_L g3892 ( 
.A1(n_3103),
.A2(n_252),
.B(n_253),
.Y(n_3892)
);

BUFx6f_ASAP7_75t_L g3893 ( 
.A(n_3467),
.Y(n_3893)
);

AOI21x1_ASAP7_75t_L g3894 ( 
.A1(n_3027),
.A2(n_252),
.B(n_254),
.Y(n_3894)
);

AO21x1_ASAP7_75t_L g3895 ( 
.A1(n_3372),
.A2(n_838),
.B(n_837),
.Y(n_3895)
);

OAI22xp5_ASAP7_75t_L g3896 ( 
.A1(n_3118),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_3896)
);

AOI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3264),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_3897)
);

AOI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_3191),
.A2(n_256),
.B(n_257),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_2890),
.B(n_258),
.Y(n_3899)
);

NOR3xp33_ASAP7_75t_L g3900 ( 
.A(n_3101),
.B(n_259),
.C(n_260),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3192),
.A2(n_259),
.B(n_260),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_2940),
.B(n_259),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3146),
.B(n_260),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3147),
.A2(n_3113),
.B(n_2993),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_2992),
.Y(n_3905)
);

A2O1A1Ixp33_ASAP7_75t_L g3906 ( 
.A1(n_3407),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3128),
.B(n_261),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3130),
.B(n_261),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3145),
.B(n_262),
.Y(n_3909)
);

OAI21xp5_ASAP7_75t_L g3910 ( 
.A1(n_3107),
.A2(n_262),
.B(n_263),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3098),
.B(n_263),
.Y(n_3911)
);

AND2x6_ASAP7_75t_L g3912 ( 
.A(n_3467),
.B(n_264),
.Y(n_3912)
);

OAI21x1_ASAP7_75t_L g3913 ( 
.A1(n_3032),
.A2(n_264),
.B(n_265),
.Y(n_3913)
);

AOI21xp5_ASAP7_75t_L g3914 ( 
.A1(n_2997),
.A2(n_264),
.B(n_265),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_3348),
.B(n_266),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_SL g3916 ( 
.A(n_3467),
.B(n_838),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3015),
.A2(n_266),
.B(n_267),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3404),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3099),
.B(n_267),
.Y(n_3919)
);

AOI21xp5_ASAP7_75t_L g3920 ( 
.A1(n_3034),
.A2(n_267),
.B(n_268),
.Y(n_3920)
);

AOI21xp5_ASAP7_75t_L g3921 ( 
.A1(n_3052),
.A2(n_268),
.B(n_269),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3104),
.B(n_268),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_2976),
.B(n_3324),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3404),
.Y(n_3924)
);

CKINVDCx6p67_ASAP7_75t_R g3925 ( 
.A(n_3480),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3043),
.B(n_2884),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_SL g3927 ( 
.A(n_3166),
.B(n_839),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3068),
.A2(n_269),
.B(n_270),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_2886),
.B(n_270),
.Y(n_3929)
);

A2O1A1Ixp33_ASAP7_75t_L g3930 ( 
.A1(n_3409),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_3930)
);

NOR2xp33_ASAP7_75t_L g3931 ( 
.A(n_3352),
.B(n_272),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3335),
.B(n_272),
.Y(n_3932)
);

BUFx2_ASAP7_75t_L g3933 ( 
.A(n_2859),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3404),
.Y(n_3934)
);

AOI22xp33_ASAP7_75t_L g3935 ( 
.A1(n_3448),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3404),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3249),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_2886),
.B(n_273),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3070),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3071),
.A2(n_273),
.B(n_274),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3249),
.Y(n_3941)
);

AOI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3083),
.A2(n_274),
.B(n_275),
.Y(n_3942)
);

OAI21xp33_ASAP7_75t_L g3943 ( 
.A1(n_2961),
.A2(n_276),
.B(n_277),
.Y(n_3943)
);

A2O1A1Ixp33_ASAP7_75t_L g3944 ( 
.A1(n_3468),
.A2(n_278),
.B(n_276),
.C(n_277),
.Y(n_3944)
);

NOR2xp33_ASAP7_75t_L g3945 ( 
.A(n_3400),
.B(n_276),
.Y(n_3945)
);

INVx2_ASAP7_75t_L g3946 ( 
.A(n_3091),
.Y(n_3946)
);

NAND3xp33_ASAP7_75t_SL g3947 ( 
.A(n_3010),
.B(n_277),
.C(n_278),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_SL g3948 ( 
.A(n_2977),
.B(n_839),
.Y(n_3948)
);

AOI21xp5_ASAP7_75t_L g3949 ( 
.A1(n_3116),
.A2(n_279),
.B(n_280),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3250),
.Y(n_3950)
);

OAI22xp5_ASAP7_75t_L g3951 ( 
.A1(n_3123),
.A2(n_3137),
.B1(n_2961),
.B2(n_3439),
.Y(n_3951)
);

A2O1A1Ixp33_ASAP7_75t_L g3952 ( 
.A1(n_3472),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_3952)
);

AOI21xp5_ASAP7_75t_L g3953 ( 
.A1(n_3117),
.A2(n_280),
.B(n_281),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_3250),
.Y(n_3954)
);

BUFx3_ASAP7_75t_L g3955 ( 
.A(n_3177),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3120),
.A2(n_282),
.B(n_283),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3273),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3160),
.A2(n_283),
.B(n_284),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3029),
.A2(n_284),
.B(n_285),
.Y(n_3959)
);

CKINVDCx20_ASAP7_75t_R g3960 ( 
.A(n_3481),
.Y(n_3960)
);

NAND2xp33_ASAP7_75t_L g3961 ( 
.A(n_3287),
.B(n_285),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_3018),
.A2(n_286),
.B(n_287),
.Y(n_3962)
);

AOI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3023),
.A2(n_286),
.B(n_287),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_2841),
.A2(n_286),
.B(n_287),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_2843),
.A2(n_288),
.B(n_289),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3287),
.Y(n_3966)
);

NOR2x1p5_ASAP7_75t_SL g3967 ( 
.A(n_3190),
.B(n_840),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_2949),
.B(n_288),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3452),
.B(n_288),
.Y(n_3969)
);

NOR2xp33_ASAP7_75t_L g3970 ( 
.A(n_3440),
.B(n_289),
.Y(n_3970)
);

OAI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_2848),
.A2(n_289),
.B(n_290),
.Y(n_3971)
);

NOR2x1_ASAP7_75t_SL g3972 ( 
.A(n_3203),
.B(n_290),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_2865),
.A2(n_291),
.B(n_292),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_2949),
.B(n_292),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_SL g3975 ( 
.A(n_3232),
.B(n_840),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3444),
.B(n_841),
.Y(n_3976)
);

A2O1A1Ixp33_ASAP7_75t_L g3977 ( 
.A1(n_3153),
.A2(n_295),
.B(n_293),
.C(n_294),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_SL g3978 ( 
.A(n_2893),
.B(n_293),
.Y(n_3978)
);

OAI22xp5_ASAP7_75t_L g3979 ( 
.A1(n_3123),
.A2(n_3137),
.B1(n_3470),
.B2(n_3452),
.Y(n_3979)
);

NOR2xp33_ASAP7_75t_L g3980 ( 
.A(n_3476),
.B(n_294),
.Y(n_3980)
);

OAI21xp33_ASAP7_75t_L g3981 ( 
.A1(n_2845),
.A2(n_295),
.B(n_296),
.Y(n_3981)
);

AOI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_2873),
.A2(n_295),
.B(n_296),
.Y(n_3982)
);

CKINVDCx11_ASAP7_75t_R g3983 ( 
.A(n_3338),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_2930),
.B(n_297),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_2875),
.A2(n_297),
.B(n_298),
.Y(n_3985)
);

AOI21xp5_ASAP7_75t_L g3986 ( 
.A1(n_3196),
.A2(n_3028),
.B(n_3026),
.Y(n_3986)
);

AOI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_2987),
.A2(n_2999),
.B(n_3198),
.Y(n_3987)
);

NAND3xp33_ASAP7_75t_L g3988 ( 
.A(n_3102),
.B(n_297),
.C(n_298),
.Y(n_3988)
);

AOI21xp5_ASAP7_75t_L g3989 ( 
.A1(n_3199),
.A2(n_298),
.B(n_299),
.Y(n_3989)
);

OAI21x1_ASAP7_75t_L g3990 ( 
.A1(n_3092),
.A2(n_299),
.B(n_300),
.Y(n_3990)
);

A2O1A1Ixp33_ASAP7_75t_L g3991 ( 
.A1(n_3334),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_3991)
);

A2O1A1Ixp33_ASAP7_75t_L g3992 ( 
.A1(n_3150),
.A2(n_3200),
.B(n_2836),
.C(n_2855),
.Y(n_3992)
);

AOI21x1_ASAP7_75t_L g3993 ( 
.A1(n_3066),
.A2(n_2874),
.B(n_2850),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3141),
.B(n_300),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_SL g3995 ( 
.A(n_2981),
.B(n_842),
.Y(n_3995)
);

AOI21xp5_ASAP7_75t_L g3996 ( 
.A1(n_3185),
.A2(n_301),
.B(n_303),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3273),
.Y(n_3997)
);

HB1xp67_ASAP7_75t_L g3998 ( 
.A(n_3152),
.Y(n_3998)
);

NAND3xp33_ASAP7_75t_L g3999 ( 
.A(n_3163),
.B(n_3231),
.C(n_3162),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_L g4000 ( 
.A(n_2836),
.B(n_301),
.Y(n_4000)
);

AO32x1_ASAP7_75t_L g4001 ( 
.A1(n_3136),
.A2(n_305),
.A3(n_303),
.B1(n_304),
.B2(n_306),
.Y(n_4001)
);

AOI21xp33_ASAP7_75t_L g4002 ( 
.A1(n_3139),
.A2(n_3172),
.B(n_3059),
.Y(n_4002)
);

AOI22x1_ASAP7_75t_L g4003 ( 
.A1(n_3095),
.A2(n_306),
.B1(n_303),
.B2(n_305),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3287),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_2981),
.B(n_843),
.Y(n_4005)
);

AOI21x1_ASAP7_75t_L g4006 ( 
.A1(n_2850),
.A2(n_305),
.B(n_306),
.Y(n_4006)
);

AOI21x1_ASAP7_75t_L g4007 ( 
.A1(n_2874),
.A2(n_307),
.B(n_308),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_L g4008 ( 
.A(n_3378),
.B(n_307),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_2844),
.B(n_307),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_L g4010 ( 
.A(n_3390),
.B(n_308),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_2844),
.B(n_309),
.Y(n_4011)
);

A2O1A1Ixp33_ASAP7_75t_L g4012 ( 
.A1(n_2855),
.A2(n_311),
.B(n_309),
.C(n_310),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3309),
.A2(n_309),
.B(n_311),
.Y(n_4013)
);

AOI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_2908),
.A2(n_311),
.B(n_312),
.Y(n_4014)
);

A2O1A1Ixp33_ASAP7_75t_L g4015 ( 
.A1(n_2863),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_4015)
);

INVx2_ASAP7_75t_L g4016 ( 
.A(n_3287),
.Y(n_4016)
);

A2O1A1Ixp33_ASAP7_75t_L g4017 ( 
.A1(n_2863),
.A2(n_314),
.B(n_312),
.C(n_313),
.Y(n_4017)
);

CKINVDCx11_ASAP7_75t_R g4018 ( 
.A(n_3155),
.Y(n_4018)
);

OAI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_3470),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3054),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3346),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_2833),
.B(n_315),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_2833),
.B(n_315),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_2847),
.B(n_316),
.Y(n_4024)
);

OAI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_3081),
.A2(n_317),
.B(n_318),
.Y(n_4025)
);

AOI21xp5_ASAP7_75t_L g4026 ( 
.A1(n_3246),
.A2(n_317),
.B(n_318),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_3259),
.A2(n_319),
.B(n_320),
.Y(n_4027)
);

NOR2xp67_ASAP7_75t_L g4028 ( 
.A(n_2926),
.B(n_319),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3361),
.B(n_319),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_2998),
.B(n_320),
.Y(n_4030)
);

CKINVDCx10_ASAP7_75t_R g4031 ( 
.A(n_3481),
.Y(n_4031)
);

AND2x2_ASAP7_75t_SL g4032 ( 
.A(n_3308),
.B(n_320),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3365),
.B(n_321),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3382),
.Y(n_4034)
);

AOI21xp5_ASAP7_75t_L g4035 ( 
.A1(n_3277),
.A2(n_321),
.B(n_322),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3384),
.Y(n_4036)
);

O2A1O1Ixp33_ASAP7_75t_L g4037 ( 
.A1(n_3240),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3396),
.B(n_322),
.Y(n_4038)
);

AOI21xp5_ASAP7_75t_L g4039 ( 
.A1(n_3304),
.A2(n_3332),
.B(n_3181),
.Y(n_4039)
);

AOI21xp5_ASAP7_75t_L g4040 ( 
.A1(n_3209),
.A2(n_3211),
.B(n_3126),
.Y(n_4040)
);

AOI21x1_ASAP7_75t_L g4041 ( 
.A1(n_3179),
.A2(n_323),
.B(n_325),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3443),
.B(n_325),
.Y(n_4042)
);

AOI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_3114),
.A2(n_3055),
.B(n_3075),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_2910),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3445),
.B(n_325),
.Y(n_4045)
);

INVx3_ASAP7_75t_L g4046 ( 
.A(n_3315),
.Y(n_4046)
);

NOR3xp33_ASAP7_75t_L g4047 ( 
.A(n_3122),
.B(n_326),
.C(n_327),
.Y(n_4047)
);

BUFx4f_ASAP7_75t_L g4048 ( 
.A(n_3397),
.Y(n_4048)
);

NOR2xp33_ASAP7_75t_L g4049 ( 
.A(n_3058),
.B(n_326),
.Y(n_4049)
);

OAI21x1_ASAP7_75t_L g4050 ( 
.A1(n_2942),
.A2(n_327),
.B(n_328),
.Y(n_4050)
);

AOI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_2947),
.A2(n_327),
.B(n_328),
.Y(n_4051)
);

NOR2x1_ASAP7_75t_L g4052 ( 
.A(n_3189),
.B(n_329),
.Y(n_4052)
);

AOI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_3061),
.A2(n_329),
.B(n_330),
.Y(n_4053)
);

OAI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3174),
.A2(n_329),
.B(n_330),
.Y(n_4054)
);

OAI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3072),
.A2(n_331),
.B(n_332),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3039),
.B(n_844),
.Y(n_4056)
);

OAI21xp33_ASAP7_75t_L g4057 ( 
.A1(n_3024),
.A2(n_331),
.B(n_332),
.Y(n_4057)
);

AOI21xp5_ASAP7_75t_L g4058 ( 
.A1(n_3062),
.A2(n_331),
.B(n_332),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3670),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_SL g4060 ( 
.A(n_3536),
.B(n_3406),
.Y(n_4060)
);

NAND3xp33_ASAP7_75t_SL g4061 ( 
.A(n_3978),
.B(n_3415),
.C(n_3457),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3509),
.Y(n_4062)
);

OAI22xp5_ASAP7_75t_L g4063 ( 
.A1(n_3536),
.A2(n_3024),
.B1(n_2870),
.B2(n_3003),
.Y(n_4063)
);

A2O1A1Ixp33_ASAP7_75t_L g4064 ( 
.A1(n_3847),
.A2(n_3162),
.B(n_3463),
.C(n_3039),
.Y(n_4064)
);

OR2x6_ASAP7_75t_SL g4065 ( 
.A(n_3712),
.B(n_3044),
.Y(n_4065)
);

HB1xp67_ASAP7_75t_L g4066 ( 
.A(n_3604),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3535),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3719),
.B(n_3156),
.Y(n_4068)
);

AOI21xp5_ASAP7_75t_L g4069 ( 
.A1(n_3847),
.A2(n_3179),
.B(n_3156),
.Y(n_4069)
);

OAI22xp5_ASAP7_75t_L g4070 ( 
.A1(n_3875),
.A2(n_3485),
.B1(n_2869),
.B2(n_2842),
.Y(n_4070)
);

A2O1A1Ixp33_ASAP7_75t_L g4071 ( 
.A1(n_3710),
.A2(n_3121),
.B(n_3187),
.C(n_2956),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3719),
.B(n_3042),
.Y(n_4072)
);

INVx3_ASAP7_75t_L g4073 ( 
.A(n_3614),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_SL g4074 ( 
.A(n_3979),
.B(n_3227),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3685),
.Y(n_4075)
);

NOR2xp33_ASAP7_75t_L g4076 ( 
.A(n_3575),
.B(n_2928),
.Y(n_4076)
);

AOI21x1_ASAP7_75t_SL g4077 ( 
.A1(n_4030),
.A2(n_3187),
.B(n_3063),
.Y(n_4077)
);

AOI21xp5_ASAP7_75t_L g4078 ( 
.A1(n_3961),
.A2(n_3041),
.B(n_3180),
.Y(n_4078)
);

HB1xp67_ASAP7_75t_L g4079 ( 
.A(n_3603),
.Y(n_4079)
);

NOR2xp33_ASAP7_75t_L g4080 ( 
.A(n_3649),
.B(n_2907),
.Y(n_4080)
);

AOI21xp5_ASAP7_75t_L g4081 ( 
.A1(n_3503),
.A2(n_3183),
.B(n_3182),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3719),
.B(n_3545),
.Y(n_4082)
);

AOI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_3527),
.A2(n_3184),
.B(n_3144),
.Y(n_4083)
);

OAI22xp5_ASAP7_75t_L g4084 ( 
.A1(n_3703),
.A2(n_3951),
.B1(n_3690),
.B2(n_4032),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_3550),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3719),
.B(n_3042),
.Y(n_4086)
);

AOI22xp33_ASAP7_75t_L g4087 ( 
.A1(n_3605),
.A2(n_3086),
.B1(n_3063),
.B2(n_3079),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_SL g4088 ( 
.A(n_4048),
.B(n_3057),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3698),
.Y(n_4089)
);

A2O1A1Ixp33_ASAP7_75t_L g4090 ( 
.A1(n_3755),
.A2(n_3121),
.B(n_2956),
.C(n_2955),
.Y(n_4090)
);

NOR2xp33_ASAP7_75t_L g4091 ( 
.A(n_3721),
.B(n_2972),
.Y(n_4091)
);

NOR2xp33_ASAP7_75t_L g4092 ( 
.A(n_3752),
.B(n_2922),
.Y(n_4092)
);

NOR2xp67_ASAP7_75t_SL g4093 ( 
.A(n_3754),
.B(n_3090),
.Y(n_4093)
);

OAI22xp5_ASAP7_75t_L g4094 ( 
.A1(n_3777),
.A2(n_3097),
.B1(n_3195),
.B2(n_3086),
.Y(n_4094)
);

HB1xp67_ASAP7_75t_L g4095 ( 
.A(n_3487),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3531),
.B(n_3089),
.Y(n_4096)
);

NOR2xp33_ASAP7_75t_L g4097 ( 
.A(n_3999),
.B(n_2954),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3564),
.B(n_3331),
.Y(n_4098)
);

O2A1O1Ixp33_ASAP7_75t_L g4099 ( 
.A1(n_3992),
.A2(n_3220),
.B(n_3002),
.C(n_3248),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_SL g4100 ( 
.A(n_4048),
.B(n_3057),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_3732),
.Y(n_4101)
);

OAI22xp5_ASAP7_75t_L g4102 ( 
.A1(n_3780),
.A2(n_3078),
.B1(n_3100),
.B2(n_2840),
.Y(n_4102)
);

AOI21xp5_ASAP7_75t_L g4103 ( 
.A1(n_3488),
.A2(n_3143),
.B(n_3206),
.Y(n_4103)
);

AOI21xp5_ASAP7_75t_L g4104 ( 
.A1(n_3547),
.A2(n_3216),
.B(n_3100),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_3706),
.B(n_3319),
.Y(n_4105)
);

AOI22xp5_ASAP7_75t_L g4106 ( 
.A1(n_3947),
.A2(n_3178),
.B1(n_3218),
.B2(n_2955),
.Y(n_4106)
);

AO32x1_ASAP7_75t_L g4107 ( 
.A1(n_3522),
.A2(n_3266),
.A3(n_3464),
.B1(n_3343),
.B2(n_3317),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_3741),
.Y(n_4108)
);

OR2x2_ASAP7_75t_L g4109 ( 
.A(n_3886),
.B(n_3319),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_3987),
.A2(n_3022),
.B(n_3217),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_3716),
.B(n_3447),
.Y(n_4111)
);

AND2x2_ASAP7_75t_L g4112 ( 
.A(n_3726),
.B(n_3447),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3508),
.B(n_3154),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_3986),
.A2(n_3022),
.B(n_3219),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3543),
.B(n_3079),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_3744),
.Y(n_4116)
);

A2O1A1Ixp33_ASAP7_75t_L g4117 ( 
.A1(n_3802),
.A2(n_3466),
.B(n_3135),
.C(n_3033),
.Y(n_4117)
);

AND2x4_ASAP7_75t_L g4118 ( 
.A(n_3918),
.B(n_3466),
.Y(n_4118)
);

INVx5_ASAP7_75t_L g4119 ( 
.A(n_3912),
.Y(n_4119)
);

O2A1O1Ixp33_ASAP7_75t_L g4120 ( 
.A1(n_3624),
.A2(n_3020),
.B(n_3222),
.C(n_3221),
.Y(n_4120)
);

BUFx12f_ASAP7_75t_L g4121 ( 
.A(n_3505),
.Y(n_4121)
);

AOI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_3687),
.A2(n_3226),
.B(n_3171),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3674),
.B(n_3140),
.Y(n_4123)
);

NAND3xp33_ASAP7_75t_SL g4124 ( 
.A(n_3611),
.B(n_3311),
.C(n_3241),
.Y(n_4124)
);

OR2x2_ASAP7_75t_L g4125 ( 
.A(n_3684),
.B(n_3082),
.Y(n_4125)
);

O2A1O1Ixp33_ASAP7_75t_SL g4126 ( 
.A1(n_4012),
.A2(n_3482),
.B(n_3251),
.C(n_3009),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3584),
.B(n_2978),
.Y(n_4127)
);

INVx2_ASAP7_75t_SL g4128 ( 
.A(n_3829),
.Y(n_4128)
);

CKINVDCx16_ASAP7_75t_R g4129 ( 
.A(n_3653),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_3626),
.B(n_3047),
.Y(n_4130)
);

NOR2xp33_ASAP7_75t_L g4131 ( 
.A(n_3923),
.B(n_3194),
.Y(n_4131)
);

AOI21xp5_ASAP7_75t_L g4132 ( 
.A1(n_3762),
.A2(n_3175),
.B(n_3170),
.Y(n_4132)
);

OAI21xp33_ASAP7_75t_L g4133 ( 
.A1(n_4057),
.A2(n_3943),
.B(n_3935),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_4028),
.B(n_3085),
.Y(n_4134)
);

AO32x2_ASAP7_75t_L g4135 ( 
.A1(n_3529),
.A2(n_3205),
.A3(n_2960),
.B1(n_335),
.B2(n_333),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_SL g4136 ( 
.A(n_3520),
.B(n_3173),
.Y(n_4136)
);

NOR2xp33_ASAP7_75t_L g4137 ( 
.A(n_3518),
.B(n_3213),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_3766),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3676),
.B(n_3036),
.Y(n_4139)
);

AOI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_3515),
.A2(n_3224),
.B(n_3257),
.Y(n_4140)
);

OA22x2_ASAP7_75t_L g4141 ( 
.A1(n_3574),
.A2(n_3109),
.B1(n_2975),
.B2(n_3124),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_3813),
.Y(n_4142)
);

AOI22xp5_ASAP7_75t_L g4143 ( 
.A1(n_3520),
.A2(n_3017),
.B1(n_3112),
.B2(n_3127),
.Y(n_4143)
);

INVx3_ASAP7_75t_L g4144 ( 
.A(n_3617),
.Y(n_4144)
);

NOR3xp33_ASAP7_75t_SL g4145 ( 
.A(n_4019),
.B(n_3149),
.C(n_3125),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3677),
.B(n_3261),
.Y(n_4146)
);

BUFx2_ASAP7_75t_L g4147 ( 
.A(n_3617),
.Y(n_4147)
);

AOI21xp5_ASAP7_75t_L g4148 ( 
.A1(n_3904),
.A2(n_3644),
.B(n_3631),
.Y(n_4148)
);

OAI22xp5_ASAP7_75t_L g4149 ( 
.A1(n_3632),
.A2(n_3620),
.B1(n_3675),
.B2(n_3573),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_3724),
.B(n_3368),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_3824),
.Y(n_4151)
);

BUFx3_ASAP7_75t_L g4152 ( 
.A(n_3634),
.Y(n_4152)
);

OAI21x1_ASAP7_75t_SL g4153 ( 
.A1(n_4041),
.A2(n_333),
.B(n_334),
.Y(n_4153)
);

AOI22xp33_ASAP7_75t_L g4154 ( 
.A1(n_3699),
.A2(n_3094),
.B1(n_3202),
.B2(n_3204),
.Y(n_4154)
);

NOR2x1_ASAP7_75t_L g4155 ( 
.A(n_4052),
.B(n_3094),
.Y(n_4155)
);

AOI21xp5_ASAP7_75t_L g4156 ( 
.A1(n_3811),
.A2(n_333),
.B(n_334),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3523),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3727),
.B(n_334),
.Y(n_4158)
);

INVx6_ASAP7_75t_L g4159 ( 
.A(n_3636),
.Y(n_4159)
);

AND2x4_ASAP7_75t_L g4160 ( 
.A(n_3924),
.B(n_335),
.Y(n_4160)
);

OAI22xp5_ASAP7_75t_L g4161 ( 
.A1(n_3632),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_4161)
);

AOI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_3794),
.A2(n_336),
.B(n_337),
.Y(n_4162)
);

AOI22xp33_ASAP7_75t_L g4163 ( 
.A1(n_3489),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3837),
.Y(n_4164)
);

AOI22xp5_ASAP7_75t_L g4165 ( 
.A1(n_3820),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_4165)
);

BUFx6f_ASAP7_75t_L g4166 ( 
.A(n_3499),
.Y(n_4166)
);

NAND2x1p5_ASAP7_75t_L g4167 ( 
.A(n_3955),
.B(n_338),
.Y(n_4167)
);

NAND3xp33_ASAP7_75t_L g4168 ( 
.A(n_3866),
.B(n_339),
.C(n_340),
.Y(n_4168)
);

NAND2xp33_ASAP7_75t_L g4169 ( 
.A(n_3912),
.B(n_3519),
.Y(n_4169)
);

AOI21xp5_ASAP7_75t_L g4170 ( 
.A1(n_4039),
.A2(n_340),
.B(n_341),
.Y(n_4170)
);

A2O1A1Ixp33_ASAP7_75t_L g4171 ( 
.A1(n_4054),
.A2(n_4055),
.B(n_3666),
.C(n_4037),
.Y(n_4171)
);

OAI22xp5_ASAP7_75t_L g4172 ( 
.A1(n_3630),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_4172)
);

A2O1A1Ixp33_ASAP7_75t_L g4173 ( 
.A1(n_3981),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_4173)
);

AOI21xp5_ASAP7_75t_L g4174 ( 
.A1(n_3580),
.A2(n_342),
.B(n_343),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_3761),
.B(n_344),
.Y(n_4175)
);

AOI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_3934),
.A2(n_344),
.B(n_345),
.Y(n_4176)
);

INVx8_ASAP7_75t_L g4177 ( 
.A(n_3693),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3876),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3863),
.Y(n_4179)
);

NAND2x1p5_ASAP7_75t_L g4180 ( 
.A(n_3551),
.B(n_345),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_3772),
.B(n_345),
.Y(n_4181)
);

BUFx6f_ASAP7_75t_L g4182 ( 
.A(n_3499),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_L g4183 ( 
.A(n_3774),
.B(n_346),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_SL g4184 ( 
.A(n_3549),
.B(n_347),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3787),
.B(n_347),
.Y(n_4185)
);

O2A1O1Ixp33_ASAP7_75t_L g4186 ( 
.A1(n_3635),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_4186)
);

OAI21x1_ASAP7_75t_L g4187 ( 
.A1(n_3561),
.A2(n_350),
.B(n_349),
.Y(n_4187)
);

NOR2xp33_ASAP7_75t_L g4188 ( 
.A(n_3933),
.B(n_348),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_R g4189 ( 
.A(n_3960),
.B(n_350),
.Y(n_4189)
);

INVx6_ASAP7_75t_L g4190 ( 
.A(n_3636),
.Y(n_4190)
);

O2A1O1Ixp33_ASAP7_75t_L g4191 ( 
.A1(n_3495),
.A2(n_353),
.B(n_351),
.C(n_352),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_3826),
.B(n_351),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_SL g4193 ( 
.A(n_3504),
.B(n_352),
.Y(n_4193)
);

BUFx2_ASAP7_75t_L g4194 ( 
.A(n_3669),
.Y(n_4194)
);

AOI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_3936),
.A2(n_4043),
.B(n_3819),
.Y(n_4195)
);

OAI22xp5_ASAP7_75t_L g4196 ( 
.A1(n_3758),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_3842),
.Y(n_4197)
);

NAND2x1p5_ASAP7_75t_L g4198 ( 
.A(n_3738),
.B(n_354),
.Y(n_4198)
);

NOR2xp33_ASAP7_75t_L g4199 ( 
.A(n_3618),
.B(n_3926),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_3834),
.B(n_3835),
.Y(n_4200)
);

INVx4_ASAP7_75t_L g4201 ( 
.A(n_3491),
.Y(n_4201)
);

INVx3_ASAP7_75t_L g4202 ( 
.A(n_3500),
.Y(n_4202)
);

O2A1O1Ixp5_ASAP7_75t_SL g4203 ( 
.A1(n_3948),
.A2(n_847),
.B(n_848),
.C(n_846),
.Y(n_4203)
);

A2O1A1Ixp33_ASAP7_75t_L g4204 ( 
.A1(n_3492),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_4204)
);

NAND3xp33_ASAP7_75t_SL g4205 ( 
.A(n_4047),
.B(n_3730),
.C(n_3897),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_3853),
.B(n_3572),
.Y(n_4206)
);

CKINVDCx6p67_ASAP7_75t_R g4207 ( 
.A(n_3860),
.Y(n_4207)
);

BUFx12f_ASAP7_75t_L g4208 ( 
.A(n_4018),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3601),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_SL g4210 ( 
.A(n_3966),
.B(n_356),
.Y(n_4210)
);

NOR3xp33_ASAP7_75t_SL g4211 ( 
.A(n_3771),
.B(n_3700),
.C(n_3789),
.Y(n_4211)
);

O2A1O1Ixp5_ASAP7_75t_L g4212 ( 
.A1(n_3621),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_4004),
.B(n_357),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_3859),
.Y(n_4214)
);

HB1xp67_ASAP7_75t_L g4215 ( 
.A(n_3998),
.Y(n_4215)
);

INVx2_ASAP7_75t_L g4216 ( 
.A(n_3867),
.Y(n_4216)
);

AOI21xp5_ASAP7_75t_L g4217 ( 
.A1(n_3646),
.A2(n_357),
.B(n_358),
.Y(n_4217)
);

INVx3_ASAP7_75t_L g4218 ( 
.A(n_3500),
.Y(n_4218)
);

NOR2xp33_ASAP7_75t_L g4219 ( 
.A(n_3907),
.B(n_359),
.Y(n_4219)
);

A2O1A1Ixp33_ASAP7_75t_L g4220 ( 
.A1(n_3728),
.A2(n_361),
.B(n_359),
.C(n_360),
.Y(n_4220)
);

NAND2xp33_ASAP7_75t_SL g4221 ( 
.A(n_3750),
.B(n_360),
.Y(n_4221)
);

AOI21xp5_ASAP7_75t_L g4222 ( 
.A1(n_3671),
.A2(n_360),
.B(n_361),
.Y(n_4222)
);

AND2x2_ASAP7_75t_L g4223 ( 
.A(n_3851),
.B(n_362),
.Y(n_4223)
);

A2O1A1Ixp33_ASAP7_75t_L g4224 ( 
.A1(n_3493),
.A2(n_364),
.B(n_362),
.C(n_363),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_SL g4225 ( 
.A(n_4016),
.B(n_362),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_SL g4226 ( 
.A(n_3993),
.B(n_363),
.Y(n_4226)
);

NOR2xp33_ASAP7_75t_L g4227 ( 
.A(n_3983),
.B(n_3709),
.Y(n_4227)
);

BUFx3_ASAP7_75t_L g4228 ( 
.A(n_3925),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3821),
.Y(n_4229)
);

NOR2xp33_ASAP7_75t_L g4230 ( 
.A(n_3843),
.B(n_363),
.Y(n_4230)
);

AOI21xp5_ASAP7_75t_L g4231 ( 
.A1(n_3840),
.A2(n_364),
.B(n_365),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_L g4232 ( 
.A(n_3862),
.B(n_364),
.Y(n_4232)
);

NOR3xp33_ASAP7_75t_SL g4233 ( 
.A(n_3858),
.B(n_365),
.C(n_366),
.Y(n_4233)
);

OAI221xp5_ASAP7_75t_L g4234 ( 
.A1(n_3889),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.C(n_368),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4021),
.B(n_367),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_3855),
.A2(n_368),
.B(n_369),
.Y(n_4236)
);

O2A1O1Ixp33_ASAP7_75t_SL g4237 ( 
.A1(n_4015),
.A2(n_370),
.B(n_368),
.C(n_369),
.Y(n_4237)
);

O2A1O1Ixp33_ASAP7_75t_SL g4238 ( 
.A1(n_4017),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_3869),
.Y(n_4239)
);

INVx4_ASAP7_75t_L g4240 ( 
.A(n_3912),
.Y(n_4240)
);

NAND3xp33_ASAP7_75t_L g4241 ( 
.A(n_3900),
.B(n_370),
.C(n_371),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_3502),
.A2(n_372),
.B(n_373),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_3742),
.A2(n_372),
.B(n_373),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_3506),
.B(n_372),
.Y(n_4244)
);

AOI21xp5_ASAP7_75t_L g4245 ( 
.A1(n_3874),
.A2(n_374),
.B(n_375),
.Y(n_4245)
);

INVx2_ASAP7_75t_SL g4246 ( 
.A(n_4031),
.Y(n_4246)
);

NOR2xp33_ASAP7_75t_R g4247 ( 
.A(n_3497),
.B(n_374),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4034),
.B(n_374),
.Y(n_4248)
);

OAI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_3988),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_4249)
);

AOI221xp5_ASAP7_75t_L g4250 ( 
.A1(n_3616),
.A2(n_379),
.B1(n_376),
.B2(n_378),
.C(n_381),
.Y(n_4250)
);

BUFx6f_ASAP7_75t_L g4251 ( 
.A(n_3499),
.Y(n_4251)
);

HB1xp67_ASAP7_75t_L g4252 ( 
.A(n_3656),
.Y(n_4252)
);

AOI21xp5_ASAP7_75t_L g4253 ( 
.A1(n_3888),
.A2(n_378),
.B(n_379),
.Y(n_4253)
);

BUFx2_ASAP7_75t_L g4254 ( 
.A(n_3669),
.Y(n_4254)
);

O2A1O1Ixp33_ASAP7_75t_L g4255 ( 
.A1(n_3885),
.A2(n_381),
.B(n_378),
.C(n_379),
.Y(n_4255)
);

AOI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_3916),
.A2(n_381),
.B(n_382),
.Y(n_4256)
);

BUFx2_ASAP7_75t_L g4257 ( 
.A(n_3747),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_4020),
.A2(n_382),
.B(n_383),
.Y(n_4258)
);

O2A1O1Ixp33_ASAP7_75t_L g4259 ( 
.A1(n_3906),
.A2(n_385),
.B(n_383),
.C(n_384),
.Y(n_4259)
);

NOR2xp33_ASAP7_75t_L g4260 ( 
.A(n_4036),
.B(n_383),
.Y(n_4260)
);

OAI22xp5_ASAP7_75t_L g4261 ( 
.A1(n_3865),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_4261)
);

O2A1O1Ixp33_ASAP7_75t_L g4262 ( 
.A1(n_3930),
.A2(n_386),
.B(n_384),
.C(n_385),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_3556),
.B(n_386),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_3905),
.Y(n_4264)
);

O2A1O1Ixp33_ASAP7_75t_L g4265 ( 
.A1(n_3944),
.A2(n_390),
.B(n_387),
.C(n_389),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_4044),
.A2(n_387),
.B(n_389),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_3490),
.B(n_387),
.Y(n_4267)
);

A2O1A1Ixp33_ASAP7_75t_L g4268 ( 
.A1(n_3696),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_4268)
);

AND2x4_ASAP7_75t_L g4269 ( 
.A(n_3734),
.B(n_391),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_3507),
.Y(n_4270)
);

AO31x2_ASAP7_75t_L g4271 ( 
.A1(n_3681),
.A2(n_393),
.A3(n_391),
.B(n_392),
.Y(n_4271)
);

CKINVDCx5p33_ASAP7_75t_R g4272 ( 
.A(n_3645),
.Y(n_4272)
);

OAI21xp33_ASAP7_75t_L g4273 ( 
.A1(n_3552),
.A2(n_392),
.B(n_393),
.Y(n_4273)
);

NOR2xp67_ASAP7_75t_SL g4274 ( 
.A(n_3747),
.B(n_394),
.Y(n_4274)
);

HB1xp67_ASAP7_75t_L g4275 ( 
.A(n_3656),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3909),
.Y(n_4276)
);

AOI222xp33_ASAP7_75t_L g4277 ( 
.A1(n_3878),
.A2(n_419),
.B1(n_402),
.B2(n_428),
.C1(n_410),
.C2(n_394),
.Y(n_4277)
);

AOI21xp5_ASAP7_75t_L g4278 ( 
.A1(n_3537),
.A2(n_394),
.B(n_395),
.Y(n_4278)
);

OAI22xp5_ASAP7_75t_L g4279 ( 
.A1(n_3890),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_4279)
);

AND2x2_ASAP7_75t_L g4280 ( 
.A(n_3932),
.B(n_396),
.Y(n_4280)
);

INVx4_ASAP7_75t_L g4281 ( 
.A(n_3912),
.Y(n_4281)
);

INVx3_ASAP7_75t_SL g4282 ( 
.A(n_3722),
.Y(n_4282)
);

BUFx2_ASAP7_75t_SL g4283 ( 
.A(n_3651),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3852),
.Y(n_4284)
);

O2A1O1Ixp33_ASAP7_75t_L g4285 ( 
.A1(n_3952),
.A2(n_399),
.B(n_397),
.C(n_398),
.Y(n_4285)
);

A2O1A1Ixp33_ASAP7_75t_L g4286 ( 
.A1(n_3717),
.A2(n_401),
.B(n_399),
.C(n_400),
.Y(n_4286)
);

NOR2xp33_ASAP7_75t_L g4287 ( 
.A(n_3770),
.B(n_3804),
.Y(n_4287)
);

OAI22xp5_ASAP7_75t_SL g4288 ( 
.A1(n_4008),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_4288)
);

INVx2_ASAP7_75t_L g4289 ( 
.A(n_3546),
.Y(n_4289)
);

BUFx2_ASAP7_75t_L g4290 ( 
.A(n_3519),
.Y(n_4290)
);

INVxp67_ASAP7_75t_SL g4291 ( 
.A(n_3501),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_3559),
.B(n_400),
.Y(n_4292)
);

BUFx6f_ASAP7_75t_L g4293 ( 
.A(n_3501),
.Y(n_4293)
);

O2A1O1Ixp33_ASAP7_75t_L g4294 ( 
.A1(n_3899),
.A2(n_403),
.B(n_401),
.C(n_402),
.Y(n_4294)
);

NOR2xp33_ASAP7_75t_L g4295 ( 
.A(n_3832),
.B(n_403),
.Y(n_4295)
);

INVx2_ASAP7_75t_L g4296 ( 
.A(n_3562),
.Y(n_4296)
);

BUFx8_ASAP7_75t_L g4297 ( 
.A(n_3969),
.Y(n_4297)
);

AOI21xp5_ASAP7_75t_L g4298 ( 
.A1(n_3563),
.A2(n_403),
.B(n_404),
.Y(n_4298)
);

AOI21xp5_ASAP7_75t_L g4299 ( 
.A1(n_3595),
.A2(n_404),
.B(n_405),
.Y(n_4299)
);

OR2x6_ASAP7_75t_L g4300 ( 
.A(n_3722),
.B(n_404),
.Y(n_4300)
);

AOI21xp5_ASAP7_75t_L g4301 ( 
.A1(n_3622),
.A2(n_405),
.B(n_406),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_3857),
.Y(n_4302)
);

INVxp67_ASAP7_75t_SL g4303 ( 
.A(n_3501),
.Y(n_4303)
);

O2A1O1Ixp33_ASAP7_75t_L g4304 ( 
.A1(n_3977),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_4304)
);

INVx2_ASAP7_75t_L g4305 ( 
.A(n_3628),
.Y(n_4305)
);

NOR2xp33_ASAP7_75t_L g4306 ( 
.A(n_3838),
.B(n_408),
.Y(n_4306)
);

OAI21xp33_ASAP7_75t_SL g4307 ( 
.A1(n_3784),
.A2(n_3990),
.B(n_3737),
.Y(n_4307)
);

OR2x6_ASAP7_75t_L g4308 ( 
.A(n_3599),
.B(n_408),
.Y(n_4308)
);

AOI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_3652),
.A2(n_408),
.B(n_409),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_3633),
.B(n_409),
.Y(n_4310)
);

NOR2x1_ASAP7_75t_L g4311 ( 
.A(n_3639),
.B(n_409),
.Y(n_4311)
);

OR2x6_ASAP7_75t_L g4312 ( 
.A(n_3871),
.B(n_410),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_3665),
.Y(n_4313)
);

OAI22xp33_ASAP7_75t_L g4314 ( 
.A1(n_4022),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_4314)
);

AOI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_3672),
.A2(n_411),
.B(n_412),
.Y(n_4315)
);

INVx2_ASAP7_75t_L g4316 ( 
.A(n_3913),
.Y(n_4316)
);

AOI21xp5_ASAP7_75t_L g4317 ( 
.A1(n_3786),
.A2(n_412),
.B(n_413),
.Y(n_4317)
);

NOR2xp33_ASAP7_75t_L g4318 ( 
.A(n_3839),
.B(n_413),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_3637),
.B(n_413),
.Y(n_4319)
);

BUFx8_ASAP7_75t_L g4320 ( 
.A(n_3519),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_3663),
.B(n_414),
.Y(n_4321)
);

O2A1O1Ixp33_ASAP7_75t_L g4322 ( 
.A1(n_3702),
.A2(n_417),
.B(n_414),
.C(n_415),
.Y(n_4322)
);

OAI22xp5_ASAP7_75t_L g4323 ( 
.A1(n_3896),
.A2(n_419),
.B1(n_415),
.B2(n_418),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_3872),
.Y(n_4324)
);

OAI22xp5_ASAP7_75t_SL g4325 ( 
.A1(n_4010),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_SL g4326 ( 
.A(n_3511),
.B(n_420),
.Y(n_4326)
);

A2O1A1Ixp33_ASAP7_75t_SL g4327 ( 
.A1(n_3892),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_4327)
);

CKINVDCx14_ASAP7_75t_R g4328 ( 
.A(n_3519),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_SL g4329 ( 
.A(n_3511),
.B(n_421),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_3733),
.B(n_421),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_SL g4331 ( 
.A(n_3511),
.B(n_422),
.Y(n_4331)
);

OAI22xp5_ASAP7_75t_L g4332 ( 
.A1(n_3714),
.A2(n_425),
.B1(n_423),
.B2(n_424),
.Y(n_4332)
);

O2A1O1Ixp5_ASAP7_75t_L g4333 ( 
.A1(n_3910),
.A2(n_425),
.B(n_423),
.C(n_424),
.Y(n_4333)
);

A2O1A1Ixp33_ASAP7_75t_L g4334 ( 
.A1(n_3971),
.A2(n_426),
.B(n_424),
.C(n_425),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_3510),
.B(n_426),
.Y(n_4335)
);

NOR2xp33_ASAP7_75t_L g4336 ( 
.A(n_4002),
.B(n_426),
.Y(n_4336)
);

AOI21xp5_ASAP7_75t_L g4337 ( 
.A1(n_3792),
.A2(n_428),
.B(n_429),
.Y(n_4337)
);

OR2x6_ASAP7_75t_SL g4338 ( 
.A(n_3707),
.B(n_3713),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_3514),
.B(n_3517),
.Y(n_4339)
);

O2A1O1Ixp33_ASAP7_75t_L g4340 ( 
.A1(n_3740),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_3521),
.B(n_430),
.Y(n_4341)
);

BUFx2_ASAP7_75t_L g4342 ( 
.A(n_3548),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_SL g4343 ( 
.A(n_3533),
.B(n_430),
.Y(n_4343)
);

A2O1A1Ixp33_ASAP7_75t_L g4344 ( 
.A1(n_3870),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_4344)
);

NOR2xp33_ASAP7_75t_L g4345 ( 
.A(n_4000),
.B(n_432),
.Y(n_4345)
);

AOI22xp5_ASAP7_75t_L g4346 ( 
.A1(n_3753),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_4346)
);

NAND2xp5_ASAP7_75t_SL g4347 ( 
.A(n_3533),
.B(n_435),
.Y(n_4347)
);

NAND2x1p5_ASAP7_75t_L g4348 ( 
.A(n_3639),
.B(n_435),
.Y(n_4348)
);

BUFx3_ASAP7_75t_L g4349 ( 
.A(n_3816),
.Y(n_4349)
);

OAI22x1_ASAP7_75t_L g4350 ( 
.A1(n_3704),
.A2(n_438),
.B1(n_435),
.B2(n_437),
.Y(n_4350)
);

OAI22xp5_ASAP7_75t_L g4351 ( 
.A1(n_3782),
.A2(n_440),
.B1(n_437),
.B2(n_439),
.Y(n_4351)
);

O2A1O1Ixp33_ASAP7_75t_L g4352 ( 
.A1(n_3995),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_4352)
);

AOI21xp5_ASAP7_75t_L g4353 ( 
.A1(n_3803),
.A2(n_439),
.B(n_441),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_SL g4354 ( 
.A(n_3533),
.B(n_441),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3873),
.Y(n_4355)
);

NOR2xp33_ASAP7_75t_R g4356 ( 
.A(n_3548),
.B(n_442),
.Y(n_4356)
);

AO32x1_ASAP7_75t_L g4357 ( 
.A1(n_3554),
.A2(n_444),
.A3(n_442),
.B1(n_443),
.B2(n_445),
.Y(n_4357)
);

BUFx2_ASAP7_75t_L g4358 ( 
.A(n_3548),
.Y(n_4358)
);

HB1xp67_ASAP7_75t_L g4359 ( 
.A(n_3749),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_3877),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_4029),
.B(n_4042),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_3526),
.B(n_3528),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_3530),
.B(n_443),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_3734),
.A2(n_444),
.B(n_445),
.Y(n_4364)
);

AO21x1_ASAP7_75t_L g4365 ( 
.A1(n_3647),
.A2(n_444),
.B(n_445),
.Y(n_4365)
);

AOI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_3764),
.A2(n_446),
.B(n_447),
.Y(n_4366)
);

NAND2x1p5_ASAP7_75t_L g4367 ( 
.A(n_3749),
.B(n_446),
.Y(n_4367)
);

AOI21xp5_ASAP7_75t_L g4368 ( 
.A1(n_3764),
.A2(n_447),
.B(n_448),
.Y(n_4368)
);

INVx3_ASAP7_75t_L g4369 ( 
.A(n_3816),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_SL g4370 ( 
.A(n_3534),
.B(n_448),
.Y(n_4370)
);

AOI21xp5_ASAP7_75t_L g4371 ( 
.A1(n_3882),
.A2(n_448),
.B(n_449),
.Y(n_4371)
);

AOI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_3760),
.A2(n_3785),
.B1(n_3915),
.B2(n_3828),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_SL g4373 ( 
.A(n_3534),
.B(n_449),
.Y(n_4373)
);

A2O1A1Ixp33_ASAP7_75t_L g4374 ( 
.A1(n_3541),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_4374)
);

HB1xp67_ASAP7_75t_L g4375 ( 
.A(n_3808),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_3539),
.B(n_450),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_3498),
.Y(n_4377)
);

BUFx6f_ASAP7_75t_L g4378 ( 
.A(n_3534),
.Y(n_4378)
);

NOR2xp33_ASAP7_75t_L g4379 ( 
.A(n_4009),
.B(n_450),
.Y(n_4379)
);

NOR2xp33_ASAP7_75t_L g4380 ( 
.A(n_4011),
.B(n_451),
.Y(n_4380)
);

INVx8_ASAP7_75t_L g4381 ( 
.A(n_3548),
.Y(n_4381)
);

AOI21xp5_ASAP7_75t_L g4382 ( 
.A1(n_3882),
.A2(n_451),
.B(n_452),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_3902),
.B(n_452),
.Y(n_4383)
);

AND2x2_ASAP7_75t_L g4384 ( 
.A(n_3931),
.B(n_453),
.Y(n_4384)
);

BUFx12f_ASAP7_75t_L g4385 ( 
.A(n_3600),
.Y(n_4385)
);

INVx1_ASAP7_75t_SL g4386 ( 
.A(n_3808),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_3879),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_3542),
.Y(n_4388)
);

NOR2xp33_ASAP7_75t_L g4389 ( 
.A(n_3887),
.B(n_453),
.Y(n_4389)
);

AOI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_4040),
.A2(n_453),
.B(n_454),
.Y(n_4390)
);

OAI22x1_ASAP7_75t_L g4391 ( 
.A1(n_4006),
.A2(n_456),
.B1(n_454),
.B2(n_455),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_SL g4392 ( 
.A(n_3705),
.B(n_455),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4024),
.B(n_455),
.Y(n_4393)
);

OAI221xp5_ASAP7_75t_L g4394 ( 
.A1(n_3903),
.A2(n_3908),
.B1(n_3994),
.B2(n_3798),
.C(n_3788),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_SL g4395 ( 
.A(n_3705),
.B(n_457),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_3689),
.B(n_457),
.Y(n_4396)
);

AOI21xp5_ASAP7_75t_L g4397 ( 
.A1(n_3705),
.A2(n_457),
.B(n_458),
.Y(n_4397)
);

O2A1O1Ixp33_ASAP7_75t_L g4398 ( 
.A1(n_4005),
.A2(n_460),
.B(n_458),
.C(n_459),
.Y(n_4398)
);

CKINVDCx5p33_ASAP7_75t_R g4399 ( 
.A(n_3600),
.Y(n_4399)
);

CKINVDCx5p33_ASAP7_75t_R g4400 ( 
.A(n_3600),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_3751),
.B(n_459),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_3566),
.B(n_459),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_3577),
.B(n_460),
.Y(n_4403)
);

AOI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_3836),
.A2(n_460),
.B(n_461),
.Y(n_4404)
);

BUFx3_ASAP7_75t_L g4405 ( 
.A(n_4046),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_3579),
.B(n_461),
.Y(n_4406)
);

AOI21xp5_ASAP7_75t_L g4407 ( 
.A1(n_3836),
.A2(n_461),
.B(n_462),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_3498),
.Y(n_4408)
);

INVx1_ASAP7_75t_SL g4409 ( 
.A(n_3836),
.Y(n_4409)
);

INVx3_ASAP7_75t_L g4410 ( 
.A(n_4046),
.Y(n_4410)
);

BUFx6f_ASAP7_75t_L g4411 ( 
.A(n_3893),
.Y(n_4411)
);

AOI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_3893),
.A2(n_462),
.B(n_463),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_3945),
.B(n_462),
.Y(n_4413)
);

OAI22xp5_ASAP7_75t_L g4414 ( 
.A1(n_3757),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_4414)
);

AOI21xp5_ASAP7_75t_L g4415 ( 
.A1(n_3893),
.A2(n_463),
.B(n_464),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_3582),
.B(n_464),
.Y(n_4416)
);

AOI21xp5_ASAP7_75t_L g4417 ( 
.A1(n_3883),
.A2(n_3708),
.B(n_3682),
.Y(n_4417)
);

AOI22xp33_ASAP7_75t_L g4418 ( 
.A1(n_3800),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_4418)
);

AND2x2_ASAP7_75t_L g4419 ( 
.A(n_3970),
.B(n_466),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_SL g4420 ( 
.A(n_3884),
.B(n_468),
.Y(n_4420)
);

AOI21x1_ASAP7_75t_L g4421 ( 
.A1(n_3524),
.A2(n_3532),
.B(n_3756),
.Y(n_4421)
);

A2O1A1Ixp33_ASAP7_75t_L g4422 ( 
.A1(n_3544),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_3586),
.B(n_3587),
.Y(n_4423)
);

OR2x2_ASAP7_75t_L g4424 ( 
.A(n_3929),
.B(n_468),
.Y(n_4424)
);

NOR2xp33_ASAP7_75t_SL g4425 ( 
.A(n_3600),
.B(n_469),
.Y(n_4425)
);

NOR2xp33_ASAP7_75t_L g4426 ( 
.A(n_3937),
.B(n_3941),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_3939),
.Y(n_4427)
);

INVx3_ASAP7_75t_L g4428 ( 
.A(n_3950),
.Y(n_4428)
);

BUFx3_ASAP7_75t_L g4429 ( 
.A(n_3954),
.Y(n_4429)
);

AOI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_3715),
.A2(n_469),
.B(n_470),
.Y(n_4430)
);

A2O1A1Ixp33_ASAP7_75t_SL g4431 ( 
.A1(n_4025),
.A2(n_472),
.B(n_470),
.C(n_471),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_3588),
.Y(n_4432)
);

NOR2xp33_ASAP7_75t_L g4433 ( 
.A(n_3957),
.B(n_471),
.Y(n_4433)
);

AOI21xp5_ASAP7_75t_L g4434 ( 
.A1(n_3597),
.A2(n_3946),
.B(n_3558),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_3894),
.Y(n_4435)
);

INVx3_ASAP7_75t_L g4436 ( 
.A(n_4050),
.Y(n_4436)
);

BUFx2_ASAP7_75t_L g4437 ( 
.A(n_3997),
.Y(n_4437)
);

AOI33xp33_ASAP7_75t_L g4438 ( 
.A1(n_3657),
.A2(n_473),
.A3(n_475),
.B1(n_471),
.B2(n_472),
.B3(n_474),
.Y(n_4438)
);

AOI21xp5_ASAP7_75t_L g4439 ( 
.A1(n_3597),
.A2(n_472),
.B(n_473),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_3589),
.B(n_473),
.Y(n_4440)
);

AO21x2_ASAP7_75t_L g4441 ( 
.A1(n_3814),
.A2(n_474),
.B(n_475),
.Y(n_4441)
);

O2A1O1Ixp33_ASAP7_75t_L g4442 ( 
.A1(n_4056),
.A2(n_477),
.B(n_474),
.C(n_475),
.Y(n_4442)
);

NOR2xp67_ASAP7_75t_L g4443 ( 
.A(n_3980),
.B(n_477),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_3593),
.B(n_477),
.Y(n_4444)
);

O2A1O1Ixp33_ASAP7_75t_L g4445 ( 
.A1(n_3881),
.A2(n_480),
.B(n_478),
.C(n_479),
.Y(n_4445)
);

AOI22xp5_ASAP7_75t_L g4446 ( 
.A1(n_3743),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_4446)
);

NOR2xp33_ASAP7_75t_L g4447 ( 
.A(n_3938),
.B(n_478),
.Y(n_4447)
);

O2A1O1Ixp5_ASAP7_75t_L g4448 ( 
.A1(n_3673),
.A2(n_482),
.B(n_479),
.C(n_481),
.Y(n_4448)
);

OAI22xp5_ASAP7_75t_L g4449 ( 
.A1(n_3880),
.A2(n_484),
.B1(n_481),
.B2(n_483),
.Y(n_4449)
);

AOI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_3568),
.A2(n_481),
.B(n_483),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_SL g4451 ( 
.A(n_3895),
.B(n_3555),
.Y(n_4451)
);

INVx3_ASAP7_75t_L g4452 ( 
.A(n_4007),
.Y(n_4452)
);

AND3x1_ASAP7_75t_SL g4453 ( 
.A(n_3972),
.B(n_483),
.C(n_485),
.Y(n_4453)
);

NOR2xp33_ASAP7_75t_L g4454 ( 
.A(n_3968),
.B(n_485),
.Y(n_4454)
);

AND2x4_ASAP7_75t_L g4455 ( 
.A(n_3967),
.B(n_485),
.Y(n_4455)
);

A2O1A1Ixp33_ASAP7_75t_SL g4456 ( 
.A1(n_3729),
.A2(n_488),
.B(n_486),
.C(n_487),
.Y(n_4456)
);

AOI22xp33_ASAP7_75t_SL g4457 ( 
.A1(n_3650),
.A2(n_488),
.B1(n_486),
.B2(n_487),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_3596),
.B(n_487),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_3602),
.B(n_489),
.Y(n_4459)
);

AOI21xp5_ASAP7_75t_L g4460 ( 
.A1(n_3759),
.A2(n_489),
.B(n_490),
.Y(n_4460)
);

INVx2_ASAP7_75t_SL g4461 ( 
.A(n_3974),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_SL g4462 ( 
.A(n_3809),
.B(n_489),
.Y(n_4462)
);

AOI21xp5_ASAP7_75t_L g4463 ( 
.A1(n_3557),
.A2(n_490),
.B(n_491),
.Y(n_4463)
);

INVx3_ASAP7_75t_L g4464 ( 
.A(n_3831),
.Y(n_4464)
);

NOR2xp33_ASAP7_75t_R g4465 ( 
.A(n_3697),
.B(n_3844),
.Y(n_4465)
);

A2O1A1Ixp33_ASAP7_75t_L g4466 ( 
.A1(n_3565),
.A2(n_3585),
.B(n_3661),
.C(n_3516),
.Y(n_4466)
);

AND2x2_ASAP7_75t_L g4467 ( 
.A(n_4023),
.B(n_491),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_3606),
.Y(n_4468)
);

AOI21xp5_ASAP7_75t_L g4469 ( 
.A1(n_3848),
.A2(n_491),
.B(n_492),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_3607),
.B(n_492),
.Y(n_4470)
);

INVx1_ASAP7_75t_SL g4471 ( 
.A(n_4033),
.Y(n_4471)
);

O2A1O1Ixp33_ASAP7_75t_SL g4472 ( 
.A1(n_3991),
.A2(n_494),
.B(n_492),
.C(n_493),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_3610),
.Y(n_4473)
);

A2O1A1Ixp33_ASAP7_75t_L g4474 ( 
.A1(n_3615),
.A2(n_3818),
.B(n_3806),
.C(n_4014),
.Y(n_4474)
);

BUFx6f_ASAP7_75t_L g4475 ( 
.A(n_3739),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_3613),
.B(n_3629),
.Y(n_4476)
);

NOR2xp33_ASAP7_75t_L g4477 ( 
.A(n_4038),
.B(n_493),
.Y(n_4477)
);

AOI222xp33_ASAP7_75t_L g4478 ( 
.A1(n_3783),
.A2(n_517),
.B1(n_501),
.B2(n_525),
.C1(n_509),
.C2(n_493),
.Y(n_4478)
);

BUFx6f_ASAP7_75t_L g4479 ( 
.A(n_4045),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_3641),
.B(n_494),
.Y(n_4480)
);

INVx3_ASAP7_75t_L g4481 ( 
.A(n_3868),
.Y(n_4481)
);

OAI22xp5_ASAP7_75t_L g4482 ( 
.A1(n_3891),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_4482)
);

HB1xp67_ASAP7_75t_L g4483 ( 
.A(n_3642),
.Y(n_4483)
);

NOR2xp33_ASAP7_75t_L g4484 ( 
.A(n_3619),
.B(n_496),
.Y(n_4484)
);

OAI21xp33_ASAP7_75t_L g4485 ( 
.A1(n_3688),
.A2(n_497),
.B(n_498),
.Y(n_4485)
);

A2O1A1Ixp33_ASAP7_75t_L g4486 ( 
.A1(n_3553),
.A2(n_499),
.B(n_497),
.C(n_498),
.Y(n_4486)
);

INVx4_ASAP7_75t_L g4487 ( 
.A(n_4003),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_3648),
.Y(n_4488)
);

NOR2xp67_ASAP7_75t_L g4489 ( 
.A(n_4049),
.B(n_497),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_3654),
.Y(n_4490)
);

AOI21xp5_ASAP7_75t_L g4491 ( 
.A1(n_3850),
.A2(n_499),
.B(n_500),
.Y(n_4491)
);

AOI21xp5_ASAP7_75t_L g4492 ( 
.A1(n_3854),
.A2(n_3861),
.B(n_3856),
.Y(n_4492)
);

NAND3xp33_ASAP7_75t_SL g4493 ( 
.A(n_3494),
.B(n_499),
.C(n_500),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_3655),
.B(n_500),
.Y(n_4494)
);

CKINVDCx5p33_ASAP7_75t_R g4495 ( 
.A(n_3927),
.Y(n_4495)
);

BUFx12f_ASAP7_75t_L g4496 ( 
.A(n_3686),
.Y(n_4496)
);

INVxp67_ASAP7_75t_L g4497 ( 
.A(n_3976),
.Y(n_4497)
);

NOR2xp33_ASAP7_75t_L g4498 ( 
.A(n_3623),
.B(n_501),
.Y(n_4498)
);

CKINVDCx5p33_ASAP7_75t_R g4499 ( 
.A(n_3638),
.Y(n_4499)
);

OAI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_3525),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_4500)
);

A2O1A1Ixp33_ASAP7_75t_L g4501 ( 
.A1(n_3746),
.A2(n_504),
.B(n_502),
.C(n_503),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_SL g4502 ( 
.A(n_4051),
.B(n_502),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_L g4503 ( 
.A(n_3658),
.B(n_503),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_3664),
.B(n_505),
.Y(n_4504)
);

OAI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_3769),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_4505)
);

A2O1A1Ixp33_ASAP7_75t_L g4506 ( 
.A1(n_3964),
.A2(n_508),
.B(n_506),
.C(n_507),
.Y(n_4506)
);

AOI21xp5_ASAP7_75t_L g4507 ( 
.A1(n_3864),
.A2(n_506),
.B(n_508),
.Y(n_4507)
);

A2O1A1Ixp33_ASAP7_75t_L g4508 ( 
.A1(n_3965),
.A2(n_510),
.B(n_508),
.C(n_509),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_SL g4509 ( 
.A(n_3975),
.B(n_509),
.Y(n_4509)
);

OAI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_3849),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_4510)
);

INVx5_ASAP7_75t_L g4511 ( 
.A(n_3686),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_3667),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_3668),
.B(n_510),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_3683),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_3691),
.B(n_511),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_SL g4516 ( 
.A(n_3598),
.B(n_512),
.Y(n_4516)
);

CKINVDCx5p33_ASAP7_75t_R g4517 ( 
.A(n_3984),
.Y(n_4517)
);

OAI22xp5_ASAP7_75t_L g4518 ( 
.A1(n_3576),
.A2(n_515),
.B1(n_513),
.B2(n_514),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_3695),
.B(n_513),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_3701),
.B(n_3731),
.Y(n_4520)
);

INVxp67_ASAP7_75t_L g4521 ( 
.A(n_3911),
.Y(n_4521)
);

AOI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_3735),
.A2(n_514),
.B(n_515),
.Y(n_4522)
);

AOI221x1_ASAP7_75t_L g4523 ( 
.A1(n_3496),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.C(n_518),
.Y(n_4523)
);

CKINVDCx5p33_ASAP7_75t_R g4524 ( 
.A(n_3919),
.Y(n_4524)
);

OAI22xp5_ASAP7_75t_L g4525 ( 
.A1(n_3745),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_3748),
.B(n_518),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_3763),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_3775),
.Y(n_4528)
);

NOR2xp33_ASAP7_75t_L g4529 ( 
.A(n_3776),
.B(n_519),
.Y(n_4529)
);

NAND2x1p5_ASAP7_75t_L g4530 ( 
.A(n_4013),
.B(n_519),
.Y(n_4530)
);

OAI21xp33_ASAP7_75t_L g4531 ( 
.A1(n_3922),
.A2(n_520),
.B(n_521),
.Y(n_4531)
);

INVx2_ASAP7_75t_L g4532 ( 
.A(n_3778),
.Y(n_4532)
);

CKINVDCx6p67_ASAP7_75t_R g4533 ( 
.A(n_3790),
.Y(n_4533)
);

AOI21xp5_ASAP7_75t_L g4534 ( 
.A1(n_3791),
.A2(n_520),
.B(n_521),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_3797),
.Y(n_4535)
);

CKINVDCx5p33_ASAP7_75t_R g4536 ( 
.A(n_3799),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_3801),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_3807),
.B(n_520),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_3812),
.Y(n_4539)
);

NOR2xp67_ASAP7_75t_L g4540 ( 
.A(n_3817),
.B(n_522),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_3822),
.B(n_522),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_SL g4542 ( 
.A(n_3959),
.B(n_522),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_SL g4543 ( 
.A(n_3512),
.B(n_523),
.Y(n_4543)
);

AOI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_3823),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_4544)
);

O2A1O1Ixp33_ASAP7_75t_L g4545 ( 
.A1(n_3827),
.A2(n_528),
.B(n_524),
.C(n_527),
.Y(n_4545)
);

INVx1_ASAP7_75t_SL g4546 ( 
.A(n_4026),
.Y(n_4546)
);

AO32x2_ASAP7_75t_L g4547 ( 
.A1(n_4001),
.A2(n_528),
.A3(n_524),
.B1(n_527),
.B2(n_529),
.Y(n_4547)
);

O2A1O1Ixp33_ASAP7_75t_L g4548 ( 
.A1(n_3973),
.A2(n_531),
.B(n_529),
.C(n_530),
.Y(n_4548)
);

INVx2_ASAP7_75t_SL g4549 ( 
.A(n_4027),
.Y(n_4549)
);

AOI21xp5_ASAP7_75t_L g4550 ( 
.A1(n_3513),
.A2(n_529),
.B(n_530),
.Y(n_4550)
);

AOI21xp5_ASAP7_75t_L g4551 ( 
.A1(n_3962),
.A2(n_530),
.B(n_532),
.Y(n_4551)
);

BUFx3_ASAP7_75t_L g4552 ( 
.A(n_3920),
.Y(n_4552)
);

AOI21xp5_ASAP7_75t_L g4553 ( 
.A1(n_3963),
.A2(n_532),
.B(n_533),
.Y(n_4553)
);

AOI22xp33_ASAP7_75t_L g4554 ( 
.A1(n_3982),
.A2(n_534),
.B1(n_532),
.B2(n_533),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_SL g4555 ( 
.A(n_3810),
.B(n_534),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_3686),
.Y(n_4556)
);

AOI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_3958),
.A2(n_534),
.B(n_535),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_SL g4558 ( 
.A(n_3725),
.B(n_535),
.Y(n_4558)
);

OAI21xp5_ASAP7_75t_L g4559 ( 
.A1(n_3985),
.A2(n_535),
.B(n_536),
.Y(n_4559)
);

AOI21xp5_ASAP7_75t_L g4560 ( 
.A1(n_4001),
.A2(n_536),
.B(n_537),
.Y(n_4560)
);

OAI22xp5_ASAP7_75t_L g4561 ( 
.A1(n_4035),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_3767),
.B(n_537),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_L g4563 ( 
.A(n_3768),
.B(n_538),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_SL g4564 ( 
.A(n_3736),
.B(n_538),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_4001),
.A2(n_539),
.B(n_540),
.Y(n_4565)
);

A2O1A1Ixp33_ASAP7_75t_L g4566 ( 
.A1(n_3917),
.A2(n_541),
.B(n_539),
.C(n_540),
.Y(n_4566)
);

NAND2xp33_ASAP7_75t_SL g4567 ( 
.A(n_3773),
.B(n_539),
.Y(n_4567)
);

OAI22xp5_ASAP7_75t_L g4568 ( 
.A1(n_3779),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_4568)
);

AOI21xp5_ASAP7_75t_L g4569 ( 
.A1(n_3538),
.A2(n_541),
.B(n_542),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_3711),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_3781),
.B(n_3793),
.Y(n_4571)
);

CKINVDCx11_ASAP7_75t_R g4572 ( 
.A(n_3694),
.Y(n_4572)
);

A2O1A1Ixp33_ASAP7_75t_L g4573 ( 
.A1(n_3989),
.A2(n_544),
.B(n_542),
.C(n_543),
.Y(n_4573)
);

AOI21xp5_ASAP7_75t_L g4574 ( 
.A1(n_3540),
.A2(n_543),
.B(n_544),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_3914),
.Y(n_4575)
);

NOR2xp33_ASAP7_75t_L g4576 ( 
.A(n_4053),
.B(n_543),
.Y(n_4576)
);

BUFx6f_ASAP7_75t_L g4577 ( 
.A(n_3921),
.Y(n_4577)
);

CKINVDCx20_ASAP7_75t_R g4578 ( 
.A(n_4058),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_3815),
.B(n_3825),
.Y(n_4579)
);

INVx4_ASAP7_75t_L g4580 ( 
.A(n_3718),
.Y(n_4580)
);

INVx4_ASAP7_75t_L g4581 ( 
.A(n_3720),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_3830),
.B(n_544),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_3833),
.B(n_545),
.Y(n_4583)
);

AOI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_3723),
.A2(n_545),
.B(n_546),
.Y(n_4584)
);

CKINVDCx5p33_ASAP7_75t_R g4585 ( 
.A(n_3996),
.Y(n_4585)
);

INVx2_ASAP7_75t_L g4586 ( 
.A(n_3560),
.Y(n_4586)
);

A2O1A1Ixp33_ASAP7_75t_L g4587 ( 
.A1(n_3841),
.A2(n_547),
.B(n_545),
.C(n_546),
.Y(n_4587)
);

OR2x2_ASAP7_75t_L g4588 ( 
.A(n_3845),
.B(n_547),
.Y(n_4588)
);

NOR2xp33_ASAP7_75t_L g4589 ( 
.A(n_3846),
.B(n_547),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_3795),
.Y(n_4590)
);

OAI22xp5_ASAP7_75t_L g4591 ( 
.A1(n_3796),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_4591)
);

HB1xp67_ASAP7_75t_L g4592 ( 
.A(n_3678),
.Y(n_4592)
);

OAI22xp5_ASAP7_75t_L g4593 ( 
.A1(n_3805),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_4593)
);

A2O1A1Ixp33_ASAP7_75t_L g4594 ( 
.A1(n_3898),
.A2(n_551),
.B(n_549),
.C(n_550),
.Y(n_4594)
);

O2A1O1Ixp33_ASAP7_75t_L g4595 ( 
.A1(n_3765),
.A2(n_553),
.B(n_551),
.C(n_552),
.Y(n_4595)
);

BUFx2_ASAP7_75t_L g4596 ( 
.A(n_3679),
.Y(n_4596)
);

NOR2x1_ASAP7_75t_L g4597 ( 
.A(n_3901),
.B(n_552),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_SL g4598 ( 
.A(n_3567),
.B(n_552),
.Y(n_4598)
);

NOR2xp33_ASAP7_75t_L g4599 ( 
.A(n_3928),
.B(n_553),
.Y(n_4599)
);

NOR2xp33_ASAP7_75t_L g4600 ( 
.A(n_3940),
.B(n_554),
.Y(n_4600)
);

AOI21x1_ASAP7_75t_L g4601 ( 
.A1(n_3569),
.A2(n_849),
.B(n_846),
.Y(n_4601)
);

OAI22xp5_ASAP7_75t_L g4602 ( 
.A1(n_3570),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.Y(n_4602)
);

AOI21xp5_ASAP7_75t_L g4603 ( 
.A1(n_3571),
.A2(n_554),
.B(n_555),
.Y(n_4603)
);

O2A1O1Ixp33_ASAP7_75t_L g4604 ( 
.A1(n_3680),
.A2(n_558),
.B(n_556),
.C(n_557),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_3692),
.B(n_556),
.Y(n_4605)
);

INVxp67_ASAP7_75t_SL g4606 ( 
.A(n_3578),
.Y(n_4606)
);

O2A1O1Ixp33_ASAP7_75t_L g4607 ( 
.A1(n_3581),
.A2(n_559),
.B(n_557),
.C(n_558),
.Y(n_4607)
);

AOI21xp5_ASAP7_75t_L g4608 ( 
.A1(n_3583),
.A2(n_557),
.B(n_558),
.Y(n_4608)
);

OAI22xp5_ASAP7_75t_L g4609 ( 
.A1(n_3590),
.A2(n_561),
.B1(n_559),
.B2(n_560),
.Y(n_4609)
);

NAND3xp33_ASAP7_75t_SL g4610 ( 
.A(n_3942),
.B(n_559),
.C(n_560),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_3591),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_3592),
.B(n_560),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_3594),
.Y(n_4613)
);

O2A1O1Ixp5_ASAP7_75t_L g4614 ( 
.A1(n_3608),
.A2(n_563),
.B(n_561),
.C(n_562),
.Y(n_4614)
);

OR2x2_ASAP7_75t_L g4615 ( 
.A(n_3609),
.B(n_561),
.Y(n_4615)
);

AND2x4_ASAP7_75t_L g4616 ( 
.A(n_3612),
.B(n_562),
.Y(n_4616)
);

NOR2xp33_ASAP7_75t_R g4617 ( 
.A(n_3625),
.B(n_562),
.Y(n_4617)
);

AOI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_3627),
.A2(n_566),
.B1(n_564),
.B2(n_565),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_3640),
.B(n_564),
.Y(n_4619)
);

HB1xp67_ASAP7_75t_L g4620 ( 
.A(n_3643),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_3659),
.B(n_565),
.Y(n_4621)
);

INVx2_ASAP7_75t_L g4622 ( 
.A(n_3660),
.Y(n_4622)
);

AND2x4_ASAP7_75t_L g4623 ( 
.A(n_3662),
.B(n_565),
.Y(n_4623)
);

BUFx3_ASAP7_75t_L g4624 ( 
.A(n_4152),
.Y(n_4624)
);

BUFx2_ASAP7_75t_L g4625 ( 
.A(n_4194),
.Y(n_4625)
);

BUFx6f_ASAP7_75t_L g4626 ( 
.A(n_4254),
.Y(n_4626)
);

BUFx3_ASAP7_75t_L g4627 ( 
.A(n_4177),
.Y(n_4627)
);

NOR2xp33_ASAP7_75t_L g4628 ( 
.A(n_4533),
.B(n_566),
.Y(n_4628)
);

BUFx6f_ASAP7_75t_L g4629 ( 
.A(n_4257),
.Y(n_4629)
);

OR2x2_ASAP7_75t_L g4630 ( 
.A(n_4361),
.B(n_566),
.Y(n_4630)
);

INVx5_ASAP7_75t_SL g4631 ( 
.A(n_4207),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4067),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4085),
.Y(n_4633)
);

INVx3_ASAP7_75t_L g4634 ( 
.A(n_4201),
.Y(n_4634)
);

INVx2_ASAP7_75t_L g4635 ( 
.A(n_4270),
.Y(n_4635)
);

BUFx6f_ASAP7_75t_L g4636 ( 
.A(n_4147),
.Y(n_4636)
);

INVx1_ASAP7_75t_SL g4637 ( 
.A(n_4272),
.Y(n_4637)
);

BUFx2_ASAP7_75t_L g4638 ( 
.A(n_4320),
.Y(n_4638)
);

BUFx3_ASAP7_75t_L g4639 ( 
.A(n_4177),
.Y(n_4639)
);

BUFx2_ASAP7_75t_L g4640 ( 
.A(n_4320),
.Y(n_4640)
);

CKINVDCx5p33_ASAP7_75t_R g4641 ( 
.A(n_4121),
.Y(n_4641)
);

INVx3_ASAP7_75t_L g4642 ( 
.A(n_4201),
.Y(n_4642)
);

BUFx6f_ASAP7_75t_L g4643 ( 
.A(n_4228),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4062),
.B(n_3949),
.Y(n_4644)
);

BUFx2_ASAP7_75t_SL g4645 ( 
.A(n_4119),
.Y(n_4645)
);

INVx2_ASAP7_75t_SL g4646 ( 
.A(n_4159),
.Y(n_4646)
);

BUFx2_ASAP7_75t_L g4647 ( 
.A(n_4144),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4157),
.Y(n_4648)
);

BUFx2_ASAP7_75t_L g4649 ( 
.A(n_4144),
.Y(n_4649)
);

AND2x4_ASAP7_75t_L g4650 ( 
.A(n_4088),
.B(n_3956),
.Y(n_4650)
);

NOR2xp33_ASAP7_75t_L g4651 ( 
.A(n_4131),
.B(n_567),
.Y(n_4651)
);

BUFx2_ASAP7_75t_SL g4652 ( 
.A(n_4119),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4178),
.Y(n_4653)
);

BUFx2_ASAP7_75t_L g4654 ( 
.A(n_4385),
.Y(n_4654)
);

BUFx12f_ASAP7_75t_L g4655 ( 
.A(n_4159),
.Y(n_4655)
);

BUFx2_ASAP7_75t_SL g4656 ( 
.A(n_4119),
.Y(n_4656)
);

BUFx12f_ASAP7_75t_L g4657 ( 
.A(n_4190),
.Y(n_4657)
);

BUFx3_ASAP7_75t_L g4658 ( 
.A(n_4073),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4179),
.Y(n_4659)
);

NAND2x1p5_ASAP7_75t_L g4660 ( 
.A(n_4093),
.B(n_3953),
.Y(n_4660)
);

INVx3_ASAP7_75t_L g4661 ( 
.A(n_4190),
.Y(n_4661)
);

INVx1_ASAP7_75t_SL g4662 ( 
.A(n_4282),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4209),
.B(n_567),
.Y(n_4663)
);

INVx1_ASAP7_75t_SL g4664 ( 
.A(n_4125),
.Y(n_4664)
);

INVx2_ASAP7_75t_SL g4665 ( 
.A(n_4129),
.Y(n_4665)
);

CKINVDCx14_ASAP7_75t_R g4666 ( 
.A(n_4189),
.Y(n_4666)
);

NAND2x1p5_ASAP7_75t_L g4667 ( 
.A(n_4246),
.B(n_567),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4200),
.Y(n_4668)
);

INVx4_ASAP7_75t_L g4669 ( 
.A(n_4300),
.Y(n_4669)
);

BUFx3_ASAP7_75t_L g4670 ( 
.A(n_4065),
.Y(n_4670)
);

INVx3_ASAP7_75t_L g4671 ( 
.A(n_4202),
.Y(n_4671)
);

BUFx6f_ASAP7_75t_L g4672 ( 
.A(n_4349),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4059),
.Y(n_4673)
);

BUFx6f_ASAP7_75t_L g4674 ( 
.A(n_4166),
.Y(n_4674)
);

CKINVDCx5p33_ASAP7_75t_R g4675 ( 
.A(n_4208),
.Y(n_4675)
);

INVx6_ASAP7_75t_L g4676 ( 
.A(n_4300),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4075),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4089),
.Y(n_4678)
);

OAI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4328),
.A2(n_4312),
.B1(n_4308),
.B2(n_4087),
.Y(n_4679)
);

NAND2x1p5_ASAP7_75t_L g4680 ( 
.A(n_4060),
.B(n_568),
.Y(n_4680)
);

BUFx3_ASAP7_75t_L g4681 ( 
.A(n_4218),
.Y(n_4681)
);

BUFx3_ASAP7_75t_L g4682 ( 
.A(n_4128),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4101),
.Y(n_4683)
);

BUFx12f_ASAP7_75t_L g4684 ( 
.A(n_4167),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4108),
.Y(n_4685)
);

BUFx10_ASAP7_75t_L g4686 ( 
.A(n_4227),
.Y(n_4686)
);

CKINVDCx16_ASAP7_75t_R g4687 ( 
.A(n_4247),
.Y(n_4687)
);

CKINVDCx6p67_ASAP7_75t_R g4688 ( 
.A(n_4283),
.Y(n_4688)
);

BUFx6f_ASAP7_75t_L g4689 ( 
.A(n_4166),
.Y(n_4689)
);

INVxp67_ASAP7_75t_L g4690 ( 
.A(n_4066),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4116),
.Y(n_4691)
);

BUFx2_ASAP7_75t_SL g4692 ( 
.A(n_4240),
.Y(n_4692)
);

INVx2_ASAP7_75t_L g4693 ( 
.A(n_4289),
.Y(n_4693)
);

INVx5_ASAP7_75t_L g4694 ( 
.A(n_4381),
.Y(n_4694)
);

INVx5_ASAP7_75t_L g4695 ( 
.A(n_4381),
.Y(n_4695)
);

INVx2_ASAP7_75t_SL g4696 ( 
.A(n_4100),
.Y(n_4696)
);

BUFx3_ASAP7_75t_L g4697 ( 
.A(n_4297),
.Y(n_4697)
);

AOI22xp5_ASAP7_75t_L g4698 ( 
.A1(n_4084),
.A2(n_4070),
.B1(n_4102),
.B2(n_4221),
.Y(n_4698)
);

BUFx3_ASAP7_75t_L g4699 ( 
.A(n_4297),
.Y(n_4699)
);

CKINVDCx16_ASAP7_75t_R g4700 ( 
.A(n_4356),
.Y(n_4700)
);

NAND2x1p5_ASAP7_75t_L g4701 ( 
.A(n_4274),
.B(n_569),
.Y(n_4701)
);

INVx2_ASAP7_75t_SL g4702 ( 
.A(n_4155),
.Y(n_4702)
);

CKINVDCx11_ASAP7_75t_R g4703 ( 
.A(n_4338),
.Y(n_4703)
);

INVxp67_ASAP7_75t_SL g4704 ( 
.A(n_4169),
.Y(n_4704)
);

BUFx12f_ASAP7_75t_L g4705 ( 
.A(n_4180),
.Y(n_4705)
);

BUFx3_ASAP7_75t_L g4706 ( 
.A(n_4215),
.Y(n_4706)
);

INVx4_ASAP7_75t_L g4707 ( 
.A(n_4240),
.Y(n_4707)
);

AO22x2_ASAP7_75t_L g4708 ( 
.A1(n_4063),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_4708)
);

NOR2xp33_ASAP7_75t_L g4709 ( 
.A(n_4517),
.B(n_569),
.Y(n_4709)
);

INVx1_ASAP7_75t_SL g4710 ( 
.A(n_4079),
.Y(n_4710)
);

BUFx2_ASAP7_75t_L g4711 ( 
.A(n_4281),
.Y(n_4711)
);

BUFx3_ASAP7_75t_L g4712 ( 
.A(n_4095),
.Y(n_4712)
);

BUFx12f_ASAP7_75t_L g4713 ( 
.A(n_4198),
.Y(n_4713)
);

AOI22xp5_ASAP7_75t_L g4714 ( 
.A1(n_4094),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_4714)
);

INVx2_ASAP7_75t_SL g4715 ( 
.A(n_4348),
.Y(n_4715)
);

INVx5_ASAP7_75t_L g4716 ( 
.A(n_4281),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4138),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4229),
.B(n_571),
.Y(n_4718)
);

INVx5_ASAP7_75t_L g4719 ( 
.A(n_4308),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4142),
.Y(n_4720)
);

AOI22xp5_ASAP7_75t_L g4721 ( 
.A1(n_4578),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.Y(n_4721)
);

INVx4_ASAP7_75t_L g4722 ( 
.A(n_4399),
.Y(n_4722)
);

INVx2_ASAP7_75t_L g4723 ( 
.A(n_4296),
.Y(n_4723)
);

CKINVDCx5p33_ASAP7_75t_R g4724 ( 
.A(n_4145),
.Y(n_4724)
);

BUFx2_ASAP7_75t_SL g4725 ( 
.A(n_4136),
.Y(n_4725)
);

NAND2x1p5_ASAP7_75t_L g4726 ( 
.A(n_4134),
.B(n_572),
.Y(n_4726)
);

INVx1_ASAP7_75t_SL g4727 ( 
.A(n_4123),
.Y(n_4727)
);

INVx5_ASAP7_75t_SL g4728 ( 
.A(n_4312),
.Y(n_4728)
);

BUFx3_ASAP7_75t_L g4729 ( 
.A(n_4405),
.Y(n_4729)
);

BUFx12f_ASAP7_75t_L g4730 ( 
.A(n_4367),
.Y(n_4730)
);

AND2x2_ASAP7_75t_L g4731 ( 
.A(n_4151),
.B(n_573),
.Y(n_4731)
);

INVx2_ASAP7_75t_SL g4732 ( 
.A(n_4269),
.Y(n_4732)
);

INVx2_ASAP7_75t_L g4733 ( 
.A(n_4305),
.Y(n_4733)
);

BUFx6f_ASAP7_75t_L g4734 ( 
.A(n_4166),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_SL g4735 ( 
.A(n_4425),
.B(n_573),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4164),
.B(n_574),
.Y(n_4736)
);

INVx2_ASAP7_75t_SL g4737 ( 
.A(n_4269),
.Y(n_4737)
);

BUFx6f_ASAP7_75t_L g4738 ( 
.A(n_4182),
.Y(n_4738)
);

AOI22xp33_ASAP7_75t_L g4739 ( 
.A1(n_4205),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4313),
.Y(n_4740)
);

CKINVDCx20_ASAP7_75t_R g4741 ( 
.A(n_4400),
.Y(n_4741)
);

BUFx2_ASAP7_75t_SL g4742 ( 
.A(n_4290),
.Y(n_4742)
);

BUFx6f_ASAP7_75t_L g4743 ( 
.A(n_4182),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4206),
.B(n_575),
.Y(n_4744)
);

INVx3_ASAP7_75t_L g4745 ( 
.A(n_4386),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4197),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4214),
.Y(n_4747)
);

CKINVDCx20_ASAP7_75t_R g4748 ( 
.A(n_4137),
.Y(n_4748)
);

INVx2_ASAP7_75t_L g4749 ( 
.A(n_4216),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_SL g4750 ( 
.A(n_4069),
.B(n_575),
.Y(n_4750)
);

CKINVDCx11_ASAP7_75t_R g4751 ( 
.A(n_4572),
.Y(n_4751)
);

BUFx3_ASAP7_75t_L g4752 ( 
.A(n_4369),
.Y(n_4752)
);

BUFx6f_ASAP7_75t_L g4753 ( 
.A(n_4182),
.Y(n_4753)
);

INVx3_ASAP7_75t_L g4754 ( 
.A(n_4239),
.Y(n_4754)
);

CKINVDCx20_ASAP7_75t_R g4755 ( 
.A(n_4536),
.Y(n_4755)
);

BUFx3_ASAP7_75t_L g4756 ( 
.A(n_4080),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4388),
.B(n_576),
.Y(n_4757)
);

BUFx3_ASAP7_75t_L g4758 ( 
.A(n_4091),
.Y(n_4758)
);

INVx1_ASAP7_75t_SL g4759 ( 
.A(n_4105),
.Y(n_4759)
);

AND2x4_ASAP7_75t_L g4760 ( 
.A(n_4311),
.B(n_577),
.Y(n_4760)
);

BUFx3_ASAP7_75t_L g4761 ( 
.A(n_4111),
.Y(n_4761)
);

AOI22xp33_ASAP7_75t_SL g4762 ( 
.A1(n_4072),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_SL g4763 ( 
.A(n_4342),
.B(n_577),
.Y(n_4763)
);

INVx2_ASAP7_75t_L g4764 ( 
.A(n_4264),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4127),
.Y(n_4765)
);

OAI22xp5_ASAP7_75t_L g4766 ( 
.A1(n_4090),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_4766)
);

NAND2x1p5_ASAP7_75t_L g4767 ( 
.A(n_4358),
.B(n_578),
.Y(n_4767)
);

NAND2x1p5_ASAP7_75t_L g4768 ( 
.A(n_4184),
.B(n_579),
.Y(n_4768)
);

INVx3_ASAP7_75t_L g4769 ( 
.A(n_4429),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4130),
.Y(n_4770)
);

BUFx2_ASAP7_75t_SL g4771 ( 
.A(n_4252),
.Y(n_4771)
);

NAND2x1p5_ASAP7_75t_L g4772 ( 
.A(n_4074),
.B(n_580),
.Y(n_4772)
);

INVx1_ASAP7_75t_SL g4773 ( 
.A(n_4112),
.Y(n_4773)
);

BUFx12f_ASAP7_75t_L g4774 ( 
.A(n_4495),
.Y(n_4774)
);

INVx2_ASAP7_75t_SL g4775 ( 
.A(n_4275),
.Y(n_4775)
);

INVx8_ASAP7_75t_L g4776 ( 
.A(n_4118),
.Y(n_4776)
);

BUFx4f_ASAP7_75t_SL g4777 ( 
.A(n_4109),
.Y(n_4777)
);

INVx5_ASAP7_75t_L g4778 ( 
.A(n_4251),
.Y(n_4778)
);

BUFx2_ASAP7_75t_L g4779 ( 
.A(n_4359),
.Y(n_4779)
);

INVx1_ASAP7_75t_SL g4780 ( 
.A(n_4409),
.Y(n_4780)
);

INVx5_ASAP7_75t_SL g4781 ( 
.A(n_4479),
.Y(n_4781)
);

INVx8_ASAP7_75t_L g4782 ( 
.A(n_4118),
.Y(n_4782)
);

BUFx2_ASAP7_75t_SL g4783 ( 
.A(n_4375),
.Y(n_4783)
);

AND2x4_ASAP7_75t_L g4784 ( 
.A(n_4064),
.B(n_581),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4467),
.B(n_4276),
.Y(n_4785)
);

BUFx3_ASAP7_75t_L g4786 ( 
.A(n_4092),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4284),
.B(n_580),
.Y(n_4787)
);

INVxp67_ASAP7_75t_SL g4788 ( 
.A(n_4291),
.Y(n_4788)
);

BUFx4_ASAP7_75t_SL g4789 ( 
.A(n_4524),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4427),
.Y(n_4790)
);

BUFx3_ASAP7_75t_L g4791 ( 
.A(n_4146),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4150),
.Y(n_4792)
);

AOI22xp33_ASAP7_75t_L g4793 ( 
.A1(n_4493),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_4793)
);

CKINVDCx5p33_ASAP7_75t_R g4794 ( 
.A(n_4188),
.Y(n_4794)
);

CKINVDCx5p33_ASAP7_75t_R g4795 ( 
.A(n_4076),
.Y(n_4795)
);

CKINVDCx5p33_ASAP7_75t_R g4796 ( 
.A(n_4499),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4158),
.Y(n_4797)
);

BUFx5_ASAP7_75t_L g4798 ( 
.A(n_4611),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4175),
.Y(n_4799)
);

INVx8_ASAP7_75t_L g4800 ( 
.A(n_4160),
.Y(n_4800)
);

BUFx4f_ASAP7_75t_L g4801 ( 
.A(n_4223),
.Y(n_4801)
);

BUFx3_ASAP7_75t_L g4802 ( 
.A(n_4251),
.Y(n_4802)
);

OR2x2_ASAP7_75t_L g4803 ( 
.A(n_4471),
.B(n_4086),
.Y(n_4803)
);

BUFx3_ASAP7_75t_L g4804 ( 
.A(n_4251),
.Y(n_4804)
);

INVx1_ASAP7_75t_SL g4805 ( 
.A(n_4292),
.Y(n_4805)
);

BUFx3_ASAP7_75t_L g4806 ( 
.A(n_4293),
.Y(n_4806)
);

BUFx6f_ASAP7_75t_L g4807 ( 
.A(n_4293),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4181),
.Y(n_4808)
);

NAND2x1p5_ASAP7_75t_L g4809 ( 
.A(n_4160),
.B(n_581),
.Y(n_4809)
);

INVx1_ASAP7_75t_SL g4810 ( 
.A(n_4293),
.Y(n_4810)
);

INVx1_ASAP7_75t_SL g4811 ( 
.A(n_4378),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_4488),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_L g4813 ( 
.A(n_4302),
.B(n_582),
.Y(n_4813)
);

BUFx6f_ASAP7_75t_L g4814 ( 
.A(n_4378),
.Y(n_4814)
);

INVx1_ASAP7_75t_SL g4815 ( 
.A(n_4378),
.Y(n_4815)
);

BUFx12f_ASAP7_75t_L g4816 ( 
.A(n_4479),
.Y(n_4816)
);

HB1xp67_ASAP7_75t_L g4817 ( 
.A(n_4479),
.Y(n_4817)
);

INVx3_ASAP7_75t_SL g4818 ( 
.A(n_4141),
.Y(n_4818)
);

BUFx6f_ASAP7_75t_L g4819 ( 
.A(n_4411),
.Y(n_4819)
);

NAND2x1p5_ASAP7_75t_L g4820 ( 
.A(n_4410),
.B(n_583),
.Y(n_4820)
);

BUFx3_ASAP7_75t_L g4821 ( 
.A(n_4411),
.Y(n_4821)
);

NOR2xp33_ASAP7_75t_L g4822 ( 
.A(n_4106),
.B(n_4124),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4183),
.Y(n_4823)
);

INVx2_ASAP7_75t_SL g4824 ( 
.A(n_4280),
.Y(n_4824)
);

BUFx2_ASAP7_75t_L g4825 ( 
.A(n_4303),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4185),
.Y(n_4826)
);

INVx1_ASAP7_75t_SL g4827 ( 
.A(n_4411),
.Y(n_4827)
);

BUFx12f_ASAP7_75t_L g4828 ( 
.A(n_4461),
.Y(n_4828)
);

BUFx6f_ASAP7_75t_L g4829 ( 
.A(n_4061),
.Y(n_4829)
);

BUFx6f_ASAP7_75t_L g4830 ( 
.A(n_4437),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_4490),
.Y(n_4831)
);

BUFx6f_ASAP7_75t_L g4832 ( 
.A(n_4428),
.Y(n_4832)
);

BUFx2_ASAP7_75t_R g4833 ( 
.A(n_4068),
.Y(n_4833)
);

INVxp67_ASAP7_75t_SL g4834 ( 
.A(n_4464),
.Y(n_4834)
);

BUFx4f_ASAP7_75t_SL g4835 ( 
.A(n_4496),
.Y(n_4835)
);

BUFx12f_ASAP7_75t_L g4836 ( 
.A(n_4585),
.Y(n_4836)
);

INVx4_ASAP7_75t_L g4837 ( 
.A(n_4455),
.Y(n_4837)
);

NAND2x1p5_ASAP7_75t_L g4838 ( 
.A(n_4326),
.B(n_583),
.Y(n_4838)
);

INVx1_ASAP7_75t_SL g4839 ( 
.A(n_4384),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4192),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4556),
.B(n_584),
.Y(n_4841)
);

INVx1_ASAP7_75t_SL g4842 ( 
.A(n_4413),
.Y(n_4842)
);

BUFx4f_ASAP7_75t_SL g4843 ( 
.A(n_4419),
.Y(n_4843)
);

INVx4_ASAP7_75t_L g4844 ( 
.A(n_4455),
.Y(n_4844)
);

INVx4_ASAP7_75t_L g4845 ( 
.A(n_4616),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4235),
.Y(n_4846)
);

BUFx2_ASAP7_75t_SL g4847 ( 
.A(n_4540),
.Y(n_4847)
);

INVx2_ASAP7_75t_L g4848 ( 
.A(n_4514),
.Y(n_4848)
);

INVx2_ASAP7_75t_L g4849 ( 
.A(n_4527),
.Y(n_4849)
);

CKINVDCx20_ASAP7_75t_R g4850 ( 
.A(n_4453),
.Y(n_4850)
);

CKINVDCx5p33_ASAP7_75t_R g4851 ( 
.A(n_4230),
.Y(n_4851)
);

NAND2x1p5_ASAP7_75t_L g4852 ( 
.A(n_4329),
.B(n_584),
.Y(n_4852)
);

BUFx3_ASAP7_75t_L g4853 ( 
.A(n_4199),
.Y(n_4853)
);

OR2x6_ASAP7_75t_L g4854 ( 
.A(n_4288),
.B(n_584),
.Y(n_4854)
);

INVx8_ASAP7_75t_L g4855 ( 
.A(n_4616),
.Y(n_4855)
);

AOI22xp33_ASAP7_75t_L g4856 ( 
.A1(n_4133),
.A2(n_4273),
.B1(n_4097),
.B2(n_4325),
.Y(n_4856)
);

AOI22xp33_ASAP7_75t_L g4857 ( 
.A1(n_4149),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4248),
.Y(n_4858)
);

BUFx12f_ASAP7_75t_L g4859 ( 
.A(n_4530),
.Y(n_4859)
);

BUFx2_ASAP7_75t_SL g4860 ( 
.A(n_4443),
.Y(n_4860)
);

INVx1_ASAP7_75t_SL g4861 ( 
.A(n_4424),
.Y(n_4861)
);

INVx1_ASAP7_75t_SL g4862 ( 
.A(n_4617),
.Y(n_4862)
);

BUFx2_ASAP7_75t_L g4863 ( 
.A(n_4483),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4528),
.Y(n_4864)
);

NAND2x1p5_ASAP7_75t_L g4865 ( 
.A(n_4331),
.B(n_585),
.Y(n_4865)
);

INVx4_ASAP7_75t_L g4866 ( 
.A(n_4623),
.Y(n_4866)
);

BUFx3_ASAP7_75t_L g4867 ( 
.A(n_4232),
.Y(n_4867)
);

BUFx12f_ASAP7_75t_L g4868 ( 
.A(n_4623),
.Y(n_4868)
);

INVx6_ASAP7_75t_SL g4869 ( 
.A(n_4077),
.Y(n_4869)
);

CKINVDCx16_ASAP7_75t_R g4870 ( 
.A(n_4161),
.Y(n_4870)
);

CKINVDCx5p33_ASAP7_75t_R g4871 ( 
.A(n_4287),
.Y(n_4871)
);

BUFx8_ASAP7_75t_L g4872 ( 
.A(n_4135),
.Y(n_4872)
);

BUFx2_ASAP7_75t_L g4873 ( 
.A(n_4465),
.Y(n_4873)
);

INVx4_ASAP7_75t_L g4874 ( 
.A(n_4436),
.Y(n_4874)
);

BUFx6f_ASAP7_75t_L g4875 ( 
.A(n_4577),
.Y(n_4875)
);

INVx2_ASAP7_75t_SL g4876 ( 
.A(n_4526),
.Y(n_4876)
);

INVx2_ASAP7_75t_L g4877 ( 
.A(n_4532),
.Y(n_4877)
);

INVx1_ASAP7_75t_SL g4878 ( 
.A(n_4396),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4539),
.Y(n_4879)
);

BUFx6f_ASAP7_75t_L g4880 ( 
.A(n_4577),
.Y(n_4880)
);

BUFx6f_ASAP7_75t_L g4881 ( 
.A(n_4577),
.Y(n_4881)
);

INVx3_ASAP7_75t_SL g4882 ( 
.A(n_4343),
.Y(n_4882)
);

INVx3_ASAP7_75t_L g4883 ( 
.A(n_4615),
.Y(n_4883)
);

BUFx12f_ASAP7_75t_L g4884 ( 
.A(n_4549),
.Y(n_4884)
);

CKINVDCx20_ASAP7_75t_R g4885 ( 
.A(n_4165),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4271),
.Y(n_4886)
);

INVx1_ASAP7_75t_SL g4887 ( 
.A(n_4113),
.Y(n_4887)
);

INVx8_ASAP7_75t_L g4888 ( 
.A(n_4605),
.Y(n_4888)
);

INVx2_ASAP7_75t_SL g4889 ( 
.A(n_4347),
.Y(n_4889)
);

INVx1_ASAP7_75t_SL g4890 ( 
.A(n_4139),
.Y(n_4890)
);

INVx1_ASAP7_75t_SL g4891 ( 
.A(n_4096),
.Y(n_4891)
);

INVx2_ASAP7_75t_SL g4892 ( 
.A(n_4354),
.Y(n_4892)
);

BUFx12f_ASAP7_75t_L g4893 ( 
.A(n_4588),
.Y(n_4893)
);

BUFx3_ASAP7_75t_L g4894 ( 
.A(n_4260),
.Y(n_4894)
);

AO22x2_ASAP7_75t_L g4895 ( 
.A1(n_4082),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_4895)
);

INVx2_ASAP7_75t_SL g4896 ( 
.A(n_4370),
.Y(n_4896)
);

BUFx2_ASAP7_75t_SL g4897 ( 
.A(n_4489),
.Y(n_4897)
);

NAND2xp5_ASAP7_75t_L g4898 ( 
.A(n_4324),
.B(n_587),
.Y(n_4898)
);

BUFx5_ASAP7_75t_L g4899 ( 
.A(n_4552),
.Y(n_4899)
);

INVxp67_ASAP7_75t_SL g4900 ( 
.A(n_4115),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4355),
.B(n_588),
.Y(n_4901)
);

INVx8_ASAP7_75t_L g4902 ( 
.A(n_4520),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4271),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_4360),
.B(n_588),
.Y(n_4904)
);

BUFx3_ASAP7_75t_L g4905 ( 
.A(n_4426),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_4387),
.B(n_588),
.Y(n_4906)
);

AOI22xp33_ASAP7_75t_L g4907 ( 
.A1(n_4394),
.A2(n_591),
.B1(n_589),
.B2(n_590),
.Y(n_4907)
);

INVx5_ASAP7_75t_L g4908 ( 
.A(n_4436),
.Y(n_4908)
);

BUFx6f_ASAP7_75t_L g4909 ( 
.A(n_4475),
.Y(n_4909)
);

OR2x6_ASAP7_75t_L g4910 ( 
.A(n_4132),
.B(n_4122),
.Y(n_4910)
);

INVx2_ASAP7_75t_SL g4911 ( 
.A(n_4373),
.Y(n_4911)
);

CKINVDCx16_ASAP7_75t_R g4912 ( 
.A(n_4143),
.Y(n_4912)
);

BUFx6f_ASAP7_75t_L g4913 ( 
.A(n_4475),
.Y(n_4913)
);

NAND2x1p5_ASAP7_75t_L g4914 ( 
.A(n_4392),
.B(n_589),
.Y(n_4914)
);

HB1xp67_ASAP7_75t_L g4915 ( 
.A(n_4596),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4511),
.B(n_589),
.Y(n_4916)
);

INVx1_ASAP7_75t_SL g4917 ( 
.A(n_4395),
.Y(n_4917)
);

INVx2_ASAP7_75t_L g4918 ( 
.A(n_4271),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4432),
.Y(n_4919)
);

INVx3_ASAP7_75t_L g4920 ( 
.A(n_4441),
.Y(n_4920)
);

CKINVDCx5p33_ASAP7_75t_R g4921 ( 
.A(n_4233),
.Y(n_4921)
);

BUFx6f_ASAP7_75t_L g4922 ( 
.A(n_4475),
.Y(n_4922)
);

BUFx2_ASAP7_75t_SL g4923 ( 
.A(n_4365),
.Y(n_4923)
);

BUFx2_ASAP7_75t_L g4924 ( 
.A(n_4307),
.Y(n_4924)
);

INVx3_ASAP7_75t_L g4925 ( 
.A(n_4487),
.Y(n_4925)
);

BUFx6f_ASAP7_75t_L g4926 ( 
.A(n_4187),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_4468),
.B(n_590),
.Y(n_4927)
);

BUFx3_ASAP7_75t_L g4928 ( 
.A(n_4477),
.Y(n_4928)
);

BUFx3_ASAP7_75t_L g4929 ( 
.A(n_4295),
.Y(n_4929)
);

BUFx3_ASAP7_75t_L g4930 ( 
.A(n_4306),
.Y(n_4930)
);

AOI22xp5_ASAP7_75t_L g4931 ( 
.A1(n_4372),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.Y(n_4931)
);

INVx2_ASAP7_75t_L g4932 ( 
.A(n_4153),
.Y(n_4932)
);

CKINVDCx8_ASAP7_75t_R g4933 ( 
.A(n_4511),
.Y(n_4933)
);

BUFx3_ASAP7_75t_L g4934 ( 
.A(n_4318),
.Y(n_4934)
);

BUFx3_ASAP7_75t_L g4935 ( 
.A(n_4473),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4512),
.Y(n_4936)
);

BUFx3_ASAP7_75t_L g4937 ( 
.A(n_4535),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4537),
.Y(n_4938)
);

NAND2x1p5_ASAP7_75t_L g4939 ( 
.A(n_4193),
.B(n_591),
.Y(n_4939)
);

CKINVDCx5p33_ASAP7_75t_R g4940 ( 
.A(n_4154),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_4377),
.Y(n_4941)
);

INVx1_ASAP7_75t_SL g4942 ( 
.A(n_4310),
.Y(n_4942)
);

NAND2x1p5_ASAP7_75t_L g4943 ( 
.A(n_4509),
.B(n_592),
.Y(n_4943)
);

INVx6_ASAP7_75t_L g4944 ( 
.A(n_4580),
.Y(n_4944)
);

BUFx2_ASAP7_75t_SL g4945 ( 
.A(n_4487),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4336),
.Y(n_4946)
);

BUFx2_ASAP7_75t_SL g4947 ( 
.A(n_4511),
.Y(n_4947)
);

INVx1_ASAP7_75t_SL g4948 ( 
.A(n_4319),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4391),
.Y(n_4949)
);

INVx3_ASAP7_75t_L g4950 ( 
.A(n_4580),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4521),
.B(n_592),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4226),
.Y(n_4952)
);

CKINVDCx20_ASAP7_75t_R g4953 ( 
.A(n_4497),
.Y(n_4953)
);

NAND2x1p5_ASAP7_75t_L g4954 ( 
.A(n_4597),
.B(n_593),
.Y(n_4954)
);

INVx8_ASAP7_75t_L g4955 ( 
.A(n_4277),
.Y(n_4955)
);

INVxp67_ASAP7_75t_SL g4956 ( 
.A(n_4452),
.Y(n_4956)
);

BUFx12f_ASAP7_75t_L g4957 ( 
.A(n_4581),
.Y(n_4957)
);

BUFx2_ASAP7_75t_L g4958 ( 
.A(n_4135),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4447),
.B(n_593),
.Y(n_4959)
);

CKINVDCx11_ASAP7_75t_R g4960 ( 
.A(n_4546),
.Y(n_4960)
);

INVx2_ASAP7_75t_L g4961 ( 
.A(n_4408),
.Y(n_4961)
);

INVx1_ASAP7_75t_SL g4962 ( 
.A(n_4321),
.Y(n_4962)
);

INVx1_ASAP7_75t_SL g4963 ( 
.A(n_4401),
.Y(n_4963)
);

BUFx3_ASAP7_75t_L g4964 ( 
.A(n_4345),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4350),
.Y(n_4965)
);

INVxp67_ASAP7_75t_SL g4966 ( 
.A(n_4481),
.Y(n_4966)
);

INVx2_ASAP7_75t_L g4967 ( 
.A(n_4547),
.Y(n_4967)
);

INVxp67_ASAP7_75t_SL g4968 ( 
.A(n_4592),
.Y(n_4968)
);

INVx4_ASAP7_75t_L g4969 ( 
.A(n_4581),
.Y(n_4969)
);

BUFx6f_ASAP7_75t_L g4970 ( 
.A(n_4612),
.Y(n_4970)
);

NAND2x1p5_ASAP7_75t_L g4971 ( 
.A(n_4446),
.B(n_594),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4435),
.Y(n_4972)
);

INVx2_ASAP7_75t_L g4973 ( 
.A(n_4547),
.Y(n_4973)
);

BUFx6f_ASAP7_75t_L g4974 ( 
.A(n_4619),
.Y(n_4974)
);

BUFx4f_ASAP7_75t_SL g4975 ( 
.A(n_4502),
.Y(n_4975)
);

BUFx2_ASAP7_75t_SL g4976 ( 
.A(n_4140),
.Y(n_4976)
);

INVxp67_ASAP7_75t_SL g4977 ( 
.A(n_4620),
.Y(n_4977)
);

BUFx2_ASAP7_75t_SL g4978 ( 
.A(n_4110),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4454),
.B(n_594),
.Y(n_4979)
);

INVx6_ASAP7_75t_L g4980 ( 
.A(n_4071),
.Y(n_4980)
);

BUFx3_ASAP7_75t_L g4981 ( 
.A(n_4379),
.Y(n_4981)
);

NAND2x1p5_ASAP7_75t_L g4982 ( 
.A(n_4210),
.B(n_594),
.Y(n_4982)
);

INVx2_ASAP7_75t_L g4983 ( 
.A(n_4547),
.Y(n_4983)
);

INVx2_ASAP7_75t_SL g4984 ( 
.A(n_4267),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4135),
.B(n_595),
.Y(n_4985)
);

BUFx2_ASAP7_75t_R g4986 ( 
.A(n_4393),
.Y(n_4986)
);

AND2x2_ASAP7_75t_L g4987 ( 
.A(n_4575),
.B(n_595),
.Y(n_4987)
);

INVx4_ASAP7_75t_L g4988 ( 
.A(n_4586),
.Y(n_4988)
);

INVx2_ASAP7_75t_SL g4989 ( 
.A(n_4330),
.Y(n_4989)
);

INVx3_ASAP7_75t_L g4990 ( 
.A(n_4601),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4438),
.Y(n_4991)
);

BUFx2_ASAP7_75t_L g4992 ( 
.A(n_4606),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_SL g4993 ( 
.A(n_4104),
.B(n_595),
.Y(n_4993)
);

HB1xp67_ASAP7_75t_L g4994 ( 
.A(n_4114),
.Y(n_4994)
);

INVx1_ASAP7_75t_SL g4995 ( 
.A(n_4263),
.Y(n_4995)
);

INVx2_ASAP7_75t_L g4996 ( 
.A(n_4421),
.Y(n_4996)
);

BUFx3_ASAP7_75t_L g4997 ( 
.A(n_4380),
.Y(n_4997)
);

INVx1_ASAP7_75t_SL g4998 ( 
.A(n_4078),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4316),
.Y(n_4999)
);

BUFx2_ASAP7_75t_SL g5000 ( 
.A(n_4332),
.Y(n_5000)
);

BUFx3_ASAP7_75t_L g5001 ( 
.A(n_4389),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4107),
.Y(n_5002)
);

INVx2_ASAP7_75t_L g5003 ( 
.A(n_4613),
.Y(n_5003)
);

BUFx6f_ASAP7_75t_L g5004 ( 
.A(n_4621),
.Y(n_5004)
);

BUFx6f_ASAP7_75t_L g5005 ( 
.A(n_4383),
.Y(n_5005)
);

AND2x4_ASAP7_75t_L g5006 ( 
.A(n_4117),
.B(n_597),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4590),
.B(n_596),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4107),
.Y(n_5008)
);

INVx3_ASAP7_75t_L g5009 ( 
.A(n_4562),
.Y(n_5009)
);

INVxp67_ASAP7_75t_SL g5010 ( 
.A(n_4244),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4402),
.Y(n_5011)
);

BUFx6f_ASAP7_75t_L g5012 ( 
.A(n_4563),
.Y(n_5012)
);

BUFx2_ASAP7_75t_L g5013 ( 
.A(n_4559),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4403),
.Y(n_5014)
);

INVx2_ASAP7_75t_SL g5015 ( 
.A(n_4213),
.Y(n_5015)
);

CKINVDCx6p67_ASAP7_75t_R g5016 ( 
.A(n_4225),
.Y(n_5016)
);

BUFx6f_ASAP7_75t_L g5017 ( 
.A(n_4582),
.Y(n_5017)
);

BUFx3_ASAP7_75t_L g5018 ( 
.A(n_4219),
.Y(n_5018)
);

BUFx6f_ASAP7_75t_SL g5019 ( 
.A(n_4478),
.Y(n_5019)
);

INVx2_ASAP7_75t_L g5020 ( 
.A(n_4622),
.Y(n_5020)
);

BUFx3_ASAP7_75t_L g5021 ( 
.A(n_4433),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4406),
.Y(n_5022)
);

INVx3_ASAP7_75t_SL g5023 ( 
.A(n_4516),
.Y(n_5023)
);

BUFx12f_ASAP7_75t_L g5024 ( 
.A(n_4457),
.Y(n_5024)
);

INVx2_ASAP7_75t_SL g5025 ( 
.A(n_4335),
.Y(n_5025)
);

INVx1_ASAP7_75t_SL g5026 ( 
.A(n_4341),
.Y(n_5026)
);

AND2x2_ASAP7_75t_L g5027 ( 
.A(n_4570),
.B(n_596),
.Y(n_5027)
);

INVx2_ASAP7_75t_L g5028 ( 
.A(n_4448),
.Y(n_5028)
);

NAND2x1p5_ASAP7_75t_L g5029 ( 
.A(n_4346),
.B(n_597),
.Y(n_5029)
);

INVx2_ASAP7_75t_L g5030 ( 
.A(n_4614),
.Y(n_5030)
);

CKINVDCx20_ASAP7_75t_R g5031 ( 
.A(n_4544),
.Y(n_5031)
);

INVx1_ASAP7_75t_SL g5032 ( 
.A(n_4363),
.Y(n_5032)
);

BUFx12f_ASAP7_75t_L g5033 ( 
.A(n_4126),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_L g5034 ( 
.A(n_4339),
.B(n_597),
.Y(n_5034)
);

BUFx12f_ASAP7_75t_L g5035 ( 
.A(n_4314),
.Y(n_5035)
);

INVx1_ASAP7_75t_SL g5036 ( 
.A(n_4376),
.Y(n_5036)
);

BUFx2_ASAP7_75t_SL g5037 ( 
.A(n_4351),
.Y(n_5037)
);

NAND2x1p5_ASAP7_75t_L g5038 ( 
.A(n_4618),
.B(n_598),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_4416),
.Y(n_5039)
);

AND2x2_ASAP7_75t_L g5040 ( 
.A(n_4560),
.B(n_598),
.Y(n_5040)
);

INVx2_ASAP7_75t_L g5041 ( 
.A(n_4362),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4423),
.B(n_599),
.Y(n_5042)
);

HB1xp67_ASAP7_75t_L g5043 ( 
.A(n_4440),
.Y(n_5043)
);

BUFx6f_ASAP7_75t_L g5044 ( 
.A(n_4583),
.Y(n_5044)
);

INVx2_ASAP7_75t_SL g5045 ( 
.A(n_4444),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_L g5046 ( 
.A(n_4476),
.B(n_599),
.Y(n_5046)
);

BUFx3_ASAP7_75t_L g5047 ( 
.A(n_4484),
.Y(n_5047)
);

BUFx4f_ASAP7_75t_SL g5048 ( 
.A(n_4462),
.Y(n_5048)
);

AND2x2_ASAP7_75t_L g5049 ( 
.A(n_4565),
.B(n_599),
.Y(n_5049)
);

BUFx3_ASAP7_75t_L g5050 ( 
.A(n_4498),
.Y(n_5050)
);

INVx8_ASAP7_75t_L g5051 ( 
.A(n_4234),
.Y(n_5051)
);

INVx1_ASAP7_75t_SL g5052 ( 
.A(n_4458),
.Y(n_5052)
);

AOI22xp33_ASAP7_75t_L g5053 ( 
.A1(n_4567),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_5053)
);

AOI22xp5_ASAP7_75t_L g5054 ( 
.A1(n_4098),
.A2(n_603),
.B1(n_600),
.B2(n_601),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4459),
.Y(n_5055)
);

INVx1_ASAP7_75t_SL g5056 ( 
.A(n_4470),
.Y(n_5056)
);

INVx5_ASAP7_75t_L g5057 ( 
.A(n_4357),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4480),
.Y(n_5058)
);

INVx2_ASAP7_75t_SL g5059 ( 
.A(n_4494),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_4529),
.B(n_600),
.Y(n_5060)
);

BUFx3_ASAP7_75t_L g5061 ( 
.A(n_4503),
.Y(n_5061)
);

BUFx12f_ASAP7_75t_L g5062 ( 
.A(n_4357),
.Y(n_5062)
);

BUFx3_ASAP7_75t_L g5063 ( 
.A(n_4504),
.Y(n_5063)
);

BUFx6f_ASAP7_75t_L g5064 ( 
.A(n_4513),
.Y(n_5064)
);

BUFx6f_ASAP7_75t_L g5065 ( 
.A(n_4515),
.Y(n_5065)
);

BUFx3_ASAP7_75t_L g5066 ( 
.A(n_4519),
.Y(n_5066)
);

BUFx6f_ASAP7_75t_L g5067 ( 
.A(n_4538),
.Y(n_5067)
);

NAND2x1p5_ASAP7_75t_L g5068 ( 
.A(n_4542),
.B(n_601),
.Y(n_5068)
);

INVx2_ASAP7_75t_L g5069 ( 
.A(n_4212),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_4541),
.B(n_603),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4420),
.Y(n_5071)
);

INVx2_ASAP7_75t_L g5072 ( 
.A(n_4333),
.Y(n_5072)
);

BUFx10_ASAP7_75t_L g5073 ( 
.A(n_4576),
.Y(n_5073)
);

BUFx2_ASAP7_75t_L g5074 ( 
.A(n_4211),
.Y(n_5074)
);

NOR2xp33_ASAP7_75t_L g5075 ( 
.A(n_4099),
.B(n_603),
.Y(n_5075)
);

BUFx6f_ASAP7_75t_L g5076 ( 
.A(n_4599),
.Y(n_5076)
);

BUFx6f_ASAP7_75t_L g5077 ( 
.A(n_4600),
.Y(n_5077)
);

BUFx6f_ASAP7_75t_SL g5078 ( 
.A(n_4250),
.Y(n_5078)
);

BUFx12f_ASAP7_75t_L g5079 ( 
.A(n_4397),
.Y(n_5079)
);

INVx3_ASAP7_75t_L g5080 ( 
.A(n_4571),
.Y(n_5080)
);

INVx2_ASAP7_75t_L g5081 ( 
.A(n_4168),
.Y(n_5081)
);

INVx1_ASAP7_75t_SL g5082 ( 
.A(n_4217),
.Y(n_5082)
);

CKINVDCx11_ASAP7_75t_R g5083 ( 
.A(n_4525),
.Y(n_5083)
);

INVx2_ASAP7_75t_L g5084 ( 
.A(n_4579),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_4294),
.Y(n_5085)
);

BUFx2_ASAP7_75t_L g5086 ( 
.A(n_4204),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4523),
.Y(n_5087)
);

INVx2_ASAP7_75t_L g5088 ( 
.A(n_4543),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4081),
.Y(n_5089)
);

BUFx2_ASAP7_75t_R g5090 ( 
.A(n_4451),
.Y(n_5090)
);

INVx3_ASAP7_75t_L g5091 ( 
.A(n_4327),
.Y(n_5091)
);

BUFx2_ASAP7_75t_L g5092 ( 
.A(n_4224),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4279),
.Y(n_5093)
);

OR2x6_ASAP7_75t_L g5094 ( 
.A(n_4222),
.B(n_604),
.Y(n_5094)
);

AND2x4_ASAP7_75t_L g5095 ( 
.A(n_4103),
.B(n_605),
.Y(n_5095)
);

BUFx12f_ASAP7_75t_L g5096 ( 
.A(n_4404),
.Y(n_5096)
);

INVx2_ASAP7_75t_L g5097 ( 
.A(n_4598),
.Y(n_5097)
);

NAND2x1p5_ASAP7_75t_L g5098 ( 
.A(n_4555),
.B(n_604),
.Y(n_5098)
);

AND2x4_ASAP7_75t_L g5099 ( 
.A(n_4625),
.B(n_4195),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_4668),
.B(n_4589),
.Y(n_5100)
);

INVx2_ASAP7_75t_SL g5101 ( 
.A(n_4902),
.Y(n_5101)
);

INVx2_ASAP7_75t_SL g5102 ( 
.A(n_4902),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_4632),
.Y(n_5103)
);

AND2x4_ASAP7_75t_L g5104 ( 
.A(n_4719),
.B(n_4083),
.Y(n_5104)
);

AO21x2_ASAP7_75t_L g5105 ( 
.A1(n_4996),
.A2(n_4148),
.B(n_4439),
.Y(n_5105)
);

OAI21x1_ASAP7_75t_L g5106 ( 
.A1(n_4990),
.A2(n_4434),
.B(n_4174),
.Y(n_5106)
);

OAI21x1_ASAP7_75t_L g5107 ( 
.A1(n_4925),
.A2(n_4492),
.B(n_4417),
.Y(n_5107)
);

NOR2xp33_ASAP7_75t_L g5108 ( 
.A(n_4669),
.B(n_605),
.Y(n_5108)
);

AOI21x1_ASAP7_75t_L g5109 ( 
.A1(n_4873),
.A2(n_4243),
.B(n_4242),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4633),
.Y(n_5110)
);

BUFx2_ASAP7_75t_L g5111 ( 
.A(n_4825),
.Y(n_5111)
);

OAI21x1_ASAP7_75t_L g5112 ( 
.A1(n_4920),
.A2(n_4203),
.B(n_4162),
.Y(n_5112)
);

OAI21x1_ASAP7_75t_L g5113 ( 
.A1(n_4950),
.A2(n_4170),
.B(n_4407),
.Y(n_5113)
);

OAI21x1_ASAP7_75t_L g5114 ( 
.A1(n_4918),
.A2(n_5020),
.B(n_5003),
.Y(n_5114)
);

OAI21x1_ASAP7_75t_L g5115 ( 
.A1(n_5080),
.A2(n_4415),
.B(n_4412),
.Y(n_5115)
);

OAI21x1_ASAP7_75t_SL g5116 ( 
.A1(n_4679),
.A2(n_4337),
.B(n_4317),
.Y(n_5116)
);

CKINVDCx20_ASAP7_75t_R g5117 ( 
.A(n_4666),
.Y(n_5117)
);

AND2x2_ASAP7_75t_L g5118 ( 
.A(n_4759),
.B(n_4773),
.Y(n_5118)
);

OA21x2_ASAP7_75t_L g5119 ( 
.A1(n_5002),
.A2(n_4531),
.B(n_4220),
.Y(n_5119)
);

A2O1A1Ixp33_ASAP7_75t_L g5120 ( 
.A1(n_4801),
.A2(n_4322),
.B(n_4340),
.C(n_4353),
.Y(n_5120)
);

OAI21xp5_ASAP7_75t_L g5121 ( 
.A1(n_4822),
.A2(n_4173),
.B(n_4171),
.Y(n_5121)
);

AOI221xp5_ASAP7_75t_L g5122 ( 
.A1(n_5019),
.A2(n_4955),
.B1(n_4946),
.B2(n_5078),
.C(n_4708),
.Y(n_5122)
);

OAI22xp5_ASAP7_75t_L g5123 ( 
.A1(n_4870),
.A2(n_4163),
.B1(n_4344),
.B2(n_4334),
.Y(n_5123)
);

AO21x2_ASAP7_75t_L g5124 ( 
.A1(n_5008),
.A2(n_4903),
.B(n_4886),
.Y(n_5124)
);

OAI21x1_ASAP7_75t_L g5125 ( 
.A1(n_4932),
.A2(n_4390),
.B(n_4450),
.Y(n_5125)
);

OAI21x1_ASAP7_75t_L g5126 ( 
.A1(n_5030),
.A2(n_4253),
.B(n_4245),
.Y(n_5126)
);

AND2x2_ASAP7_75t_L g5127 ( 
.A(n_4824),
.B(n_606),
.Y(n_5127)
);

INVx2_ASAP7_75t_L g5128 ( 
.A(n_4635),
.Y(n_5128)
);

AND2x2_ASAP7_75t_L g5129 ( 
.A(n_4839),
.B(n_606),
.Y(n_5129)
);

AND2x2_ASAP7_75t_L g5130 ( 
.A(n_4842),
.B(n_606),
.Y(n_5130)
);

AOI22xp33_ASAP7_75t_L g5131 ( 
.A1(n_4955),
.A2(n_4485),
.B1(n_4241),
.B2(n_4610),
.Y(n_5131)
);

AOI22xp5_ASAP7_75t_L g5132 ( 
.A1(n_4912),
.A2(n_4196),
.B1(n_4261),
.B2(n_4414),
.Y(n_5132)
);

INVx1_ASAP7_75t_SL g5133 ( 
.A(n_4624),
.Y(n_5133)
);

OAI21x1_ASAP7_75t_L g5134 ( 
.A1(n_4993),
.A2(n_4256),
.B(n_4278),
.Y(n_5134)
);

AND2x2_ASAP7_75t_L g5135 ( 
.A(n_4761),
.B(n_607),
.Y(n_5135)
);

AO21x2_ASAP7_75t_L g5136 ( 
.A1(n_4965),
.A2(n_4431),
.B(n_4456),
.Y(n_5136)
);

AO32x2_ASAP7_75t_L g5137 ( 
.A1(n_4969),
.A2(n_4323),
.A3(n_4249),
.B1(n_4482),
.B2(n_4449),
.Y(n_5137)
);

BUFx6f_ASAP7_75t_L g5138 ( 
.A(n_4626),
.Y(n_5138)
);

OA21x2_ASAP7_75t_L g5139 ( 
.A1(n_5089),
.A2(n_4924),
.B(n_4967),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_4648),
.Y(n_5140)
);

OAI21x1_ASAP7_75t_L g5141 ( 
.A1(n_5084),
.A2(n_4299),
.B(n_4298),
.Y(n_5141)
);

OAI21x1_ASAP7_75t_L g5142 ( 
.A1(n_4956),
.A2(n_4309),
.B(n_4301),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_4653),
.Y(n_5143)
);

OAI21xp5_ASAP7_75t_L g5144 ( 
.A1(n_5075),
.A2(n_4735),
.B(n_4714),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4659),
.Y(n_5145)
);

BUFx2_ASAP7_75t_L g5146 ( 
.A(n_4626),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_4919),
.Y(n_5147)
);

NAND2x1p5_ASAP7_75t_L g5148 ( 
.A(n_4627),
.B(n_4639),
.Y(n_5148)
);

INVx1_ASAP7_75t_L g5149 ( 
.A(n_4936),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4938),
.Y(n_5150)
);

OA21x2_ASAP7_75t_L g5151 ( 
.A1(n_4973),
.A2(n_4156),
.B(n_4374),
.Y(n_5151)
);

INVx2_ASAP7_75t_SL g5152 ( 
.A(n_4629),
.Y(n_5152)
);

OAI21x1_ASAP7_75t_L g5153 ( 
.A1(n_5069),
.A2(n_4366),
.B(n_4364),
.Y(n_5153)
);

OAI21xp5_ASAP7_75t_L g5154 ( 
.A1(n_4854),
.A2(n_4286),
.B(n_4268),
.Y(n_5154)
);

INVx3_ASAP7_75t_L g5155 ( 
.A(n_4629),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4863),
.Y(n_5156)
);

OAI21x1_ASAP7_75t_L g5157 ( 
.A1(n_5072),
.A2(n_4371),
.B(n_4368),
.Y(n_5157)
);

OAI21xp5_ASAP7_75t_L g5158 ( 
.A1(n_4854),
.A2(n_4534),
.B(n_4522),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_5041),
.B(n_4474),
.Y(n_5159)
);

OAI21x1_ASAP7_75t_L g5160 ( 
.A1(n_4834),
.A2(n_4382),
.B(n_4550),
.Y(n_5160)
);

OAI21xp5_ASAP7_75t_L g5161 ( 
.A1(n_4701),
.A2(n_4120),
.B(n_4422),
.Y(n_5161)
);

AO31x2_ASAP7_75t_L g5162 ( 
.A1(n_4874),
.A2(n_4172),
.A3(n_4505),
.B(n_4602),
.Y(n_5162)
);

INVx2_ASAP7_75t_L g5163 ( 
.A(n_4693),
.Y(n_5163)
);

AOI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_4855),
.A2(n_4472),
.B(n_4466),
.Y(n_5164)
);

OAI21x1_ASAP7_75t_L g5165 ( 
.A1(n_4966),
.A2(n_4603),
.B(n_4584),
.Y(n_5165)
);

BUFx6f_ASAP7_75t_L g5166 ( 
.A(n_4636),
.Y(n_5166)
);

AOI22xp33_ASAP7_75t_L g5167 ( 
.A1(n_5024),
.A2(n_4510),
.B1(n_4518),
.B2(n_4500),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_4879),
.Y(n_5168)
);

OAI21x1_ASAP7_75t_L g5169 ( 
.A1(n_4972),
.A2(n_4608),
.B(n_4236),
.Y(n_5169)
);

OAI21x1_ASAP7_75t_L g5170 ( 
.A1(n_4999),
.A2(n_4231),
.B(n_4430),
.Y(n_5170)
);

CKINVDCx20_ASAP7_75t_R g5171 ( 
.A(n_4755),
.Y(n_5171)
);

BUFx3_ASAP7_75t_L g5172 ( 
.A(n_4655),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_4812),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_4831),
.Y(n_5174)
);

NOR2x1_ASAP7_75t_SL g5175 ( 
.A(n_4692),
.B(n_4719),
.Y(n_5175)
);

AND2x4_ASAP7_75t_L g5176 ( 
.A(n_4845),
.B(n_4176),
.Y(n_5176)
);

OAI21x1_ASAP7_75t_L g5177 ( 
.A1(n_5091),
.A2(n_4266),
.B(n_4258),
.Y(n_5177)
);

AND2x4_ASAP7_75t_L g5178 ( 
.A(n_4866),
.B(n_4486),
.Y(n_5178)
);

OAI22xp33_ASAP7_75t_L g5179 ( 
.A1(n_4700),
.A2(n_4591),
.B1(n_4568),
.B2(n_4593),
.Y(n_5179)
);

BUFx6f_ASAP7_75t_L g5180 ( 
.A(n_4636),
.Y(n_5180)
);

OAI21x1_ASAP7_75t_L g5181 ( 
.A1(n_4952),
.A2(n_4463),
.B(n_4604),
.Y(n_5181)
);

A2O1A1Ixp33_ASAP7_75t_L g5182 ( 
.A1(n_4855),
.A2(n_4352),
.B(n_4442),
.C(n_4398),
.Y(n_5182)
);

AND2x4_ASAP7_75t_L g5183 ( 
.A(n_4706),
.B(n_4501),
.Y(n_5183)
);

OAI21x1_ASAP7_75t_L g5184 ( 
.A1(n_5071),
.A2(n_4607),
.B(n_4315),
.Y(n_5184)
);

AO21x2_ASAP7_75t_L g5185 ( 
.A1(n_5027),
.A2(n_4238),
.B(n_4237),
.Y(n_5185)
);

INVx2_ASAP7_75t_L g5186 ( 
.A(n_4723),
.Y(n_5186)
);

OAI21x1_ASAP7_75t_L g5187 ( 
.A1(n_5087),
.A2(n_4191),
.B(n_4545),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_4890),
.B(n_4554),
.Y(n_5188)
);

CKINVDCx5p33_ASAP7_75t_R g5189 ( 
.A(n_4789),
.Y(n_5189)
);

AOI211xp5_ASAP7_75t_L g5190 ( 
.A1(n_4818),
.A2(n_4561),
.B(n_4186),
.C(n_4259),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_4848),
.Y(n_5191)
);

NAND3xp33_ASAP7_75t_L g5192 ( 
.A(n_5074),
.B(n_4508),
.C(n_4506),
.Y(n_5192)
);

OAI21x1_ASAP7_75t_L g5193 ( 
.A1(n_4772),
.A2(n_4553),
.B(n_4551),
.Y(n_5193)
);

OAI21x1_ASAP7_75t_L g5194 ( 
.A1(n_5088),
.A2(n_4557),
.B(n_4460),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_L g5195 ( 
.A(n_4887),
.B(n_4255),
.Y(n_5195)
);

OR2x2_ASAP7_75t_L g5196 ( 
.A(n_4710),
.B(n_607),
.Y(n_5196)
);

OA21x2_ASAP7_75t_L g5197 ( 
.A1(n_4983),
.A2(n_4594),
.B(n_4587),
.Y(n_5197)
);

AO31x2_ASAP7_75t_L g5198 ( 
.A1(n_4988),
.A2(n_4609),
.A3(n_4573),
.B(n_4566),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_L g5199 ( 
.A(n_4849),
.B(n_4262),
.Y(n_5199)
);

AOI222xp33_ASAP7_75t_L g5200 ( 
.A1(n_4703),
.A2(n_4418),
.B1(n_4558),
.B2(n_4564),
.C1(n_4548),
.C2(n_4285),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_4864),
.Y(n_5201)
);

OAI21x1_ASAP7_75t_L g5202 ( 
.A1(n_5097),
.A2(n_4491),
.B(n_4469),
.Y(n_5202)
);

NOR2xp33_ASAP7_75t_L g5203 ( 
.A(n_4676),
.B(n_607),
.Y(n_5203)
);

INVx4_ASAP7_75t_L g5204 ( 
.A(n_4688),
.Y(n_5204)
);

OAI221xp5_ASAP7_75t_L g5205 ( 
.A1(n_4698),
.A2(n_4265),
.B1(n_4445),
.B2(n_4304),
.C(n_4595),
.Y(n_5205)
);

OAI22xp5_ASAP7_75t_L g5206 ( 
.A1(n_4728),
.A2(n_4507),
.B1(n_4574),
.B2(n_4569),
.Y(n_5206)
);

AOI21x1_ASAP7_75t_L g5207 ( 
.A1(n_4647),
.A2(n_608),
.B(n_609),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_4877),
.Y(n_5208)
);

INVx3_ASAP7_75t_L g5209 ( 
.A(n_4657),
.Y(n_5209)
);

OAI21x1_ASAP7_75t_L g5210 ( 
.A1(n_4941),
.A2(n_851),
.B(n_850),
.Y(n_5210)
);

OAI21x1_ASAP7_75t_L g5211 ( 
.A1(n_4961),
.A2(n_853),
.B(n_852),
.Y(n_5211)
);

INVx3_ASAP7_75t_L g5212 ( 
.A(n_4634),
.Y(n_5212)
);

NOR2xp33_ASAP7_75t_L g5213 ( 
.A(n_4676),
.B(n_608),
.Y(n_5213)
);

CKINVDCx5p33_ASAP7_75t_R g5214 ( 
.A(n_4641),
.Y(n_5214)
);

BUFx2_ASAP7_75t_L g5215 ( 
.A(n_4884),
.Y(n_5215)
);

INVx4_ASAP7_75t_L g5216 ( 
.A(n_4694),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_4891),
.B(n_608),
.Y(n_5217)
);

BUFx2_ASAP7_75t_R g5218 ( 
.A(n_4697),
.Y(n_5218)
);

OAI22xp5_ASAP7_75t_R g5219 ( 
.A1(n_4675),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.Y(n_5219)
);

NOR2xp33_ASAP7_75t_L g5220 ( 
.A(n_4843),
.B(n_4665),
.Y(n_5220)
);

OAI21x1_ASAP7_75t_L g5221 ( 
.A1(n_5028),
.A2(n_853),
.B(n_852),
.Y(n_5221)
);

INVx2_ASAP7_75t_L g5222 ( 
.A(n_4733),
.Y(n_5222)
);

INVx2_ASAP7_75t_L g5223 ( 
.A(n_4740),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_4673),
.B(n_4677),
.Y(n_5224)
);

NAND2x1p5_ASAP7_75t_L g5225 ( 
.A(n_4694),
.B(n_610),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4935),
.Y(n_5226)
);

AND2x2_ASAP7_75t_L g5227 ( 
.A(n_4727),
.B(n_611),
.Y(n_5227)
);

AOI22x1_ASAP7_75t_L g5228 ( 
.A1(n_4687),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.Y(n_5228)
);

OAI21x1_ASAP7_75t_L g5229 ( 
.A1(n_4644),
.A2(n_855),
.B(n_854),
.Y(n_5229)
);

OAI21x1_ASAP7_75t_L g5230 ( 
.A1(n_4660),
.A2(n_857),
.B(n_855),
.Y(n_5230)
);

CKINVDCx8_ASAP7_75t_R g5231 ( 
.A(n_4638),
.Y(n_5231)
);

INVx3_ASAP7_75t_L g5232 ( 
.A(n_4642),
.Y(n_5232)
);

AND2x2_ASAP7_75t_L g5233 ( 
.A(n_4712),
.B(n_4937),
.Y(n_5233)
);

OAI21x1_ASAP7_75t_L g5234 ( 
.A1(n_4968),
.A2(n_858),
.B(n_857),
.Y(n_5234)
);

NAND2x1p5_ASAP7_75t_L g5235 ( 
.A(n_4695),
.B(n_612),
.Y(n_5235)
);

INVx2_ASAP7_75t_L g5236 ( 
.A(n_4749),
.Y(n_5236)
);

INVx2_ASAP7_75t_SL g5237 ( 
.A(n_4658),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_4764),
.Y(n_5238)
);

OR2x6_ASAP7_75t_L g5239 ( 
.A(n_4800),
.B(n_612),
.Y(n_5239)
);

BUFx3_ASAP7_75t_L g5240 ( 
.A(n_4643),
.Y(n_5240)
);

CKINVDCx16_ASAP7_75t_R g5241 ( 
.A(n_4699),
.Y(n_5241)
);

INVx1_ASAP7_75t_L g5242 ( 
.A(n_4678),
.Y(n_5242)
);

OA21x2_ASAP7_75t_L g5243 ( 
.A1(n_4992),
.A2(n_613),
.B(n_614),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_4754),
.Y(n_5244)
);

OAI21xp5_ASAP7_75t_L g5245 ( 
.A1(n_4739),
.A2(n_613),
.B(n_614),
.Y(n_5245)
);

INVx6_ASAP7_75t_L g5246 ( 
.A(n_4695),
.Y(n_5246)
);

OAI21x1_ASAP7_75t_L g5247 ( 
.A1(n_4977),
.A2(n_860),
.B(n_859),
.Y(n_5247)
);

BUFx3_ASAP7_75t_L g5248 ( 
.A(n_4643),
.Y(n_5248)
);

AND2x2_ASAP7_75t_L g5249 ( 
.A(n_4876),
.B(n_615),
.Y(n_5249)
);

AOI22xp5_ASAP7_75t_L g5250 ( 
.A1(n_5035),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_5250)
);

OAI21xp33_ASAP7_75t_SL g5251 ( 
.A1(n_4837),
.A2(n_615),
.B(n_616),
.Y(n_5251)
);

INVxp67_ASAP7_75t_L g5252 ( 
.A(n_4853),
.Y(n_5252)
);

INVx3_ASAP7_75t_L g5253 ( 
.A(n_4730),
.Y(n_5253)
);

OAI21xp5_ASAP7_75t_L g5254 ( 
.A1(n_5006),
.A2(n_4809),
.B(n_5010),
.Y(n_5254)
);

O2A1O1Ixp33_ASAP7_75t_SL g5255 ( 
.A1(n_4862),
.A2(n_4662),
.B(n_4850),
.C(n_4646),
.Y(n_5255)
);

AND2x2_ASAP7_75t_L g5256 ( 
.A(n_4905),
.B(n_616),
.Y(n_5256)
);

OAI21x1_ASAP7_75t_L g5257 ( 
.A1(n_5081),
.A2(n_860),
.B(n_859),
.Y(n_5257)
);

INVx5_ASAP7_75t_SL g5258 ( 
.A(n_4829),
.Y(n_5258)
);

INVx1_ASAP7_75t_L g5259 ( 
.A(n_4683),
.Y(n_5259)
);

AO21x2_ASAP7_75t_L g5260 ( 
.A1(n_5027),
.A2(n_617),
.B(n_618),
.Y(n_5260)
);

AND2x4_ASAP7_75t_L g5261 ( 
.A(n_4649),
.B(n_617),
.Y(n_5261)
);

INVx2_ASAP7_75t_L g5262 ( 
.A(n_4685),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_4691),
.Y(n_5263)
);

AOI22xp33_ASAP7_75t_L g5264 ( 
.A1(n_5051),
.A2(n_620),
.B1(n_618),
.B2(n_619),
.Y(n_5264)
);

OAI21x1_ASAP7_75t_L g5265 ( 
.A1(n_4704),
.A2(n_862),
.B(n_861),
.Y(n_5265)
);

AOI22xp33_ASAP7_75t_L g5266 ( 
.A1(n_5051),
.A2(n_620),
.B1(n_618),
.B2(n_619),
.Y(n_5266)
);

NAND2x1p5_ASAP7_75t_L g5267 ( 
.A(n_4640),
.B(n_620),
.Y(n_5267)
);

AOI21xp5_ASAP7_75t_L g5268 ( 
.A1(n_4994),
.A2(n_621),
.B(n_622),
.Y(n_5268)
);

HB1xp67_ASAP7_75t_L g5269 ( 
.A(n_4830),
.Y(n_5269)
);

AO21x2_ASAP7_75t_L g5270 ( 
.A1(n_4750),
.A2(n_622),
.B(n_623),
.Y(n_5270)
);

AOI22xp33_ASAP7_75t_L g5271 ( 
.A1(n_4980),
.A2(n_625),
.B1(n_623),
.B2(n_624),
.Y(n_5271)
);

INVx3_ASAP7_75t_L g5272 ( 
.A(n_4684),
.Y(n_5272)
);

OAI21xp5_ASAP7_75t_L g5273 ( 
.A1(n_4784),
.A2(n_624),
.B(n_625),
.Y(n_5273)
);

NOR2xp33_ASAP7_75t_L g5274 ( 
.A(n_4940),
.B(n_624),
.Y(n_5274)
);

OR2x2_ASAP7_75t_L g5275 ( 
.A(n_4803),
.B(n_625),
.Y(n_5275)
);

HB1xp67_ASAP7_75t_L g5276 ( 
.A(n_4830),
.Y(n_5276)
);

INVx2_ASAP7_75t_L g5277 ( 
.A(n_4717),
.Y(n_5277)
);

BUFx3_ASAP7_75t_L g5278 ( 
.A(n_4681),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_4720),
.Y(n_5279)
);

INVx2_ASAP7_75t_L g5280 ( 
.A(n_4746),
.Y(n_5280)
);

AOI222xp33_ASAP7_75t_L g5281 ( 
.A1(n_4991),
.A2(n_628),
.B1(n_631),
.B2(n_626),
.C1(n_627),
.C2(n_630),
.Y(n_5281)
);

OR2x6_ASAP7_75t_L g5282 ( 
.A(n_4800),
.B(n_626),
.Y(n_5282)
);

AO21x2_ASAP7_75t_L g5283 ( 
.A1(n_4916),
.A2(n_626),
.B(n_627),
.Y(n_5283)
);

AOI21xp5_ASAP7_75t_L g5284 ( 
.A1(n_5013),
.A2(n_628),
.B(n_630),
.Y(n_5284)
);

NOR2x1_ASAP7_75t_SL g5285 ( 
.A(n_4868),
.B(n_630),
.Y(n_5285)
);

NAND2xp5_ASAP7_75t_L g5286 ( 
.A(n_4747),
.B(n_631),
.Y(n_5286)
);

AOI22xp5_ASAP7_75t_SL g5287 ( 
.A1(n_4670),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.Y(n_5287)
);

OR2x2_ASAP7_75t_L g5288 ( 
.A(n_4803),
.B(n_632),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_4690),
.Y(n_5289)
);

AOI21xp5_ASAP7_75t_L g5290 ( 
.A1(n_5082),
.A2(n_4910),
.B(n_4908),
.Y(n_5290)
);

OAI21x1_ASAP7_75t_L g5291 ( 
.A1(n_4949),
.A2(n_5009),
.B(n_4769),
.Y(n_5291)
);

AO31x2_ASAP7_75t_L g5292 ( 
.A1(n_4958),
.A2(n_634),
.A3(n_632),
.B(n_633),
.Y(n_5292)
);

OAI21x1_ASAP7_75t_L g5293 ( 
.A1(n_4915),
.A2(n_862),
.B(n_861),
.Y(n_5293)
);

BUFx3_ASAP7_75t_L g5294 ( 
.A(n_4682),
.Y(n_5294)
);

HB1xp67_ASAP7_75t_L g5295 ( 
.A(n_4779),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4790),
.Y(n_5296)
);

INVx5_ASAP7_75t_L g5297 ( 
.A(n_4859),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_4765),
.Y(n_5298)
);

OAI21x1_ASAP7_75t_L g5299 ( 
.A1(n_4788),
.A2(n_864),
.B(n_863),
.Y(n_5299)
);

A2O1A1Ixp33_ASAP7_75t_L g5300 ( 
.A1(n_4888),
.A2(n_637),
.B(n_635),
.C(n_636),
.Y(n_5300)
);

OR2x6_ASAP7_75t_L g5301 ( 
.A(n_4888),
.B(n_635),
.Y(n_5301)
);

AO21x2_ASAP7_75t_L g5302 ( 
.A1(n_4916),
.A2(n_635),
.B(n_636),
.Y(n_5302)
);

INVx2_ASAP7_75t_L g5303 ( 
.A(n_4731),
.Y(n_5303)
);

AOI21xp5_ASAP7_75t_L g5304 ( 
.A1(n_4910),
.A2(n_636),
.B(n_637),
.Y(n_5304)
);

CKINVDCx20_ASAP7_75t_R g5305 ( 
.A(n_4631),
.Y(n_5305)
);

INVx3_ASAP7_75t_L g5306 ( 
.A(n_4729),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_4770),
.Y(n_5307)
);

AO21x2_ASAP7_75t_L g5308 ( 
.A1(n_4763),
.A2(n_637),
.B(n_638),
.Y(n_5308)
);

OAI21x1_ASAP7_75t_L g5309 ( 
.A1(n_4987),
.A2(n_865),
.B(n_863),
.Y(n_5309)
);

OAI21x1_ASAP7_75t_L g5310 ( 
.A1(n_4987),
.A2(n_866),
.B(n_865),
.Y(n_5310)
);

OAI21x1_ASAP7_75t_L g5311 ( 
.A1(n_5007),
.A2(n_868),
.B(n_867),
.Y(n_5311)
);

AO21x2_ASAP7_75t_L g5312 ( 
.A1(n_4721),
.A2(n_638),
.B(n_639),
.Y(n_5312)
);

INVx2_ASAP7_75t_L g5313 ( 
.A(n_4731),
.Y(n_5313)
);

OAI21x1_ASAP7_75t_L g5314 ( 
.A1(n_5007),
.A2(n_868),
.B(n_867),
.Y(n_5314)
);

OA21x2_ASAP7_75t_L g5315 ( 
.A1(n_4998),
.A2(n_638),
.B(n_639),
.Y(n_5315)
);

OR2x6_ASAP7_75t_L g5316 ( 
.A(n_4847),
.B(n_639),
.Y(n_5316)
);

BUFx8_ASAP7_75t_SL g5317 ( 
.A(n_4661),
.Y(n_5317)
);

NOR2xp33_ASAP7_75t_L g5318 ( 
.A(n_4637),
.B(n_640),
.Y(n_5318)
);

NAND2x1p5_ASAP7_75t_L g5319 ( 
.A(n_4716),
.B(n_640),
.Y(n_5319)
);

OAI21xp5_ASAP7_75t_L g5320 ( 
.A1(n_4856),
.A2(n_640),
.B(n_641),
.Y(n_5320)
);

OAI21x1_ASAP7_75t_L g5321 ( 
.A1(n_4954),
.A2(n_870),
.B(n_869),
.Y(n_5321)
);

NOR2xp33_ASAP7_75t_SL g5322 ( 
.A(n_4705),
.B(n_641),
.Y(n_5322)
);

OA21x2_ASAP7_75t_L g5323 ( 
.A1(n_5093),
.A2(n_641),
.B(n_642),
.Y(n_5323)
);

AND2x2_ASAP7_75t_L g5324 ( 
.A(n_4664),
.B(n_642),
.Y(n_5324)
);

OAI21x1_ASAP7_75t_L g5325 ( 
.A1(n_5085),
.A2(n_871),
.B(n_869),
.Y(n_5325)
);

INVx2_ASAP7_75t_L g5326 ( 
.A(n_4736),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_4792),
.Y(n_5327)
);

AND2x4_ASAP7_75t_L g5328 ( 
.A(n_4844),
.B(n_643),
.Y(n_5328)
);

AOI21x1_ASAP7_75t_L g5329 ( 
.A1(n_4711),
.A2(n_643),
.B(n_644),
.Y(n_5329)
);

NAND2xp5_ASAP7_75t_L g5330 ( 
.A(n_4841),
.B(n_644),
.Y(n_5330)
);

INVx2_ASAP7_75t_L g5331 ( 
.A(n_4736),
.Y(n_5331)
);

OAI21x1_ASAP7_75t_L g5332 ( 
.A1(n_5068),
.A2(n_5098),
.B(n_4852),
.Y(n_5332)
);

NAND2xp5_ASAP7_75t_L g5333 ( 
.A(n_4841),
.B(n_644),
.Y(n_5333)
);

OAI21x1_ASAP7_75t_L g5334 ( 
.A1(n_4838),
.A2(n_872),
.B(n_871),
.Y(n_5334)
);

NAND3xp33_ASAP7_75t_L g5335 ( 
.A(n_5076),
.B(n_645),
.C(n_646),
.Y(n_5335)
);

BUFx2_ASAP7_75t_L g5336 ( 
.A(n_4957),
.Y(n_5336)
);

NOR2xp33_ASAP7_75t_SL g5337 ( 
.A(n_4713),
.B(n_645),
.Y(n_5337)
);

BUFx6f_ASAP7_75t_L g5338 ( 
.A(n_4816),
.Y(n_5338)
);

AOI21xp5_ASAP7_75t_L g5339 ( 
.A1(n_4908),
.A2(n_645),
.B(n_647),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_4775),
.Y(n_5340)
);

AOI22xp33_ASAP7_75t_L g5341 ( 
.A1(n_4980),
.A2(n_649),
.B1(n_647),
.B2(n_648),
.Y(n_5341)
);

OAI21xp5_ASAP7_75t_L g5342 ( 
.A1(n_4651),
.A2(n_648),
.B(n_649),
.Y(n_5342)
);

CKINVDCx11_ASAP7_75t_R g5343 ( 
.A(n_4686),
.Y(n_5343)
);

OAI21x1_ASAP7_75t_L g5344 ( 
.A1(n_4865),
.A2(n_873),
.B(n_872),
.Y(n_5344)
);

HB1xp67_ASAP7_75t_L g5345 ( 
.A(n_4791),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_4785),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4883),
.Y(n_5347)
);

BUFx2_ASAP7_75t_L g5348 ( 
.A(n_4899),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_4817),
.Y(n_5349)
);

OAI21x1_ASAP7_75t_SL g5350 ( 
.A1(n_4707),
.A2(n_648),
.B(n_649),
.Y(n_5350)
);

OAI21x1_ASAP7_75t_L g5351 ( 
.A1(n_4914),
.A2(n_876),
.B(n_875),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5043),
.Y(n_5352)
);

OAI21xp5_ASAP7_75t_L g5353 ( 
.A1(n_4931),
.A2(n_650),
.B(n_651),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_L g5354 ( 
.A(n_4797),
.B(n_650),
.Y(n_5354)
);

BUFx2_ASAP7_75t_SL g5355 ( 
.A(n_4716),
.Y(n_5355)
);

INVx2_ASAP7_75t_L g5356 ( 
.A(n_4970),
.Y(n_5356)
);

INVx2_ASAP7_75t_L g5357 ( 
.A(n_4970),
.Y(n_5357)
);

OAI21x1_ASAP7_75t_L g5358 ( 
.A1(n_4982),
.A2(n_877),
.B(n_876),
.Y(n_5358)
);

HB1xp67_ASAP7_75t_L g5359 ( 
.A(n_4780),
.Y(n_5359)
);

AOI22xp5_ASAP7_75t_L g5360 ( 
.A1(n_4921),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.Y(n_5360)
);

OAI21x1_ASAP7_75t_L g5361 ( 
.A1(n_5038),
.A2(n_878),
.B(n_877),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4771),
.Y(n_5362)
);

NAND2xp5_ASAP7_75t_SL g5363 ( 
.A(n_4829),
.B(n_651),
.Y(n_5363)
);

AOI21xp5_ASAP7_75t_L g5364 ( 
.A1(n_4810),
.A2(n_652),
.B(n_653),
.Y(n_5364)
);

NAND2xp5_ASAP7_75t_SL g5365 ( 
.A(n_4728),
.B(n_652),
.Y(n_5365)
);

AOI21xp5_ASAP7_75t_L g5366 ( 
.A1(n_4811),
.A2(n_653),
.B(n_654),
.Y(n_5366)
);

AOI21xp5_ASAP7_75t_L g5367 ( 
.A1(n_4815),
.A2(n_653),
.B(n_654),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_4783),
.Y(n_5368)
);

OAI21x1_ASAP7_75t_L g5369 ( 
.A1(n_4767),
.A2(n_879),
.B(n_878),
.Y(n_5369)
);

OAI22xp5_ASAP7_75t_L g5370 ( 
.A1(n_4857),
.A2(n_656),
.B1(n_654),
.B2(n_655),
.Y(n_5370)
);

OR2x2_ASAP7_75t_L g5371 ( 
.A(n_4805),
.B(n_4630),
.Y(n_5371)
);

NOR2xp33_ASAP7_75t_L g5372 ( 
.A(n_4928),
.B(n_656),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_4745),
.Y(n_5373)
);

OAI21x1_ASAP7_75t_L g5374 ( 
.A1(n_4943),
.A2(n_4939),
.B(n_4971),
.Y(n_5374)
);

AND2x2_ASAP7_75t_L g5375 ( 
.A(n_4861),
.B(n_656),
.Y(n_5375)
);

BUFx3_ASAP7_75t_L g5376 ( 
.A(n_4828),
.Y(n_5376)
);

NAND2xp5_ASAP7_75t_L g5377 ( 
.A(n_4799),
.B(n_657),
.Y(n_5377)
);

AND2x4_ASAP7_75t_L g5378 ( 
.A(n_4732),
.B(n_657),
.Y(n_5378)
);

INVx1_ASAP7_75t_L g5379 ( 
.A(n_5011),
.Y(n_5379)
);

HB1xp67_ASAP7_75t_L g5380 ( 
.A(n_4832),
.Y(n_5380)
);

OR2x2_ASAP7_75t_L g5381 ( 
.A(n_4900),
.B(n_657),
.Y(n_5381)
);

AND2x2_ASAP7_75t_L g5382 ( 
.A(n_4942),
.B(n_658),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_5014),
.Y(n_5383)
);

OAI21x1_ASAP7_75t_L g5384 ( 
.A1(n_4768),
.A2(n_880),
.B(n_879),
.Y(n_5384)
);

OR2x2_ASAP7_75t_L g5385 ( 
.A(n_4786),
.B(n_658),
.Y(n_5385)
);

INVx2_ASAP7_75t_L g5386 ( 
.A(n_4974),
.Y(n_5386)
);

AND2x2_ASAP7_75t_L g5387 ( 
.A(n_4948),
.B(n_659),
.Y(n_5387)
);

OAI21x1_ASAP7_75t_L g5388 ( 
.A1(n_5029),
.A2(n_882),
.B(n_881),
.Y(n_5388)
);

OAI221xp5_ASAP7_75t_L g5389 ( 
.A1(n_4628),
.A2(n_661),
.B1(n_659),
.B2(n_660),
.C(n_662),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_4808),
.B(n_659),
.Y(n_5390)
);

OA21x2_ASAP7_75t_L g5391 ( 
.A1(n_5086),
.A2(n_660),
.B(n_661),
.Y(n_5391)
);

BUFx3_ASAP7_75t_L g5392 ( 
.A(n_4671),
.Y(n_5392)
);

BUFx3_ASAP7_75t_L g5393 ( 
.A(n_4672),
.Y(n_5393)
);

AO31x2_ASAP7_75t_L g5394 ( 
.A1(n_5092),
.A2(n_663),
.A3(n_661),
.B(n_662),
.Y(n_5394)
);

OAI21x1_ASAP7_75t_L g5395 ( 
.A1(n_4726),
.A2(n_882),
.B(n_881),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_5022),
.Y(n_5396)
);

INVx3_ASAP7_75t_L g5397 ( 
.A(n_4631),
.Y(n_5397)
);

AO21x2_ASAP7_75t_L g5398 ( 
.A1(n_4985),
.A2(n_662),
.B(n_663),
.Y(n_5398)
);

OAI21x1_ASAP7_75t_L g5399 ( 
.A1(n_4820),
.A2(n_884),
.B(n_883),
.Y(n_5399)
);

OAI21x1_ASAP7_75t_L g5400 ( 
.A1(n_4680),
.A2(n_886),
.B(n_885),
.Y(n_5400)
);

INVx2_ASAP7_75t_L g5401 ( 
.A(n_4974),
.Y(n_5401)
);

OAI21x1_ASAP7_75t_L g5402 ( 
.A1(n_5040),
.A2(n_886),
.B(n_885),
.Y(n_5402)
);

BUFx6f_ASAP7_75t_L g5403 ( 
.A(n_4672),
.Y(n_5403)
);

OA21x2_ASAP7_75t_L g5404 ( 
.A1(n_5095),
.A2(n_663),
.B(n_664),
.Y(n_5404)
);

OAI21x1_ASAP7_75t_L g5405 ( 
.A1(n_5040),
.A2(n_891),
.B(n_890),
.Y(n_5405)
);

INVx2_ASAP7_75t_L g5406 ( 
.A(n_5004),
.Y(n_5406)
);

OAI21x1_ASAP7_75t_L g5407 ( 
.A1(n_5049),
.A2(n_891),
.B(n_890),
.Y(n_5407)
);

AOI211x1_ASAP7_75t_L g5408 ( 
.A1(n_4951),
.A2(n_667),
.B(n_665),
.C(n_666),
.Y(n_5408)
);

NAND2xp5_ASAP7_75t_L g5409 ( 
.A(n_4823),
.B(n_666),
.Y(n_5409)
);

AOI22xp33_ASAP7_75t_L g5410 ( 
.A1(n_5083),
.A2(n_668),
.B1(n_666),
.B2(n_667),
.Y(n_5410)
);

O2A1O1Ixp33_ASAP7_75t_L g5411 ( 
.A1(n_5060),
.A2(n_670),
.B(n_668),
.C(n_669),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_5039),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_5055),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_5352),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5103),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5110),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5111),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5140),
.Y(n_5418)
);

INVx5_ASAP7_75t_L g5419 ( 
.A(n_5246),
.Y(n_5419)
);

NAND2xp5_ASAP7_75t_L g5420 ( 
.A(n_5346),
.B(n_5058),
.Y(n_5420)
);

AND2x2_ASAP7_75t_L g5421 ( 
.A(n_5118),
.B(n_4758),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_5143),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_5379),
.B(n_4962),
.Y(n_5423)
);

AOI22xp33_ASAP7_75t_SL g5424 ( 
.A1(n_5345),
.A2(n_4872),
.B1(n_4835),
.B2(n_5048),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5145),
.Y(n_5425)
);

INVx2_ASAP7_75t_L g5426 ( 
.A(n_5111),
.Y(n_5426)
);

INVx1_ASAP7_75t_L g5427 ( 
.A(n_5147),
.Y(n_5427)
);

INVx2_ASAP7_75t_L g5428 ( 
.A(n_5128),
.Y(n_5428)
);

CKINVDCx20_ASAP7_75t_R g5429 ( 
.A(n_5171),
.Y(n_5429)
);

OAI221xp5_ASAP7_75t_L g5430 ( 
.A1(n_5122),
.A2(n_4667),
.B1(n_4897),
.B2(n_5023),
.C(n_4860),
.Y(n_5430)
);

BUFx2_ASAP7_75t_L g5431 ( 
.A(n_5348),
.Y(n_5431)
);

INVx2_ASAP7_75t_L g5432 ( 
.A(n_5163),
.Y(n_5432)
);

INVx3_ASAP7_75t_SL g5433 ( 
.A(n_5297),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_5149),
.Y(n_5434)
);

OAI21x1_ASAP7_75t_SL g5435 ( 
.A1(n_5175),
.A2(n_5285),
.B(n_5254),
.Y(n_5435)
);

NAND2xp5_ASAP7_75t_L g5436 ( 
.A(n_5383),
.B(n_4963),
.Y(n_5436)
);

OA21x2_ASAP7_75t_L g5437 ( 
.A1(n_5290),
.A2(n_4985),
.B(n_4840),
.Y(n_5437)
);

INVx3_ASAP7_75t_L g5438 ( 
.A(n_5231),
.Y(n_5438)
);

AND2x4_ASAP7_75t_L g5439 ( 
.A(n_5233),
.B(n_4737),
.Y(n_5439)
);

BUFx4f_ASAP7_75t_SL g5440 ( 
.A(n_5305),
.Y(n_5440)
);

BUFx6f_ASAP7_75t_L g5441 ( 
.A(n_5278),
.Y(n_5441)
);

AOI22xp5_ASAP7_75t_L g5442 ( 
.A1(n_5179),
.A2(n_5031),
.B1(n_4885),
.B2(n_4893),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5150),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_5396),
.B(n_4995),
.Y(n_5444)
);

AOI21x1_ASAP7_75t_L g5445 ( 
.A1(n_5243),
.A2(n_4895),
.B(n_4654),
.Y(n_5445)
);

INVx2_ASAP7_75t_L g5446 ( 
.A(n_5186),
.Y(n_5446)
);

INVx1_ASAP7_75t_L g5447 ( 
.A(n_5412),
.Y(n_5447)
);

AND2x2_ASAP7_75t_L g5448 ( 
.A(n_5269),
.B(n_4756),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5413),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5327),
.Y(n_5450)
);

INVx1_ASAP7_75t_L g5451 ( 
.A(n_5298),
.Y(n_5451)
);

INVx1_ASAP7_75t_L g5452 ( 
.A(n_5307),
.Y(n_5452)
);

INVx2_ASAP7_75t_L g5453 ( 
.A(n_5222),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_5242),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_5259),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_5263),
.Y(n_5456)
);

BUFx2_ASAP7_75t_L g5457 ( 
.A(n_5348),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_5223),
.Y(n_5458)
);

INVxp67_ASAP7_75t_L g5459 ( 
.A(n_5276),
.Y(n_5459)
);

AO21x2_ASAP7_75t_L g5460 ( 
.A1(n_5291),
.A2(n_4787),
.B(n_4757),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5279),
.Y(n_5461)
);

INVx2_ASAP7_75t_L g5462 ( 
.A(n_5236),
.Y(n_5462)
);

INVx1_ASAP7_75t_L g5463 ( 
.A(n_5296),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_5262),
.Y(n_5464)
);

INVx2_ASAP7_75t_L g5465 ( 
.A(n_5238),
.Y(n_5465)
);

INVx2_ASAP7_75t_SL g5466 ( 
.A(n_5297),
.Y(n_5466)
);

AOI22xp33_ASAP7_75t_L g5467 ( 
.A1(n_5123),
.A2(n_5037),
.B1(n_5000),
.B2(n_5076),
.Y(n_5467)
);

AND2x4_ASAP7_75t_L g5468 ( 
.A(n_5146),
.B(n_4832),
.Y(n_5468)
);

NAND2xp5_ASAP7_75t_L g5469 ( 
.A(n_5303),
.B(n_5026),
.Y(n_5469)
);

AND2x4_ASAP7_75t_L g5470 ( 
.A(n_5215),
.B(n_4722),
.Y(n_5470)
);

BUFx2_ASAP7_75t_L g5471 ( 
.A(n_5138),
.Y(n_5471)
);

AOI22xp33_ASAP7_75t_L g5472 ( 
.A1(n_5116),
.A2(n_5077),
.B1(n_4929),
.B2(n_4934),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_5277),
.Y(n_5473)
);

OAI21xp5_ASAP7_75t_L g5474 ( 
.A1(n_5251),
.A2(n_4709),
.B(n_4760),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_5280),
.Y(n_5475)
);

INVx4_ASAP7_75t_L g5476 ( 
.A(n_5297),
.Y(n_5476)
);

OAI21x1_ASAP7_75t_L g5477 ( 
.A1(n_5107),
.A2(n_5106),
.B(n_5112),
.Y(n_5477)
);

INVx4_ASAP7_75t_L g5478 ( 
.A(n_5204),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5168),
.Y(n_5479)
);

CKINVDCx5p33_ASAP7_75t_R g5480 ( 
.A(n_5189),
.Y(n_5480)
);

INVx4_ASAP7_75t_SL g5481 ( 
.A(n_5246),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5224),
.Y(n_5482)
);

BUFx2_ASAP7_75t_R g5483 ( 
.A(n_5172),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_5289),
.Y(n_5484)
);

INVx3_ASAP7_75t_L g5485 ( 
.A(n_5216),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5156),
.Y(n_5486)
);

HB1xp67_ASAP7_75t_L g5487 ( 
.A(n_5295),
.Y(n_5487)
);

HB1xp67_ASAP7_75t_L g5488 ( 
.A(n_5359),
.Y(n_5488)
);

NAND2x1p5_ASAP7_75t_L g5489 ( 
.A(n_5253),
.B(n_5272),
.Y(n_5489)
);

CKINVDCx5p33_ASAP7_75t_R g5490 ( 
.A(n_5343),
.Y(n_5490)
);

BUFx3_ASAP7_75t_L g5491 ( 
.A(n_5148),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5173),
.Y(n_5492)
);

AND2x2_ASAP7_75t_L g5493 ( 
.A(n_5226),
.B(n_5077),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_5347),
.Y(n_5494)
);

INVx2_ASAP7_75t_L g5495 ( 
.A(n_5174),
.Y(n_5495)
);

OAI221xp5_ASAP7_75t_L g5496 ( 
.A1(n_5250),
.A2(n_5050),
.B1(n_5047),
.B2(n_4715),
.C(n_5036),
.Y(n_5496)
);

INVx2_ASAP7_75t_L g5497 ( 
.A(n_5191),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5201),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5208),
.Y(n_5499)
);

AOI21x1_ASAP7_75t_L g5500 ( 
.A1(n_5243),
.A2(n_4895),
.B(n_4708),
.Y(n_5500)
);

INVx3_ASAP7_75t_L g5501 ( 
.A(n_5338),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_5349),
.Y(n_5502)
);

INVx2_ASAP7_75t_L g5503 ( 
.A(n_5356),
.Y(n_5503)
);

INVx3_ASAP7_75t_L g5504 ( 
.A(n_5338),
.Y(n_5504)
);

AND2x4_ASAP7_75t_L g5505 ( 
.A(n_5215),
.B(n_4702),
.Y(n_5505)
);

AO21x1_ASAP7_75t_L g5506 ( 
.A1(n_5261),
.A2(n_4766),
.B(n_4826),
.Y(n_5506)
);

INVx2_ASAP7_75t_SL g5507 ( 
.A(n_5101),
.Y(n_5507)
);

INVx3_ASAP7_75t_L g5508 ( 
.A(n_5294),
.Y(n_5508)
);

AOI22xp33_ASAP7_75t_SL g5509 ( 
.A1(n_5287),
.A2(n_4777),
.B1(n_4742),
.B2(n_4975),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_5357),
.Y(n_5510)
);

BUFx3_ASAP7_75t_L g5511 ( 
.A(n_5102),
.Y(n_5511)
);

INVx2_ASAP7_75t_SL g5512 ( 
.A(n_5240),
.Y(n_5512)
);

A2O1A1Ixp33_ASAP7_75t_L g5513 ( 
.A1(n_5300),
.A2(n_4945),
.B(n_4724),
.C(n_4894),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_5340),
.Y(n_5514)
);

CKINVDCx5p33_ASAP7_75t_R g5515 ( 
.A(n_5214),
.Y(n_5515)
);

INVx2_ASAP7_75t_L g5516 ( 
.A(n_5386),
.Y(n_5516)
);

BUFx3_ASAP7_75t_L g5517 ( 
.A(n_5306),
.Y(n_5517)
);

AOI21x1_ASAP7_75t_L g5518 ( 
.A1(n_5207),
.A2(n_5049),
.B(n_4892),
.Y(n_5518)
);

NOR2x1_ASAP7_75t_R g5519 ( 
.A(n_5336),
.B(n_4751),
.Y(n_5519)
);

NAND2x1p5_ASAP7_75t_L g5520 ( 
.A(n_5376),
.B(n_4778),
.Y(n_5520)
);

INVx4_ASAP7_75t_L g5521 ( 
.A(n_5301),
.Y(n_5521)
);

BUFx3_ASAP7_75t_L g5522 ( 
.A(n_5317),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5244),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_5401),
.Y(n_5524)
);

INVx1_ASAP7_75t_L g5525 ( 
.A(n_5373),
.Y(n_5525)
);

BUFx3_ASAP7_75t_L g5526 ( 
.A(n_5248),
.Y(n_5526)
);

BUFx3_ASAP7_75t_L g5527 ( 
.A(n_5209),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5313),
.Y(n_5528)
);

INVx2_ASAP7_75t_L g5529 ( 
.A(n_5406),
.Y(n_5529)
);

INVx2_ASAP7_75t_L g5530 ( 
.A(n_5326),
.Y(n_5530)
);

INVxp67_ASAP7_75t_L g5531 ( 
.A(n_5380),
.Y(n_5531)
);

INVx2_ASAP7_75t_L g5532 ( 
.A(n_5331),
.Y(n_5532)
);

INVx2_ASAP7_75t_L g5533 ( 
.A(n_5124),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_5139),
.Y(n_5534)
);

AOI22xp33_ASAP7_75t_L g5535 ( 
.A1(n_5205),
.A2(n_4930),
.B1(n_5018),
.B2(n_4981),
.Y(n_5535)
);

AND2x2_ASAP7_75t_L g5536 ( 
.A(n_5362),
.B(n_4960),
.Y(n_5536)
);

OAI22xp33_ASAP7_75t_L g5537 ( 
.A1(n_5301),
.A2(n_5239),
.B1(n_5282),
.B2(n_5316),
.Y(n_5537)
);

AND2x2_ASAP7_75t_L g5538 ( 
.A(n_5368),
.B(n_5032),
.Y(n_5538)
);

OAI21x1_ASAP7_75t_L g5539 ( 
.A1(n_5114),
.A2(n_4793),
.B(n_4718),
.Y(n_5539)
);

INVx2_ASAP7_75t_L g5540 ( 
.A(n_5139),
.Y(n_5540)
);

BUFx2_ASAP7_75t_L g5541 ( 
.A(n_5138),
.Y(n_5541)
);

INVx1_ASAP7_75t_L g5542 ( 
.A(n_5275),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_5288),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_5371),
.Y(n_5544)
);

AND2x4_ASAP7_75t_L g5545 ( 
.A(n_5152),
.B(n_4752),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5159),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_5166),
.Y(n_5547)
);

INVx2_ASAP7_75t_L g5548 ( 
.A(n_5166),
.Y(n_5548)
);

AND2x2_ASAP7_75t_L g5549 ( 
.A(n_5252),
.B(n_5052),
.Y(n_5549)
);

INVx2_ASAP7_75t_L g5550 ( 
.A(n_5180),
.Y(n_5550)
);

BUFx2_ASAP7_75t_L g5551 ( 
.A(n_5180),
.Y(n_5551)
);

OAI22xp5_ASAP7_75t_L g5552 ( 
.A1(n_5239),
.A2(n_5090),
.B1(n_4882),
.B2(n_4869),
.Y(n_5552)
);

BUFx3_ASAP7_75t_L g5553 ( 
.A(n_5237),
.Y(n_5553)
);

AOI22xp33_ASAP7_75t_SL g5554 ( 
.A1(n_5228),
.A2(n_4923),
.B1(n_4725),
.B2(n_4836),
.Y(n_5554)
);

INVxp67_ASAP7_75t_L g5555 ( 
.A(n_5336),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5196),
.Y(n_5556)
);

OAI21x1_ASAP7_75t_SL g5557 ( 
.A1(n_5350),
.A2(n_4896),
.B(n_4889),
.Y(n_5557)
);

AND2x2_ASAP7_75t_L g5558 ( 
.A(n_5155),
.B(n_5056),
.Y(n_5558)
);

HB1xp67_ASAP7_75t_L g5559 ( 
.A(n_5135),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5381),
.Y(n_5560)
);

NAND2xp5_ASAP7_75t_L g5561 ( 
.A(n_5100),
.B(n_4878),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_5292),
.Y(n_5562)
);

OAI21x1_ASAP7_75t_L g5563 ( 
.A1(n_5109),
.A2(n_4663),
.B(n_4813),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5292),
.Y(n_5564)
);

INVx2_ASAP7_75t_L g5565 ( 
.A(n_5099),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_5385),
.Y(n_5566)
);

INVx3_ASAP7_75t_L g5567 ( 
.A(n_5241),
.Y(n_5567)
);

HB1xp67_ASAP7_75t_L g5568 ( 
.A(n_5133),
.Y(n_5568)
);

INVx2_ASAP7_75t_L g5569 ( 
.A(n_5315),
.Y(n_5569)
);

OR2x6_ASAP7_75t_L g5570 ( 
.A(n_5355),
.B(n_4645),
.Y(n_5570)
);

INVx2_ASAP7_75t_L g5571 ( 
.A(n_5315),
.Y(n_5571)
);

NAND2xp5_ASAP7_75t_L g5572 ( 
.A(n_5382),
.B(n_5387),
.Y(n_5572)
);

INVx2_ASAP7_75t_L g5573 ( 
.A(n_5404),
.Y(n_5573)
);

OR2x6_ASAP7_75t_L g5574 ( 
.A(n_5282),
.B(n_4652),
.Y(n_5574)
);

OAI21x1_ASAP7_75t_L g5575 ( 
.A1(n_5374),
.A2(n_4901),
.B(n_4898),
.Y(n_5575)
);

CKINVDCx9p33_ASAP7_75t_R g5576 ( 
.A(n_5220),
.Y(n_5576)
);

OA21x2_ASAP7_75t_L g5577 ( 
.A1(n_5121),
.A2(n_4858),
.B(n_4846),
.Y(n_5577)
);

CKINVDCx5p33_ASAP7_75t_R g5578 ( 
.A(n_5117),
.Y(n_5578)
);

NAND2xp5_ASAP7_75t_L g5579 ( 
.A(n_5227),
.B(n_4989),
.Y(n_5579)
);

OR2x2_ASAP7_75t_L g5580 ( 
.A(n_5544),
.B(n_5129),
.Y(n_5580)
);

AND2x2_ASAP7_75t_L g5581 ( 
.A(n_5421),
.B(n_4947),
.Y(n_5581)
);

NOR2x1_ASAP7_75t_R g5582 ( 
.A(n_5478),
.B(n_4774),
.Y(n_5582)
);

NAND2xp5_ASAP7_75t_L g5583 ( 
.A(n_5546),
.B(n_5398),
.Y(n_5583)
);

NOR2xp33_ASAP7_75t_R g5584 ( 
.A(n_5490),
.B(n_5322),
.Y(n_5584)
);

NAND2xp33_ASAP7_75t_L g5585 ( 
.A(n_5433),
.B(n_5267),
.Y(n_5585)
);

AND2x2_ASAP7_75t_L g5586 ( 
.A(n_5487),
.B(n_5393),
.Y(n_5586)
);

HB1xp67_ASAP7_75t_L g5587 ( 
.A(n_5568),
.Y(n_5587)
);

OAI22xp5_ASAP7_75t_L g5588 ( 
.A1(n_5574),
.A2(n_5316),
.B1(n_4833),
.B2(n_5410),
.Y(n_5588)
);

INVx8_ASAP7_75t_L g5589 ( 
.A(n_5570),
.Y(n_5589)
);

AND2x2_ASAP7_75t_L g5590 ( 
.A(n_5488),
.B(n_5256),
.Y(n_5590)
);

NOR2xp33_ASAP7_75t_R g5591 ( 
.A(n_5578),
.B(n_5337),
.Y(n_5591)
);

INVx2_ASAP7_75t_L g5592 ( 
.A(n_5431),
.Y(n_5592)
);

CKINVDCx16_ASAP7_75t_R g5593 ( 
.A(n_5522),
.Y(n_5593)
);

OR2x2_ASAP7_75t_L g5594 ( 
.A(n_5417),
.B(n_5130),
.Y(n_5594)
);

AND2x2_ASAP7_75t_L g5595 ( 
.A(n_5448),
.B(n_5258),
.Y(n_5595)
);

AOI22xp33_ASAP7_75t_SL g5596 ( 
.A1(n_5521),
.A2(n_5435),
.B1(n_5552),
.B2(n_5574),
.Y(n_5596)
);

HB1xp67_ASAP7_75t_L g5597 ( 
.A(n_5431),
.Y(n_5597)
);

NAND2xp5_ASAP7_75t_L g5598 ( 
.A(n_5528),
.B(n_5482),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5415),
.Y(n_5599)
);

OAI22xp5_ASAP7_75t_L g5600 ( 
.A1(n_5509),
.A2(n_5131),
.B1(n_4953),
.B2(n_5319),
.Y(n_5600)
);

AND2x2_ASAP7_75t_L g5601 ( 
.A(n_5493),
.B(n_5258),
.Y(n_5601)
);

NAND2xp33_ASAP7_75t_R g5602 ( 
.A(n_5570),
.B(n_5397),
.Y(n_5602)
);

AND2x2_ASAP7_75t_L g5603 ( 
.A(n_5559),
.B(n_5324),
.Y(n_5603)
);

OAI22xp5_ASAP7_75t_L g5604 ( 
.A1(n_5467),
.A2(n_5235),
.B1(n_5225),
.B2(n_5164),
.Y(n_5604)
);

INVxp67_ASAP7_75t_L g5605 ( 
.A(n_5441),
.Y(n_5605)
);

NAND2xp5_ASAP7_75t_L g5606 ( 
.A(n_5542),
.B(n_5375),
.Y(n_5606)
);

HB1xp67_ASAP7_75t_L g5607 ( 
.A(n_5457),
.Y(n_5607)
);

HB1xp67_ASAP7_75t_L g5608 ( 
.A(n_5457),
.Y(n_5608)
);

INVx3_ASAP7_75t_L g5609 ( 
.A(n_5476),
.Y(n_5609)
);

AND2x2_ASAP7_75t_L g5610 ( 
.A(n_5565),
.B(n_4933),
.Y(n_5610)
);

AND2x4_ASAP7_75t_L g5611 ( 
.A(n_5481),
.B(n_5392),
.Y(n_5611)
);

AOI22xp33_ASAP7_75t_SL g5612 ( 
.A1(n_5435),
.A2(n_5178),
.B1(n_5328),
.B2(n_5183),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5416),
.Y(n_5613)
);

AOI22xp33_ASAP7_75t_L g5614 ( 
.A1(n_5506),
.A2(n_5096),
.B1(n_5079),
.B2(n_4997),
.Y(n_5614)
);

NAND2xp5_ASAP7_75t_L g5615 ( 
.A(n_5543),
.B(n_5283),
.Y(n_5615)
);

AND2x2_ASAP7_75t_L g5616 ( 
.A(n_5558),
.B(n_5104),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5418),
.Y(n_5617)
);

INVx3_ASAP7_75t_L g5618 ( 
.A(n_5441),
.Y(n_5618)
);

OR2x2_ASAP7_75t_L g5619 ( 
.A(n_5426),
.B(n_5217),
.Y(n_5619)
);

INVx2_ASAP7_75t_L g5620 ( 
.A(n_5428),
.Y(n_5620)
);

HB1xp67_ASAP7_75t_L g5621 ( 
.A(n_5459),
.Y(n_5621)
);

BUFx3_ASAP7_75t_L g5622 ( 
.A(n_5511),
.Y(n_5622)
);

AOI22xp5_ASAP7_75t_L g5623 ( 
.A1(n_5442),
.A2(n_5274),
.B1(n_5108),
.B2(n_5372),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5422),
.Y(n_5624)
);

OR2x2_ASAP7_75t_L g5625 ( 
.A(n_5530),
.B(n_5188),
.Y(n_5625)
);

NAND3xp33_ASAP7_75t_SL g5626 ( 
.A(n_5554),
.B(n_5365),
.C(n_5320),
.Y(n_5626)
);

NAND2xp5_ASAP7_75t_L g5627 ( 
.A(n_5556),
.B(n_5302),
.Y(n_5627)
);

NAND2xp33_ASAP7_75t_R g5628 ( 
.A(n_5567),
.B(n_5404),
.Y(n_5628)
);

NOR2xp33_ASAP7_75t_L g5629 ( 
.A(n_5519),
.B(n_5218),
.Y(n_5629)
);

HB1xp67_ASAP7_75t_L g5630 ( 
.A(n_5531),
.Y(n_5630)
);

HB1xp67_ASAP7_75t_L g5631 ( 
.A(n_5464),
.Y(n_5631)
);

AO21x2_ASAP7_75t_L g5632 ( 
.A1(n_5533),
.A2(n_5477),
.B(n_5537),
.Y(n_5632)
);

NAND2xp5_ASAP7_75t_L g5633 ( 
.A(n_5560),
.B(n_5195),
.Y(n_5633)
);

AOI22xp33_ASAP7_75t_L g5634 ( 
.A1(n_5474),
.A2(n_5001),
.B1(n_4964),
.B2(n_5200),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5425),
.Y(n_5635)
);

AND2x2_ASAP7_75t_L g5636 ( 
.A(n_5538),
.B(n_5403),
.Y(n_5636)
);

BUFx3_ASAP7_75t_L g5637 ( 
.A(n_5553),
.Y(n_5637)
);

NAND2xp5_ASAP7_75t_L g5638 ( 
.A(n_5532),
.B(n_5162),
.Y(n_5638)
);

AND2x4_ASAP7_75t_L g5639 ( 
.A(n_5481),
.B(n_5212),
.Y(n_5639)
);

INVxp67_ASAP7_75t_L g5640 ( 
.A(n_5517),
.Y(n_5640)
);

INVx1_ASAP7_75t_SL g5641 ( 
.A(n_5483),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_5484),
.B(n_5162),
.Y(n_5642)
);

HB1xp67_ASAP7_75t_L g5643 ( 
.A(n_5473),
.Y(n_5643)
);

BUFx2_ASAP7_75t_L g5644 ( 
.A(n_5508),
.Y(n_5644)
);

AOI22xp33_ASAP7_75t_L g5645 ( 
.A1(n_5496),
.A2(n_5192),
.B1(n_5154),
.B2(n_4867),
.Y(n_5645)
);

NOR3xp33_ASAP7_75t_SL g5646 ( 
.A(n_5430),
.B(n_5389),
.C(n_4796),
.Y(n_5646)
);

NAND2xp33_ASAP7_75t_R g5647 ( 
.A(n_5438),
.B(n_5391),
.Y(n_5647)
);

BUFx3_ASAP7_75t_L g5648 ( 
.A(n_5527),
.Y(n_5648)
);

AO31x2_ASAP7_75t_L g5649 ( 
.A1(n_5562),
.A2(n_5213),
.A3(n_5203),
.B(n_5304),
.Y(n_5649)
);

CKINVDCx5p33_ASAP7_75t_R g5650 ( 
.A(n_5480),
.Y(n_5650)
);

INVx2_ASAP7_75t_L g5651 ( 
.A(n_5432),
.Y(n_5651)
);

NOR2xp33_ASAP7_75t_R g5652 ( 
.A(n_5440),
.B(n_4741),
.Y(n_5652)
);

OR2x2_ASAP7_75t_L g5653 ( 
.A(n_5502),
.B(n_5469),
.Y(n_5653)
);

NAND3xp33_ASAP7_75t_L g5654 ( 
.A(n_5535),
.B(n_5408),
.C(n_5335),
.Y(n_5654)
);

NOR2xp33_ASAP7_75t_R g5655 ( 
.A(n_5429),
.B(n_4748),
.Y(n_5655)
);

NAND2xp33_ASAP7_75t_R g5656 ( 
.A(n_5485),
.B(n_5391),
.Y(n_5656)
);

AOI21xp33_ASAP7_75t_L g5657 ( 
.A1(n_5472),
.A2(n_5411),
.B(n_5136),
.Y(n_5657)
);

NAND2xp5_ASAP7_75t_L g5658 ( 
.A(n_5486),
.B(n_5025),
.Y(n_5658)
);

INVx2_ASAP7_75t_L g5659 ( 
.A(n_5446),
.Y(n_5659)
);

INVx1_ASAP7_75t_L g5660 ( 
.A(n_5427),
.Y(n_5660)
);

INVx1_ASAP7_75t_L g5661 ( 
.A(n_5434),
.Y(n_5661)
);

CKINVDCx16_ASAP7_75t_R g5662 ( 
.A(n_5491),
.Y(n_5662)
);

INVx1_ASAP7_75t_L g5663 ( 
.A(n_5443),
.Y(n_5663)
);

AOI21xp33_ASAP7_75t_L g5664 ( 
.A1(n_5557),
.A2(n_5281),
.B(n_5363),
.Y(n_5664)
);

NAND3xp33_ASAP7_75t_SL g5665 ( 
.A(n_5513),
.B(n_5273),
.C(n_5342),
.Y(n_5665)
);

INVx1_ASAP7_75t_SL g5666 ( 
.A(n_5526),
.Y(n_5666)
);

AOI211xp5_ASAP7_75t_L g5667 ( 
.A1(n_5466),
.A2(n_5255),
.B(n_5318),
.C(n_5161),
.Y(n_5667)
);

NOR2xp33_ASAP7_75t_R g5668 ( 
.A(n_5515),
.B(n_5232),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5454),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_5455),
.Y(n_5670)
);

AND2x2_ASAP7_75t_L g5671 ( 
.A(n_5549),
.B(n_5403),
.Y(n_5671)
);

OAI22xp5_ASAP7_75t_L g5672 ( 
.A1(n_5424),
.A2(n_4986),
.B1(n_5132),
.B2(n_5167),
.Y(n_5672)
);

AOI22xp33_ASAP7_75t_L g5673 ( 
.A1(n_5566),
.A2(n_5017),
.B1(n_5044),
.B2(n_5012),
.Y(n_5673)
);

NOR3xp33_ASAP7_75t_SL g5674 ( 
.A(n_5579),
.B(n_4795),
.C(n_4794),
.Y(n_5674)
);

NOR2xp33_ASAP7_75t_R g5675 ( 
.A(n_5501),
.B(n_4871),
.Y(n_5675)
);

NAND2xp33_ASAP7_75t_R g5676 ( 
.A(n_5504),
.B(n_5323),
.Y(n_5676)
);

AND2x2_ASAP7_75t_L g5677 ( 
.A(n_5439),
.B(n_4899),
.Y(n_5677)
);

NOR2xp33_ASAP7_75t_R g5678 ( 
.A(n_5419),
.B(n_5329),
.Y(n_5678)
);

NAND3xp33_ASAP7_75t_L g5679 ( 
.A(n_5577),
.B(n_5190),
.C(n_5354),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5456),
.Y(n_5680)
);

OAI21xp5_ASAP7_75t_SL g5681 ( 
.A1(n_5489),
.A2(n_5158),
.B(n_5284),
.Y(n_5681)
);

HB1xp67_ASAP7_75t_L g5682 ( 
.A(n_5475),
.Y(n_5682)
);

INVx2_ASAP7_75t_L g5683 ( 
.A(n_5453),
.Y(n_5683)
);

OR2x2_ASAP7_75t_L g5684 ( 
.A(n_5492),
.B(n_5330),
.Y(n_5684)
);

AND2x2_ASAP7_75t_L g5685 ( 
.A(n_5514),
.B(n_4899),
.Y(n_5685)
);

BUFx6f_ASAP7_75t_L g5686 ( 
.A(n_5419),
.Y(n_5686)
);

NAND2xp5_ASAP7_75t_L g5687 ( 
.A(n_5414),
.B(n_5045),
.Y(n_5687)
);

HB1xp67_ASAP7_75t_L g5688 ( 
.A(n_5495),
.Y(n_5688)
);

O2A1O1Ixp33_ASAP7_75t_SL g5689 ( 
.A1(n_5555),
.A2(n_5120),
.B(n_5182),
.C(n_5333),
.Y(n_5689)
);

OAI222xp33_ASAP7_75t_L g5690 ( 
.A1(n_5445),
.A2(n_5127),
.B1(n_5378),
.B2(n_5249),
.C1(n_5360),
.C2(n_5339),
.Y(n_5690)
);

NOR3xp33_ASAP7_75t_SL g5691 ( 
.A(n_5561),
.B(n_4851),
.C(n_5144),
.Y(n_5691)
);

INVx2_ASAP7_75t_L g5692 ( 
.A(n_5458),
.Y(n_5692)
);

AND2x2_ASAP7_75t_L g5693 ( 
.A(n_5536),
.B(n_4899),
.Y(n_5693)
);

INVx2_ASAP7_75t_L g5694 ( 
.A(n_5462),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_L g5695 ( 
.A(n_5497),
.B(n_5059),
.Y(n_5695)
);

OR2x2_ASAP7_75t_SL g5696 ( 
.A(n_5437),
.B(n_5323),
.Y(n_5696)
);

INVx2_ASAP7_75t_L g5697 ( 
.A(n_5465),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5461),
.Y(n_5698)
);

BUFx4_ASAP7_75t_SL g5699 ( 
.A(n_5471),
.Y(n_5699)
);

NAND2xp33_ASAP7_75t_R g5700 ( 
.A(n_5505),
.B(n_5219),
.Y(n_5700)
);

AND2x2_ASAP7_75t_L g5701 ( 
.A(n_5494),
.B(n_4944),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5463),
.Y(n_5702)
);

INVx1_ASAP7_75t_L g5703 ( 
.A(n_5631),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5643),
.Y(n_5704)
);

HB1xp67_ASAP7_75t_L g5705 ( 
.A(n_5688),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5682),
.Y(n_5706)
);

AOI221xp5_ASAP7_75t_L g5707 ( 
.A1(n_5689),
.A2(n_5525),
.B1(n_5523),
.B2(n_5572),
.C(n_5436),
.Y(n_5707)
);

AND2x4_ASAP7_75t_L g5708 ( 
.A(n_5632),
.B(n_5471),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_5615),
.B(n_5564),
.Y(n_5709)
);

OR2x2_ASAP7_75t_L g5710 ( 
.A(n_5625),
.B(n_5423),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5598),
.Y(n_5711)
);

BUFx2_ASAP7_75t_SL g5712 ( 
.A(n_5611),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5599),
.Y(n_5713)
);

OR2x2_ASAP7_75t_SL g5714 ( 
.A(n_5662),
.B(n_5437),
.Y(n_5714)
);

AND2x4_ASAP7_75t_L g5715 ( 
.A(n_5616),
.B(n_5541),
.Y(n_5715)
);

AND2x2_ASAP7_75t_L g5716 ( 
.A(n_5590),
.B(n_5541),
.Y(n_5716)
);

INVx2_ASAP7_75t_L g5717 ( 
.A(n_5597),
.Y(n_5717)
);

INVx2_ASAP7_75t_L g5718 ( 
.A(n_5607),
.Y(n_5718)
);

NAND2xp33_ASAP7_75t_L g5719 ( 
.A(n_5589),
.B(n_5419),
.Y(n_5719)
);

BUFx2_ASAP7_75t_L g5720 ( 
.A(n_5648),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5613),
.Y(n_5721)
);

INVx2_ASAP7_75t_L g5722 ( 
.A(n_5608),
.Y(n_5722)
);

INVx3_ASAP7_75t_L g5723 ( 
.A(n_5589),
.Y(n_5723)
);

AND2x2_ASAP7_75t_L g5724 ( 
.A(n_5671),
.B(n_5551),
.Y(n_5724)
);

NAND2xp5_ASAP7_75t_L g5725 ( 
.A(n_5627),
.B(n_5444),
.Y(n_5725)
);

INVx2_ASAP7_75t_L g5726 ( 
.A(n_5620),
.Y(n_5726)
);

AND2x2_ASAP7_75t_L g5727 ( 
.A(n_5636),
.B(n_5551),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_5617),
.Y(n_5728)
);

INVx2_ASAP7_75t_SL g5729 ( 
.A(n_5699),
.Y(n_5729)
);

AND2x4_ASAP7_75t_SL g5730 ( 
.A(n_5639),
.B(n_5470),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5624),
.Y(n_5731)
);

INVx2_ASAP7_75t_L g5732 ( 
.A(n_5651),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_5635),
.Y(n_5733)
);

AND2x2_ASAP7_75t_L g5734 ( 
.A(n_5586),
.B(n_5512),
.Y(n_5734)
);

AOI22xp5_ASAP7_75t_L g5735 ( 
.A1(n_5672),
.A2(n_5460),
.B1(n_5073),
.B2(n_5061),
.Y(n_5735)
);

AND2x2_ASAP7_75t_L g5736 ( 
.A(n_5587),
.B(n_5547),
.Y(n_5736)
);

OR2x2_ASAP7_75t_L g5737 ( 
.A(n_5653),
.B(n_5447),
.Y(n_5737)
);

AND2x2_ASAP7_75t_L g5738 ( 
.A(n_5644),
.B(n_5548),
.Y(n_5738)
);

OR2x2_ASAP7_75t_L g5739 ( 
.A(n_5594),
.B(n_5449),
.Y(n_5739)
);

INVx1_ASAP7_75t_L g5740 ( 
.A(n_5660),
.Y(n_5740)
);

INVx2_ASAP7_75t_L g5741 ( 
.A(n_5659),
.Y(n_5741)
);

INVx2_ASAP7_75t_L g5742 ( 
.A(n_5683),
.Y(n_5742)
);

HB1xp67_ASAP7_75t_L g5743 ( 
.A(n_5621),
.Y(n_5743)
);

NAND2x1p5_ASAP7_75t_L g5744 ( 
.A(n_5622),
.B(n_5507),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_5661),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5663),
.Y(n_5746)
);

INVxp67_ASAP7_75t_SL g5747 ( 
.A(n_5628),
.Y(n_5747)
);

AND2x4_ASAP7_75t_L g5748 ( 
.A(n_5610),
.B(n_5550),
.Y(n_5748)
);

BUFx2_ASAP7_75t_L g5749 ( 
.A(n_5637),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_5669),
.Y(n_5750)
);

INVx1_ASAP7_75t_L g5751 ( 
.A(n_5670),
.Y(n_5751)
);

AOI22xp33_ASAP7_75t_SL g5752 ( 
.A1(n_5600),
.A2(n_5557),
.B1(n_5577),
.B2(n_5545),
.Y(n_5752)
);

AND2x4_ASAP7_75t_L g5753 ( 
.A(n_5685),
.B(n_5573),
.Y(n_5753)
);

AND2x2_ASAP7_75t_L g5754 ( 
.A(n_5630),
.B(n_5468),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_5680),
.Y(n_5755)
);

AND2x2_ASAP7_75t_L g5756 ( 
.A(n_5603),
.B(n_5581),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5698),
.Y(n_5757)
);

BUFx3_ASAP7_75t_L g5758 ( 
.A(n_5666),
.Y(n_5758)
);

NAND2xp5_ASAP7_75t_L g5759 ( 
.A(n_5583),
.B(n_5498),
.Y(n_5759)
);

NAND2xp5_ASAP7_75t_L g5760 ( 
.A(n_5642),
.B(n_5638),
.Y(n_5760)
);

AND2x2_ASAP7_75t_L g5761 ( 
.A(n_5677),
.B(n_5503),
.Y(n_5761)
);

AND2x2_ASAP7_75t_L g5762 ( 
.A(n_5693),
.B(n_5592),
.Y(n_5762)
);

OAI222xp33_ASAP7_75t_L g5763 ( 
.A1(n_5596),
.A2(n_5500),
.B1(n_5518),
.B2(n_5520),
.C1(n_5420),
.C2(n_5450),
.Y(n_5763)
);

HB1xp67_ASAP7_75t_L g5764 ( 
.A(n_5692),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5702),
.Y(n_5765)
);

INVx2_ASAP7_75t_L g5766 ( 
.A(n_5694),
.Y(n_5766)
);

AND2x2_ASAP7_75t_L g5767 ( 
.A(n_5701),
.B(n_5510),
.Y(n_5767)
);

AND2x2_ASAP7_75t_L g5768 ( 
.A(n_5640),
.B(n_5516),
.Y(n_5768)
);

AND2x4_ASAP7_75t_L g5769 ( 
.A(n_5639),
.B(n_5569),
.Y(n_5769)
);

NAND2xp5_ASAP7_75t_L g5770 ( 
.A(n_5633),
.B(n_5499),
.Y(n_5770)
);

AND2x2_ASAP7_75t_L g5771 ( 
.A(n_5595),
.B(n_5524),
.Y(n_5771)
);

INVx2_ASAP7_75t_L g5772 ( 
.A(n_5697),
.Y(n_5772)
);

HB1xp67_ASAP7_75t_L g5773 ( 
.A(n_5619),
.Y(n_5773)
);

INVx2_ASAP7_75t_L g5774 ( 
.A(n_5696),
.Y(n_5774)
);

AND2x2_ASAP7_75t_L g5775 ( 
.A(n_5605),
.B(n_5529),
.Y(n_5775)
);

NAND2xp5_ASAP7_75t_L g5776 ( 
.A(n_5684),
.B(n_5451),
.Y(n_5776)
);

AO31x2_ASAP7_75t_L g5777 ( 
.A1(n_5629),
.A2(n_5534),
.A3(n_5540),
.B(n_5571),
.Y(n_5777)
);

AND2x2_ASAP7_75t_L g5778 ( 
.A(n_5601),
.B(n_5452),
.Y(n_5778)
);

OR2x2_ASAP7_75t_L g5779 ( 
.A(n_5580),
.B(n_5479),
.Y(n_5779)
);

INVx2_ASAP7_75t_L g5780 ( 
.A(n_5609),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_5695),
.Y(n_5781)
);

INVxp67_ASAP7_75t_SL g5782 ( 
.A(n_5656),
.Y(n_5782)
);

NAND2xp5_ASAP7_75t_L g5783 ( 
.A(n_5606),
.B(n_5563),
.Y(n_5783)
);

AOI22xp5_ASAP7_75t_L g5784 ( 
.A1(n_5665),
.A2(n_5063),
.B1(n_5066),
.B2(n_5021),
.Y(n_5784)
);

INVx3_ASAP7_75t_L g5785 ( 
.A(n_5686),
.Y(n_5785)
);

INVx3_ASAP7_75t_L g5786 ( 
.A(n_5686),
.Y(n_5786)
);

INVx5_ASAP7_75t_L g5787 ( 
.A(n_5686),
.Y(n_5787)
);

INVx2_ASAP7_75t_L g5788 ( 
.A(n_5658),
.Y(n_5788)
);

AOI221xp5_ASAP7_75t_L g5789 ( 
.A1(n_5679),
.A2(n_5264),
.B1(n_5266),
.B2(n_4984),
.C(n_5377),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_5687),
.Y(n_5790)
);

AND2x2_ASAP7_75t_L g5791 ( 
.A(n_5618),
.B(n_5575),
.Y(n_5791)
);

INVx3_ASAP7_75t_L g5792 ( 
.A(n_5593),
.Y(n_5792)
);

NAND2x1p5_ASAP7_75t_L g5793 ( 
.A(n_5641),
.B(n_4778),
.Y(n_5793)
);

INVx2_ASAP7_75t_SL g5794 ( 
.A(n_5675),
.Y(n_5794)
);

HB1xp67_ASAP7_75t_L g5795 ( 
.A(n_5602),
.Y(n_5795)
);

AO21x2_ASAP7_75t_L g5796 ( 
.A1(n_5678),
.A2(n_5591),
.B(n_5584),
.Y(n_5796)
);

INVx1_ASAP7_75t_L g5797 ( 
.A(n_5649),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5649),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5649),
.Y(n_5799)
);

INVx2_ASAP7_75t_SL g5800 ( 
.A(n_5668),
.Y(n_5800)
);

INVx1_ASAP7_75t_L g5801 ( 
.A(n_5673),
.Y(n_5801)
);

INVx1_ASAP7_75t_SL g5802 ( 
.A(n_5720),
.Y(n_5802)
);

AND2x2_ASAP7_75t_L g5803 ( 
.A(n_5795),
.B(n_5612),
.Y(n_5803)
);

INVxp67_ASAP7_75t_SL g5804 ( 
.A(n_5705),
.Y(n_5804)
);

INVx2_ASAP7_75t_L g5805 ( 
.A(n_5720),
.Y(n_5805)
);

OAI21x1_ASAP7_75t_L g5806 ( 
.A1(n_5744),
.A2(n_5614),
.B(n_5588),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5743),
.Y(n_5807)
);

NAND3xp33_ASAP7_75t_L g5808 ( 
.A(n_5752),
.B(n_5634),
.C(n_5645),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5773),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5764),
.Y(n_5810)
);

INVx2_ASAP7_75t_L g5811 ( 
.A(n_5749),
.Y(n_5811)
);

INVx2_ASAP7_75t_L g5812 ( 
.A(n_5749),
.Y(n_5812)
);

BUFx3_ASAP7_75t_L g5813 ( 
.A(n_5758),
.Y(n_5813)
);

OAI221xp5_ASAP7_75t_L g5814 ( 
.A1(n_5735),
.A2(n_5667),
.B1(n_5681),
.B2(n_5700),
.C(n_5691),
.Y(n_5814)
);

OAI21x1_ASAP7_75t_L g5815 ( 
.A1(n_5782),
.A2(n_5604),
.B(n_5690),
.Y(n_5815)
);

AOI22xp33_ASAP7_75t_L g5816 ( 
.A1(n_5796),
.A2(n_5626),
.B1(n_5657),
.B2(n_5664),
.Y(n_5816)
);

INVx2_ASAP7_75t_L g5817 ( 
.A(n_5717),
.Y(n_5817)
);

INVx2_ASAP7_75t_L g5818 ( 
.A(n_5718),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5722),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_5703),
.Y(n_5820)
);

NAND2xp5_ASAP7_75t_L g5821 ( 
.A(n_5704),
.B(n_5539),
.Y(n_5821)
);

OAI22xp5_ASAP7_75t_L g5822 ( 
.A1(n_5712),
.A2(n_5674),
.B1(n_5646),
.B2(n_5623),
.Y(n_5822)
);

AOI21xp5_ASAP7_75t_L g5823 ( 
.A1(n_5719),
.A2(n_5585),
.B(n_5582),
.Y(n_5823)
);

AOI22xp33_ASAP7_75t_L g5824 ( 
.A1(n_5801),
.A2(n_5654),
.B1(n_5176),
.B2(n_5017),
.Y(n_5824)
);

AND2x2_ASAP7_75t_L g5825 ( 
.A(n_5715),
.B(n_5655),
.Y(n_5825)
);

OR2x2_ASAP7_75t_L g5826 ( 
.A(n_5725),
.B(n_5105),
.Y(n_5826)
);

OAI211xp5_ASAP7_75t_SL g5827 ( 
.A1(n_5707),
.A2(n_5341),
.B(n_5271),
.C(n_4959),
.Y(n_5827)
);

AOI22xp5_ASAP7_75t_L g5828 ( 
.A1(n_5747),
.A2(n_5647),
.B1(n_5676),
.B2(n_5312),
.Y(n_5828)
);

AO21x2_ASAP7_75t_L g5829 ( 
.A1(n_5763),
.A2(n_5774),
.B(n_5797),
.Y(n_5829)
);

INVxp67_ASAP7_75t_L g5830 ( 
.A(n_5712),
.Y(n_5830)
);

AOI21xp5_ASAP7_75t_SL g5831 ( 
.A1(n_5729),
.A2(n_5576),
.B(n_5650),
.Y(n_5831)
);

AND2x4_ASAP7_75t_L g5832 ( 
.A(n_5730),
.B(n_5004),
.Y(n_5832)
);

AOI21xp5_ASAP7_75t_L g5833 ( 
.A1(n_5794),
.A2(n_5268),
.B(n_5286),
.Y(n_5833)
);

INVxp67_ASAP7_75t_L g5834 ( 
.A(n_5792),
.Y(n_5834)
);

INVx2_ASAP7_75t_L g5835 ( 
.A(n_5726),
.Y(n_5835)
);

OAI21xp33_ASAP7_75t_L g5836 ( 
.A1(n_5798),
.A2(n_5652),
.B(n_4979),
.Y(n_5836)
);

AND2x2_ASAP7_75t_L g5837 ( 
.A(n_5715),
.B(n_4976),
.Y(n_5837)
);

BUFx2_ASAP7_75t_L g5838 ( 
.A(n_5793),
.Y(n_5838)
);

NAND2xp5_ASAP7_75t_L g5839 ( 
.A(n_5706),
.B(n_5119),
.Y(n_5839)
);

NAND2xp5_ASAP7_75t_L g5840 ( 
.A(n_5783),
.B(n_5119),
.Y(n_5840)
);

INVx2_ASAP7_75t_L g5841 ( 
.A(n_5732),
.Y(n_5841)
);

OR2x6_ASAP7_75t_L g5842 ( 
.A(n_5800),
.B(n_4656),
.Y(n_5842)
);

INVx2_ASAP7_75t_L g5843 ( 
.A(n_5741),
.Y(n_5843)
);

INVx2_ASAP7_75t_L g5844 ( 
.A(n_5742),
.Y(n_5844)
);

NAND2xp5_ASAP7_75t_L g5845 ( 
.A(n_5760),
.B(n_5260),
.Y(n_5845)
);

HB1xp67_ASAP7_75t_L g5846 ( 
.A(n_5759),
.Y(n_5846)
);

INVx4_ASAP7_75t_SL g5847 ( 
.A(n_5777),
.Y(n_5847)
);

INVx1_ASAP7_75t_L g5848 ( 
.A(n_5713),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5737),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_5766),
.Y(n_5850)
);

INVx1_ASAP7_75t_L g5851 ( 
.A(n_5721),
.Y(n_5851)
);

INVx1_ASAP7_75t_L g5852 ( 
.A(n_5728),
.Y(n_5852)
);

OA21x2_ASAP7_75t_L g5853 ( 
.A1(n_5708),
.A2(n_5126),
.B(n_5165),
.Y(n_5853)
);

AND2x4_ASAP7_75t_L g5854 ( 
.A(n_5791),
.B(n_5332),
.Y(n_5854)
);

AOI22xp5_ASAP7_75t_L g5855 ( 
.A1(n_5784),
.A2(n_5065),
.B1(n_5067),
.B2(n_5064),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5731),
.Y(n_5856)
);

BUFx2_ASAP7_75t_L g5857 ( 
.A(n_5723),
.Y(n_5857)
);

HB1xp67_ASAP7_75t_L g5858 ( 
.A(n_5777),
.Y(n_5858)
);

OAI22xp5_ASAP7_75t_L g5859 ( 
.A1(n_5714),
.A2(n_4944),
.B1(n_5033),
.B2(n_4781),
.Y(n_5859)
);

OR2x2_ASAP7_75t_L g5860 ( 
.A(n_5709),
.B(n_5394),
.Y(n_5860)
);

AND2x2_ASAP7_75t_L g5861 ( 
.A(n_5724),
.B(n_4978),
.Y(n_5861)
);

INVx2_ASAP7_75t_L g5862 ( 
.A(n_5772),
.Y(n_5862)
);

AND2x2_ASAP7_75t_L g5863 ( 
.A(n_5727),
.B(n_4781),
.Y(n_5863)
);

NOR2xp33_ASAP7_75t_L g5864 ( 
.A(n_5711),
.B(n_5390),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5733),
.Y(n_5865)
);

BUFx2_ASAP7_75t_L g5866 ( 
.A(n_5787),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5740),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5745),
.Y(n_5868)
);

INVx2_ASAP7_75t_L g5869 ( 
.A(n_5746),
.Y(n_5869)
);

AND2x2_ASAP7_75t_L g5870 ( 
.A(n_5716),
.B(n_5137),
.Y(n_5870)
);

INVx2_ASAP7_75t_L g5871 ( 
.A(n_5750),
.Y(n_5871)
);

AOI22xp5_ASAP7_75t_SL g5872 ( 
.A1(n_5734),
.A2(n_5708),
.B1(n_5769),
.B2(n_5754),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5751),
.Y(n_5873)
);

OA21x2_ASAP7_75t_L g5874 ( 
.A1(n_5799),
.A2(n_5293),
.B(n_5202),
.Y(n_5874)
);

NAND2xp5_ASAP7_75t_L g5875 ( 
.A(n_5781),
.B(n_5394),
.Y(n_5875)
);

INVx2_ASAP7_75t_L g5876 ( 
.A(n_5805),
.Y(n_5876)
);

INVx2_ASAP7_75t_L g5877 ( 
.A(n_5811),
.Y(n_5877)
);

AND2x2_ASAP7_75t_L g5878 ( 
.A(n_5838),
.B(n_5769),
.Y(n_5878)
);

OAI33xp33_ASAP7_75t_L g5879 ( 
.A1(n_5822),
.A2(n_5790),
.A3(n_5770),
.B1(n_5757),
.B2(n_5755),
.B3(n_5765),
.Y(n_5879)
);

OAI33xp33_ASAP7_75t_L g5880 ( 
.A1(n_5808),
.A2(n_5776),
.A3(n_5779),
.B1(n_5788),
.B2(n_5710),
.B3(n_5780),
.Y(n_5880)
);

NOR2x1_ASAP7_75t_L g5881 ( 
.A(n_5842),
.B(n_5308),
.Y(n_5881)
);

INVx1_ASAP7_75t_SL g5882 ( 
.A(n_5813),
.Y(n_5882)
);

INVxp67_ASAP7_75t_L g5883 ( 
.A(n_5857),
.Y(n_5883)
);

AND2x2_ASAP7_75t_L g5884 ( 
.A(n_5872),
.B(n_5738),
.Y(n_5884)
);

AND2x4_ASAP7_75t_L g5885 ( 
.A(n_5842),
.B(n_5830),
.Y(n_5885)
);

INVx2_ASAP7_75t_L g5886 ( 
.A(n_5812),
.Y(n_5886)
);

OAI21xp33_ASAP7_75t_L g5887 ( 
.A1(n_5816),
.A2(n_5736),
.B(n_5768),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5804),
.Y(n_5888)
);

INVx1_ASAP7_75t_L g5889 ( 
.A(n_5809),
.Y(n_5889)
);

INVx5_ASAP7_75t_L g5890 ( 
.A(n_5866),
.Y(n_5890)
);

NOR2xp33_ASAP7_75t_R g5891 ( 
.A(n_5834),
.B(n_5787),
.Y(n_5891)
);

HB1xp67_ASAP7_75t_L g5892 ( 
.A(n_5802),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5807),
.Y(n_5893)
);

INVx2_ASAP7_75t_L g5894 ( 
.A(n_5810),
.Y(n_5894)
);

HB1xp67_ASAP7_75t_L g5895 ( 
.A(n_5869),
.Y(n_5895)
);

BUFx2_ASAP7_75t_L g5896 ( 
.A(n_5806),
.Y(n_5896)
);

AND2x2_ASAP7_75t_L g5897 ( 
.A(n_5803),
.B(n_5748),
.Y(n_5897)
);

AOI22xp5_ASAP7_75t_L g5898 ( 
.A1(n_5814),
.A2(n_5789),
.B1(n_5748),
.B2(n_5775),
.Y(n_5898)
);

INVx2_ASAP7_75t_L g5899 ( 
.A(n_5835),
.Y(n_5899)
);

BUFx2_ASAP7_75t_L g5900 ( 
.A(n_5847),
.Y(n_5900)
);

AND2x2_ASAP7_75t_L g5901 ( 
.A(n_5825),
.B(n_5756),
.Y(n_5901)
);

OR2x2_ASAP7_75t_L g5902 ( 
.A(n_5845),
.B(n_5739),
.Y(n_5902)
);

BUFx2_ASAP7_75t_L g5903 ( 
.A(n_5847),
.Y(n_5903)
);

AND2x4_ASAP7_75t_SL g5904 ( 
.A(n_5832),
.B(n_5771),
.Y(n_5904)
);

OAI31xp33_ASAP7_75t_SL g5905 ( 
.A1(n_5815),
.A2(n_5778),
.A3(n_5753),
.B(n_5767),
.Y(n_5905)
);

AND2x2_ASAP7_75t_L g5906 ( 
.A(n_5846),
.B(n_5761),
.Y(n_5906)
);

AND2x2_ASAP7_75t_L g5907 ( 
.A(n_5870),
.B(n_5762),
.Y(n_5907)
);

INVx4_ASAP7_75t_L g5908 ( 
.A(n_5832),
.Y(n_5908)
);

OAI221xp5_ASAP7_75t_L g5909 ( 
.A1(n_5828),
.A2(n_5785),
.B1(n_5786),
.B2(n_4762),
.C(n_5353),
.Y(n_5909)
);

NAND2xp5_ASAP7_75t_L g5910 ( 
.A(n_5820),
.B(n_5753),
.Y(n_5910)
);

HB1xp67_ASAP7_75t_L g5911 ( 
.A(n_5871),
.Y(n_5911)
);

AND2x2_ASAP7_75t_L g5912 ( 
.A(n_5854),
.B(n_5787),
.Y(n_5912)
);

AND2x4_ASAP7_75t_L g5913 ( 
.A(n_5823),
.B(n_5012),
.Y(n_5913)
);

NAND3xp33_ASAP7_75t_L g5914 ( 
.A(n_5858),
.B(n_5409),
.C(n_5065),
.Y(n_5914)
);

BUFx3_ASAP7_75t_L g5915 ( 
.A(n_5863),
.Y(n_5915)
);

INVx2_ASAP7_75t_SL g5916 ( 
.A(n_5849),
.Y(n_5916)
);

AND2x4_ASAP7_75t_L g5917 ( 
.A(n_5854),
.B(n_5044),
.Y(n_5917)
);

NAND2xp5_ASAP7_75t_SL g5918 ( 
.A(n_5859),
.B(n_4674),
.Y(n_5918)
);

OAI222xp33_ASAP7_75t_L g5919 ( 
.A1(n_5824),
.A2(n_5860),
.B1(n_5855),
.B2(n_5821),
.C1(n_5840),
.C2(n_5875),
.Y(n_5919)
);

INVx3_ASAP7_75t_L g5920 ( 
.A(n_5841),
.Y(n_5920)
);

INVx1_ASAP7_75t_L g5921 ( 
.A(n_5848),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_5843),
.Y(n_5922)
);

INVxp67_ASAP7_75t_L g5923 ( 
.A(n_5864),
.Y(n_5923)
);

INVx2_ASAP7_75t_L g5924 ( 
.A(n_5844),
.Y(n_5924)
);

INVx2_ASAP7_75t_L g5925 ( 
.A(n_5850),
.Y(n_5925)
);

AOI33xp33_ASAP7_75t_L g5926 ( 
.A1(n_5851),
.A2(n_4907),
.A3(n_5053),
.B1(n_5054),
.B2(n_4917),
.B3(n_4911),
.Y(n_5926)
);

AND2x2_ASAP7_75t_L g5927 ( 
.A(n_5837),
.B(n_5137),
.Y(n_5927)
);

INVx2_ASAP7_75t_L g5928 ( 
.A(n_5862),
.Y(n_5928)
);

OAI31xp33_ASAP7_75t_L g5929 ( 
.A1(n_5836),
.A2(n_5206),
.A3(n_5370),
.B(n_5199),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5817),
.Y(n_5930)
);

HB1xp67_ASAP7_75t_L g5931 ( 
.A(n_5848),
.Y(n_5931)
);

AND2x2_ASAP7_75t_SL g5932 ( 
.A(n_5853),
.B(n_5151),
.Y(n_5932)
);

AND2x4_ASAP7_75t_L g5933 ( 
.A(n_5829),
.B(n_5005),
.Y(n_5933)
);

AOI211xp5_ASAP7_75t_L g5934 ( 
.A1(n_5831),
.A2(n_5364),
.B(n_5367),
.C(n_5366),
.Y(n_5934)
);

AND2x2_ASAP7_75t_L g5935 ( 
.A(n_5861),
.B(n_5818),
.Y(n_5935)
);

AOI21xp5_ASAP7_75t_L g5936 ( 
.A1(n_5833),
.A2(n_4744),
.B(n_5034),
.Y(n_5936)
);

INVx3_ASAP7_75t_L g5937 ( 
.A(n_5819),
.Y(n_5937)
);

INVx1_ASAP7_75t_L g5938 ( 
.A(n_5856),
.Y(n_5938)
);

INVx2_ASAP7_75t_L g5939 ( 
.A(n_5856),
.Y(n_5939)
);

INVx2_ASAP7_75t_L g5940 ( 
.A(n_5873),
.Y(n_5940)
);

AND2x4_ASAP7_75t_L g5941 ( 
.A(n_5852),
.B(n_5005),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5873),
.Y(n_5942)
);

AND2x4_ASAP7_75t_L g5943 ( 
.A(n_5865),
.B(n_5867),
.Y(n_5943)
);

INVxp67_ASAP7_75t_L g5944 ( 
.A(n_5868),
.Y(n_5944)
);

OR2x2_ASAP7_75t_L g5945 ( 
.A(n_5888),
.B(n_5839),
.Y(n_5945)
);

INVx2_ASAP7_75t_L g5946 ( 
.A(n_5892),
.Y(n_5946)
);

NAND2xp5_ASAP7_75t_L g5947 ( 
.A(n_5923),
.B(n_5826),
.Y(n_5947)
);

OR2x6_ASAP7_75t_L g5948 ( 
.A(n_5885),
.B(n_5369),
.Y(n_5948)
);

AND2x2_ASAP7_75t_L g5949 ( 
.A(n_5878),
.B(n_5853),
.Y(n_5949)
);

NAND2xp5_ASAP7_75t_L g5950 ( 
.A(n_5883),
.B(n_5874),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5931),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5889),
.Y(n_5952)
);

AND2x2_ASAP7_75t_L g5953 ( 
.A(n_5884),
.B(n_5908),
.Y(n_5953)
);

INVx2_ASAP7_75t_L g5954 ( 
.A(n_5937),
.Y(n_5954)
);

NOR4xp25_ASAP7_75t_SL g5955 ( 
.A(n_5896),
.B(n_5827),
.C(n_5016),
.D(n_5405),
.Y(n_5955)
);

INVx2_ASAP7_75t_SL g5956 ( 
.A(n_5904),
.Y(n_5956)
);

NAND3xp33_ASAP7_75t_L g5957 ( 
.A(n_5905),
.B(n_5874),
.C(n_5067),
.Y(n_5957)
);

OR2x2_ASAP7_75t_L g5958 ( 
.A(n_5902),
.B(n_5197),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5920),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5893),
.Y(n_5960)
);

INVx2_ASAP7_75t_L g5961 ( 
.A(n_5876),
.Y(n_5961)
);

INVx2_ASAP7_75t_L g5962 ( 
.A(n_5877),
.Y(n_5962)
);

AND2x2_ASAP7_75t_L g5963 ( 
.A(n_5897),
.B(n_5064),
.Y(n_5963)
);

INVx2_ASAP7_75t_L g5964 ( 
.A(n_5886),
.Y(n_5964)
);

INVxp33_ASAP7_75t_L g5965 ( 
.A(n_5891),
.Y(n_5965)
);

INVx3_ASAP7_75t_L g5966 ( 
.A(n_5890),
.Y(n_5966)
);

NAND2xp5_ASAP7_75t_L g5967 ( 
.A(n_5916),
.B(n_5187),
.Y(n_5967)
);

AND2x4_ASAP7_75t_L g5968 ( 
.A(n_5882),
.B(n_4696),
.Y(n_5968)
);

HB1xp67_ASAP7_75t_L g5969 ( 
.A(n_5894),
.Y(n_5969)
);

INVx3_ASAP7_75t_L g5970 ( 
.A(n_5890),
.Y(n_5970)
);

INVx2_ASAP7_75t_L g5971 ( 
.A(n_5890),
.Y(n_5971)
);

INVx2_ASAP7_75t_L g5972 ( 
.A(n_5899),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5939),
.Y(n_5973)
);

INVx1_ASAP7_75t_L g5974 ( 
.A(n_5921),
.Y(n_5974)
);

INVxp67_ASAP7_75t_L g5975 ( 
.A(n_5896),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_SL g5976 ( 
.A(n_5881),
.B(n_5057),
.Y(n_5976)
);

AND2x2_ASAP7_75t_L g5977 ( 
.A(n_5913),
.B(n_5402),
.Y(n_5977)
);

AND2x2_ASAP7_75t_L g5978 ( 
.A(n_5913),
.B(n_5407),
.Y(n_5978)
);

NOR2x1_ASAP7_75t_SL g5979 ( 
.A(n_5918),
.B(n_5270),
.Y(n_5979)
);

INVx2_ASAP7_75t_SL g5980 ( 
.A(n_5915),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5940),
.Y(n_5981)
);

INVx1_ASAP7_75t_L g5982 ( 
.A(n_5938),
.Y(n_5982)
);

NAND2xp5_ASAP7_75t_L g5983 ( 
.A(n_5929),
.B(n_5198),
.Y(n_5983)
);

HB1xp67_ASAP7_75t_L g5984 ( 
.A(n_5944),
.Y(n_5984)
);

AND2x4_ASAP7_75t_SL g5985 ( 
.A(n_5901),
.B(n_5094),
.Y(n_5985)
);

NAND2xp5_ASAP7_75t_L g5986 ( 
.A(n_5927),
.B(n_5198),
.Y(n_5986)
);

NAND2xp5_ASAP7_75t_L g5987 ( 
.A(n_5943),
.B(n_5181),
.Y(n_5987)
);

AOI21xp33_ASAP7_75t_SL g5988 ( 
.A1(n_5909),
.A2(n_5388),
.B(n_5361),
.Y(n_5988)
);

AND2x4_ASAP7_75t_L g5989 ( 
.A(n_5956),
.B(n_5980),
.Y(n_5989)
);

NAND2xp5_ASAP7_75t_L g5990 ( 
.A(n_5946),
.B(n_5943),
.Y(n_5990)
);

NAND2xp5_ASAP7_75t_L g5991 ( 
.A(n_5988),
.B(n_5898),
.Y(n_5991)
);

AND2x2_ASAP7_75t_L g5992 ( 
.A(n_5953),
.B(n_5912),
.Y(n_5992)
);

INVxp67_ASAP7_75t_L g5993 ( 
.A(n_5971),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5984),
.Y(n_5994)
);

OR2x2_ASAP7_75t_L g5995 ( 
.A(n_5945),
.B(n_5895),
.Y(n_5995)
);

OR2x6_ASAP7_75t_L g5996 ( 
.A(n_5948),
.B(n_5900),
.Y(n_5996)
);

AOI21xp33_ASAP7_75t_SL g5997 ( 
.A1(n_5965),
.A2(n_5903),
.B(n_5900),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5951),
.Y(n_5998)
);

AND2x2_ASAP7_75t_L g5999 ( 
.A(n_5954),
.B(n_5907),
.Y(n_5999)
);

INVx1_ASAP7_75t_L g6000 ( 
.A(n_5947),
.Y(n_6000)
);

OR2x2_ASAP7_75t_L g6001 ( 
.A(n_5969),
.B(n_5911),
.Y(n_6001)
);

INVx1_ASAP7_75t_L g6002 ( 
.A(n_5982),
.Y(n_6002)
);

AND2x2_ASAP7_75t_L g6003 ( 
.A(n_5959),
.B(n_5966),
.Y(n_6003)
);

AND2x2_ASAP7_75t_L g6004 ( 
.A(n_5966),
.B(n_5906),
.Y(n_6004)
);

HB1xp67_ASAP7_75t_L g6005 ( 
.A(n_5961),
.Y(n_6005)
);

BUFx2_ASAP7_75t_L g6006 ( 
.A(n_5970),
.Y(n_6006)
);

INVx1_ASAP7_75t_SL g6007 ( 
.A(n_5968),
.Y(n_6007)
);

OR2x2_ASAP7_75t_L g6008 ( 
.A(n_5962),
.B(n_5930),
.Y(n_6008)
);

NAND2xp5_ASAP7_75t_L g6009 ( 
.A(n_5983),
.B(n_5936),
.Y(n_6009)
);

NAND2xp5_ASAP7_75t_L g6010 ( 
.A(n_5975),
.B(n_5887),
.Y(n_6010)
);

NOR2x1_ASAP7_75t_L g6011 ( 
.A(n_5970),
.B(n_5903),
.Y(n_6011)
);

NAND2xp5_ASAP7_75t_L g6012 ( 
.A(n_5952),
.B(n_5941),
.Y(n_6012)
);

AND2x2_ASAP7_75t_L g6013 ( 
.A(n_5977),
.B(n_5935),
.Y(n_6013)
);

INVx2_ASAP7_75t_L g6014 ( 
.A(n_5964),
.Y(n_6014)
);

NAND2xp5_ASAP7_75t_L g6015 ( 
.A(n_5960),
.B(n_5941),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5982),
.Y(n_6016)
);

AND2x2_ASAP7_75t_L g6017 ( 
.A(n_5978),
.B(n_5917),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5974),
.Y(n_6018)
);

NAND2xp5_ASAP7_75t_L g6019 ( 
.A(n_5972),
.B(n_5942),
.Y(n_6019)
);

NOR2xp33_ASAP7_75t_L g6020 ( 
.A(n_5968),
.B(n_5880),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5973),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_5973),
.Y(n_6022)
);

AND2x2_ASAP7_75t_L g6023 ( 
.A(n_5949),
.B(n_5917),
.Y(n_6023)
);

INVx1_ASAP7_75t_L g6024 ( 
.A(n_5981),
.Y(n_6024)
);

INVxp67_ASAP7_75t_L g6025 ( 
.A(n_5979),
.Y(n_6025)
);

AND2x2_ASAP7_75t_L g6026 ( 
.A(n_5989),
.B(n_5992),
.Y(n_6026)
);

BUFx3_ASAP7_75t_L g6027 ( 
.A(n_5989),
.Y(n_6027)
);

NAND2xp5_ASAP7_75t_L g6028 ( 
.A(n_5993),
.B(n_5948),
.Y(n_6028)
);

NAND2xp5_ASAP7_75t_L g6029 ( 
.A(n_6020),
.B(n_5950),
.Y(n_6029)
);

INVx4_ASAP7_75t_L g6030 ( 
.A(n_6006),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_6005),
.Y(n_6031)
);

AND2x2_ASAP7_75t_L g6032 ( 
.A(n_6004),
.B(n_5985),
.Y(n_6032)
);

AND2x4_ASAP7_75t_L g6033 ( 
.A(n_6007),
.B(n_5963),
.Y(n_6033)
);

HB1xp67_ASAP7_75t_L g6034 ( 
.A(n_5994),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_6021),
.Y(n_6035)
);

BUFx2_ASAP7_75t_L g6036 ( 
.A(n_6011),
.Y(n_6036)
);

INVx1_ASAP7_75t_SL g6037 ( 
.A(n_6003),
.Y(n_6037)
);

INVx2_ASAP7_75t_L g6038 ( 
.A(n_6001),
.Y(n_6038)
);

NAND2xp33_ASAP7_75t_L g6039 ( 
.A(n_6000),
.B(n_5990),
.Y(n_6039)
);

BUFx3_ASAP7_75t_L g6040 ( 
.A(n_6014),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5999),
.B(n_6023),
.Y(n_6041)
);

AND3x1_ASAP7_75t_L g6042 ( 
.A(n_5991),
.B(n_5955),
.C(n_5934),
.Y(n_6042)
);

INVx2_ASAP7_75t_L g6043 ( 
.A(n_6008),
.Y(n_6043)
);

OR2x6_ASAP7_75t_L g6044 ( 
.A(n_5996),
.B(n_5933),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_6022),
.Y(n_6045)
);

INVx1_ASAP7_75t_L g6046 ( 
.A(n_6024),
.Y(n_6046)
);

CKINVDCx16_ASAP7_75t_R g6047 ( 
.A(n_5996),
.Y(n_6047)
);

OR2x2_ASAP7_75t_L g6048 ( 
.A(n_5995),
.B(n_5986),
.Y(n_6048)
);

AOI22xp33_ASAP7_75t_L g6049 ( 
.A1(n_6009),
.A2(n_5879),
.B1(n_5957),
.B2(n_5933),
.Y(n_6049)
);

INVx1_ASAP7_75t_SL g6050 ( 
.A(n_5998),
.Y(n_6050)
);

OR2x2_ASAP7_75t_L g6051 ( 
.A(n_6019),
.B(n_5958),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_6002),
.Y(n_6052)
);

OR2x2_ASAP7_75t_L g6053 ( 
.A(n_6010),
.B(n_5967),
.Y(n_6053)
);

AND2x2_ASAP7_75t_L g6054 ( 
.A(n_6013),
.B(n_5979),
.Y(n_6054)
);

NAND3x1_ASAP7_75t_L g6055 ( 
.A(n_5997),
.B(n_5981),
.C(n_5987),
.Y(n_6055)
);

INVx2_ASAP7_75t_SL g6056 ( 
.A(n_6012),
.Y(n_6056)
);

INVx2_ASAP7_75t_L g6057 ( 
.A(n_6015),
.Y(n_6057)
);

INVx2_ASAP7_75t_L g6058 ( 
.A(n_6018),
.Y(n_6058)
);

INVx2_ASAP7_75t_L g6059 ( 
.A(n_6017),
.Y(n_6059)
);

OR2x2_ASAP7_75t_L g6060 ( 
.A(n_6016),
.B(n_5922),
.Y(n_6060)
);

AND2x2_ASAP7_75t_L g6061 ( 
.A(n_6025),
.B(n_5910),
.Y(n_6061)
);

AND2x2_ASAP7_75t_L g6062 ( 
.A(n_5989),
.B(n_5924),
.Y(n_6062)
);

A2O1A1Ixp33_ASAP7_75t_SL g6063 ( 
.A1(n_6025),
.A2(n_5925),
.B(n_5928),
.C(n_5070),
.Y(n_6063)
);

AND2x2_ASAP7_75t_L g6064 ( 
.A(n_5989),
.B(n_5914),
.Y(n_6064)
);

AND2x2_ASAP7_75t_L g6065 ( 
.A(n_5989),
.B(n_5932),
.Y(n_6065)
);

INVx2_ASAP7_75t_L g6066 ( 
.A(n_5989),
.Y(n_6066)
);

INVxp67_ASAP7_75t_SL g6067 ( 
.A(n_6027),
.Y(n_6067)
);

OR2x2_ASAP7_75t_L g6068 ( 
.A(n_6038),
.B(n_5976),
.Y(n_6068)
);

BUFx2_ASAP7_75t_L g6069 ( 
.A(n_6066),
.Y(n_6069)
);

INVx2_ASAP7_75t_SL g6070 ( 
.A(n_6062),
.Y(n_6070)
);

AND2x2_ASAP7_75t_L g6071 ( 
.A(n_6026),
.B(n_5926),
.Y(n_6071)
);

INVxp67_ASAP7_75t_L g6072 ( 
.A(n_6036),
.Y(n_6072)
);

NAND2xp33_ASAP7_75t_L g6073 ( 
.A(n_6037),
.B(n_5042),
.Y(n_6073)
);

OR2x2_ASAP7_75t_L g6074 ( 
.A(n_6031),
.B(n_668),
.Y(n_6074)
);

NAND2xp5_ASAP7_75t_L g6075 ( 
.A(n_6030),
.B(n_669),
.Y(n_6075)
);

INVxp67_ASAP7_75t_L g6076 ( 
.A(n_6040),
.Y(n_6076)
);

AND2x2_ASAP7_75t_L g6077 ( 
.A(n_6041),
.B(n_5919),
.Y(n_6077)
);

NAND4xp25_ASAP7_75t_SL g6078 ( 
.A(n_6029),
.B(n_5245),
.C(n_5046),
.D(n_4904),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_6034),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_6043),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_6030),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_6060),
.Y(n_6082)
);

NAND2xp5_ASAP7_75t_L g6083 ( 
.A(n_6056),
.B(n_669),
.Y(n_6083)
);

AND2x2_ASAP7_75t_L g6084 ( 
.A(n_6032),
.B(n_5321),
.Y(n_6084)
);

NAND2xp5_ASAP7_75t_L g6085 ( 
.A(n_6057),
.B(n_670),
.Y(n_6085)
);

NOR2xp33_ASAP7_75t_L g6086 ( 
.A(n_6047),
.B(n_671),
.Y(n_6086)
);

AND2x2_ASAP7_75t_L g6087 ( 
.A(n_6064),
.B(n_5309),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_6051),
.Y(n_6088)
);

NAND2xp33_ASAP7_75t_L g6089 ( 
.A(n_6028),
.B(n_4906),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_6039),
.Y(n_6090)
);

AND2x2_ASAP7_75t_L g6091 ( 
.A(n_6065),
.B(n_5310),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_6035),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_6035),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_6045),
.Y(n_6094)
);

HB1xp67_ASAP7_75t_L g6095 ( 
.A(n_6045),
.Y(n_6095)
);

BUFx2_ASAP7_75t_L g6096 ( 
.A(n_6033),
.Y(n_6096)
);

NAND2xp5_ASAP7_75t_L g6097 ( 
.A(n_6050),
.B(n_671),
.Y(n_6097)
);

INVx1_ASAP7_75t_L g6098 ( 
.A(n_6046),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_6046),
.Y(n_6099)
);

AND2x2_ASAP7_75t_L g6100 ( 
.A(n_6033),
.B(n_5311),
.Y(n_6100)
);

INVx1_ASAP7_75t_L g6101 ( 
.A(n_6061),
.Y(n_6101)
);

INVx1_ASAP7_75t_L g6102 ( 
.A(n_6048),
.Y(n_6102)
);

AND2x2_ASAP7_75t_L g6103 ( 
.A(n_6054),
.B(n_5314),
.Y(n_6103)
);

INVx2_ASAP7_75t_L g6104 ( 
.A(n_6059),
.Y(n_6104)
);

INVx2_ASAP7_75t_L g6105 ( 
.A(n_6058),
.Y(n_6105)
);

NAND2xp5_ASAP7_75t_L g6106 ( 
.A(n_6052),
.B(n_671),
.Y(n_6106)
);

INVxp67_ASAP7_75t_SL g6107 ( 
.A(n_6076),
.Y(n_6107)
);

AOI22xp5_ASAP7_75t_L g6108 ( 
.A1(n_6067),
.A2(n_6042),
.B1(n_6055),
.B2(n_6053),
.Y(n_6108)
);

NOR2xp33_ASAP7_75t_L g6109 ( 
.A(n_6096),
.B(n_6052),
.Y(n_6109)
);

INVx1_ASAP7_75t_L g6110 ( 
.A(n_6081),
.Y(n_6110)
);

INVx1_ASAP7_75t_SL g6111 ( 
.A(n_6069),
.Y(n_6111)
);

AOI211xp5_ASAP7_75t_L g6112 ( 
.A1(n_6072),
.A2(n_6063),
.B(n_6049),
.C(n_6044),
.Y(n_6112)
);

NOR2xp33_ASAP7_75t_L g6113 ( 
.A(n_6070),
.B(n_6044),
.Y(n_6113)
);

INVx1_ASAP7_75t_L g6114 ( 
.A(n_6075),
.Y(n_6114)
);

OAI22xp5_ASAP7_75t_L g6115 ( 
.A1(n_6090),
.A2(n_5094),
.B1(n_4927),
.B2(n_5015),
.Y(n_6115)
);

OAI211xp5_ASAP7_75t_L g6116 ( 
.A1(n_6080),
.A2(n_5399),
.B(n_5384),
.C(n_5400),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_6068),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_6086),
.Y(n_6118)
);

NAND2xp5_ASAP7_75t_L g6119 ( 
.A(n_6077),
.B(n_6071),
.Y(n_6119)
);

INVxp67_ASAP7_75t_L g6120 ( 
.A(n_6097),
.Y(n_6120)
);

AOI21xp5_ASAP7_75t_L g6121 ( 
.A1(n_6097),
.A2(n_5395),
.B(n_5344),
.Y(n_6121)
);

NOR2xp33_ASAP7_75t_L g6122 ( 
.A(n_6101),
.B(n_672),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_6083),
.Y(n_6123)
);

OR2x2_ASAP7_75t_L g6124 ( 
.A(n_6104),
.B(n_672),
.Y(n_6124)
);

AOI21xp5_ASAP7_75t_L g6125 ( 
.A1(n_6106),
.A2(n_5351),
.B(n_5334),
.Y(n_6125)
);

INVx3_ASAP7_75t_L g6126 ( 
.A(n_6105),
.Y(n_6126)
);

INVx1_ASAP7_75t_L g6127 ( 
.A(n_6074),
.Y(n_6127)
);

NAND2xp5_ASAP7_75t_L g6128 ( 
.A(n_6100),
.B(n_672),
.Y(n_6128)
);

INVx1_ASAP7_75t_L g6129 ( 
.A(n_6082),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_6088),
.Y(n_6130)
);

OR2x2_ASAP7_75t_L g6131 ( 
.A(n_6085),
.B(n_673),
.Y(n_6131)
);

AOI22xp5_ASAP7_75t_L g6132 ( 
.A1(n_6102),
.A2(n_4650),
.B1(n_5062),
.B2(n_5358),
.Y(n_6132)
);

AOI22xp5_ASAP7_75t_L g6133 ( 
.A1(n_6084),
.A2(n_5184),
.B1(n_5185),
.B2(n_5193),
.Y(n_6133)
);

NAND2xp5_ASAP7_75t_L g6134 ( 
.A(n_6087),
.B(n_673),
.Y(n_6134)
);

NAND2xp5_ASAP7_75t_SL g6135 ( 
.A(n_6079),
.B(n_5265),
.Y(n_6135)
);

AOI221xp5_ASAP7_75t_L g6136 ( 
.A1(n_6095),
.A2(n_4926),
.B1(n_4881),
.B2(n_4880),
.C(n_4875),
.Y(n_6136)
);

INVx2_ASAP7_75t_SL g6137 ( 
.A(n_6103),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_6106),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_6073),
.Y(n_6139)
);

OR2x2_ASAP7_75t_L g6140 ( 
.A(n_6091),
.B(n_674),
.Y(n_6140)
);

NAND2xp5_ASAP7_75t_L g6141 ( 
.A(n_6089),
.B(n_6092),
.Y(n_6141)
);

O2A1O1Ixp33_ASAP7_75t_L g6142 ( 
.A1(n_6093),
.A2(n_676),
.B(n_674),
.C(n_675),
.Y(n_6142)
);

O2A1O1Ixp33_ASAP7_75t_L g6143 ( 
.A1(n_6094),
.A2(n_677),
.B(n_675),
.C(n_676),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_6098),
.Y(n_6144)
);

INVx2_ASAP7_75t_SL g6145 ( 
.A(n_6099),
.Y(n_6145)
);

NAND2x1p5_ASAP7_75t_L g6146 ( 
.A(n_6078),
.B(n_5230),
.Y(n_6146)
);

INVx2_ASAP7_75t_SL g6147 ( 
.A(n_6069),
.Y(n_6147)
);

OAI322xp33_ASAP7_75t_L g6148 ( 
.A1(n_6072),
.A2(n_4827),
.A3(n_4926),
.B1(n_683),
.B2(n_680),
.C1(n_682),
.C2(n_678),
.Y(n_6148)
);

HB1xp67_ASAP7_75t_L g6149 ( 
.A(n_6081),
.Y(n_6149)
);

AOI21xp5_ASAP7_75t_L g6150 ( 
.A1(n_6067),
.A2(n_5325),
.B(n_5299),
.Y(n_6150)
);

AOI222xp33_ASAP7_75t_L g6151 ( 
.A1(n_6067),
.A2(n_5234),
.B1(n_5247),
.B2(n_5257),
.C1(n_5229),
.C2(n_5057),
.Y(n_6151)
);

AOI21xp33_ASAP7_75t_SL g6152 ( 
.A1(n_6076),
.A2(n_679),
.B(n_680),
.Y(n_6152)
);

AOI221xp5_ASAP7_75t_L g6153 ( 
.A1(n_6067),
.A2(n_4875),
.B1(n_4881),
.B2(n_4880),
.C(n_4782),
.Y(n_6153)
);

AOI222xp33_ASAP7_75t_L g6154 ( 
.A1(n_6067),
.A2(n_5221),
.B1(n_5134),
.B2(n_5211),
.C1(n_5210),
.C2(n_5113),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_6096),
.Y(n_6155)
);

NOR2x1_ASAP7_75t_L g6156 ( 
.A(n_6075),
.B(n_681),
.Y(n_6156)
);

NOR3xp33_ASAP7_75t_SL g6157 ( 
.A(n_6067),
.B(n_682),
.C(n_683),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_6067),
.Y(n_6158)
);

INVx1_ASAP7_75t_L g6159 ( 
.A(n_6067),
.Y(n_6159)
);

NAND2x1_ASAP7_75t_L g6160 ( 
.A(n_6096),
.B(n_5151),
.Y(n_6160)
);

INVxp67_ASAP7_75t_L g6161 ( 
.A(n_6113),
.Y(n_6161)
);

INVx2_ASAP7_75t_SL g6162 ( 
.A(n_6158),
.Y(n_6162)
);

NAND2xp5_ASAP7_75t_L g6163 ( 
.A(n_6159),
.B(n_682),
.Y(n_6163)
);

INVx1_ASAP7_75t_L g6164 ( 
.A(n_6107),
.Y(n_6164)
);

OR2x2_ASAP7_75t_L g6165 ( 
.A(n_6111),
.B(n_683),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_6149),
.Y(n_6166)
);

NAND2xp5_ASAP7_75t_L g6167 ( 
.A(n_6147),
.B(n_684),
.Y(n_6167)
);

INVx2_ASAP7_75t_L g6168 ( 
.A(n_6155),
.Y(n_6168)
);

NAND2xp5_ASAP7_75t_L g6169 ( 
.A(n_6119),
.B(n_684),
.Y(n_6169)
);

INVx1_ASAP7_75t_L g6170 ( 
.A(n_6126),
.Y(n_6170)
);

INVxp67_ASAP7_75t_SL g6171 ( 
.A(n_6126),
.Y(n_6171)
);

OR2x2_ASAP7_75t_L g6172 ( 
.A(n_6117),
.B(n_6124),
.Y(n_6172)
);

INVx2_ASAP7_75t_L g6173 ( 
.A(n_6110),
.Y(n_6173)
);

AND2x2_ASAP7_75t_L g6174 ( 
.A(n_6157),
.B(n_684),
.Y(n_6174)
);

NAND2xp5_ASAP7_75t_L g6175 ( 
.A(n_6112),
.B(n_685),
.Y(n_6175)
);

OR2x2_ASAP7_75t_L g6176 ( 
.A(n_6134),
.B(n_685),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_6128),
.Y(n_6177)
);

NAND2xp5_ASAP7_75t_L g6178 ( 
.A(n_6152),
.B(n_685),
.Y(n_6178)
);

NOR2xp33_ASAP7_75t_L g6179 ( 
.A(n_6108),
.B(n_686),
.Y(n_6179)
);

INVx1_ASAP7_75t_L g6180 ( 
.A(n_6131),
.Y(n_6180)
);

NOR2xp33_ASAP7_75t_L g6181 ( 
.A(n_6137),
.B(n_686),
.Y(n_6181)
);

INVx2_ASAP7_75t_SL g6182 ( 
.A(n_6129),
.Y(n_6182)
);

NAND2xp5_ASAP7_75t_L g6183 ( 
.A(n_6109),
.B(n_686),
.Y(n_6183)
);

AND2x2_ASAP7_75t_L g6184 ( 
.A(n_6118),
.B(n_6139),
.Y(n_6184)
);

NAND2xp5_ASAP7_75t_L g6185 ( 
.A(n_6146),
.B(n_687),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_6140),
.Y(n_6186)
);

AOI21xp5_ASAP7_75t_SL g6187 ( 
.A1(n_6142),
.A2(n_687),
.B(n_688),
.Y(n_6187)
);

NAND2xp5_ASAP7_75t_SL g6188 ( 
.A(n_6130),
.B(n_4674),
.Y(n_6188)
);

AOI21xp5_ASAP7_75t_L g6189 ( 
.A1(n_6143),
.A2(n_5177),
.B(n_687),
.Y(n_6189)
);

NAND2xp5_ASAP7_75t_L g6190 ( 
.A(n_6125),
.B(n_688),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_6156),
.Y(n_6191)
);

NAND2xp5_ASAP7_75t_L g6192 ( 
.A(n_6121),
.B(n_688),
.Y(n_6192)
);

AND2x2_ASAP7_75t_L g6193 ( 
.A(n_6127),
.B(n_689),
.Y(n_6193)
);

INVx1_ASAP7_75t_L g6194 ( 
.A(n_6141),
.Y(n_6194)
);

NAND2xp5_ASAP7_75t_L g6195 ( 
.A(n_6122),
.B(n_689),
.Y(n_6195)
);

NAND2xp5_ASAP7_75t_SL g6196 ( 
.A(n_6145),
.B(n_4689),
.Y(n_6196)
);

NAND2xp5_ASAP7_75t_SL g6197 ( 
.A(n_6138),
.B(n_6120),
.Y(n_6197)
);

AND2x2_ASAP7_75t_L g6198 ( 
.A(n_6114),
.B(n_690),
.Y(n_6198)
);

INVxp67_ASAP7_75t_L g6199 ( 
.A(n_6144),
.Y(n_6199)
);

AND2x2_ASAP7_75t_L g6200 ( 
.A(n_6123),
.B(n_690),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_6148),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_6135),
.Y(n_6202)
);

NOR2xp33_ASAP7_75t_L g6203 ( 
.A(n_6115),
.B(n_690),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_6150),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_6171),
.Y(n_6205)
);

AOI221xp5_ASAP7_75t_L g6206 ( 
.A1(n_6201),
.A2(n_6153),
.B1(n_6160),
.B2(n_6133),
.C(n_6116),
.Y(n_6206)
);

INVx2_ASAP7_75t_L g6207 ( 
.A(n_6168),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_6165),
.Y(n_6208)
);

NOR3x1_ASAP7_75t_L g6209 ( 
.A(n_6169),
.B(n_6132),
.C(n_6154),
.Y(n_6209)
);

NAND2xp5_ASAP7_75t_L g6210 ( 
.A(n_6174),
.B(n_6164),
.Y(n_6210)
);

INVxp67_ASAP7_75t_L g6211 ( 
.A(n_6181),
.Y(n_6211)
);

AND2x4_ASAP7_75t_L g6212 ( 
.A(n_6162),
.B(n_6136),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_6167),
.Y(n_6213)
);

NAND2xp5_ASAP7_75t_L g6214 ( 
.A(n_6170),
.B(n_6151),
.Y(n_6214)
);

NAND2xp5_ASAP7_75t_L g6215 ( 
.A(n_6166),
.B(n_691),
.Y(n_6215)
);

NAND2xp5_ASAP7_75t_SL g6216 ( 
.A(n_6175),
.B(n_6183),
.Y(n_6216)
);

OR2x2_ASAP7_75t_L g6217 ( 
.A(n_6185),
.B(n_691),
.Y(n_6217)
);

NAND2xp5_ASAP7_75t_SL g6218 ( 
.A(n_6183),
.B(n_4689),
.Y(n_6218)
);

NAND2xp5_ASAP7_75t_L g6219 ( 
.A(n_6179),
.B(n_691),
.Y(n_6219)
);

INVx1_ASAP7_75t_L g6220 ( 
.A(n_6172),
.Y(n_6220)
);

INVx2_ASAP7_75t_L g6221 ( 
.A(n_6173),
.Y(n_6221)
);

NAND2xp5_ASAP7_75t_L g6222 ( 
.A(n_6161),
.B(n_692),
.Y(n_6222)
);

OR2x2_ASAP7_75t_L g6223 ( 
.A(n_6163),
.B(n_692),
.Y(n_6223)
);

OA22x2_ASAP7_75t_L g6224 ( 
.A1(n_6187),
.A2(n_5115),
.B1(n_5160),
.B2(n_5194),
.Y(n_6224)
);

AND2x2_ASAP7_75t_L g6225 ( 
.A(n_6193),
.B(n_692),
.Y(n_6225)
);

NAND3xp33_ASAP7_75t_L g6226 ( 
.A(n_6194),
.B(n_693),
.C(n_694),
.Y(n_6226)
);

INVx1_ASAP7_75t_L g6227 ( 
.A(n_6198),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_6200),
.B(n_693),
.Y(n_6228)
);

A2O1A1Ixp33_ASAP7_75t_L g6229 ( 
.A1(n_6203),
.A2(n_5169),
.B(n_5153),
.C(n_5157),
.Y(n_6229)
);

NAND2xp5_ASAP7_75t_L g6230 ( 
.A(n_6204),
.B(n_6189),
.Y(n_6230)
);

NAND2xp5_ASAP7_75t_L g6231 ( 
.A(n_6184),
.B(n_694),
.Y(n_6231)
);

AOI31xp67_ASAP7_75t_SL g6232 ( 
.A1(n_6190),
.A2(n_6192),
.A3(n_6186),
.B(n_6202),
.Y(n_6232)
);

AOI211x1_ASAP7_75t_L g6233 ( 
.A1(n_6197),
.A2(n_696),
.B(n_694),
.C(n_695),
.Y(n_6233)
);

OR3x1_ASAP7_75t_L g6234 ( 
.A(n_6180),
.B(n_695),
.C(n_696),
.Y(n_6234)
);

NAND2x1_ASAP7_75t_SL g6235 ( 
.A(n_6191),
.B(n_696),
.Y(n_6235)
);

NAND2x1_ASAP7_75t_SL g6236 ( 
.A(n_6177),
.B(n_697),
.Y(n_6236)
);

INVx1_ASAP7_75t_L g6237 ( 
.A(n_6178),
.Y(n_6237)
);

NAND2xp5_ASAP7_75t_L g6238 ( 
.A(n_6182),
.B(n_697),
.Y(n_6238)
);

AND2x2_ASAP7_75t_L g6239 ( 
.A(n_6176),
.B(n_698),
.Y(n_6239)
);

AOI22xp33_ASAP7_75t_SL g6240 ( 
.A1(n_6199),
.A2(n_4782),
.B1(n_4776),
.B2(n_4802),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_6195),
.Y(n_6241)
);

INVx1_ASAP7_75t_L g6242 ( 
.A(n_6188),
.Y(n_6242)
);

NAND2xp5_ASAP7_75t_L g6243 ( 
.A(n_6196),
.B(n_698),
.Y(n_6243)
);

AOI21xp5_ASAP7_75t_L g6244 ( 
.A1(n_6187),
.A2(n_698),
.B(n_699),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_6171),
.Y(n_6245)
);

NOR2xp33_ASAP7_75t_L g6246 ( 
.A(n_6201),
.B(n_699),
.Y(n_6246)
);

NAND2xp5_ASAP7_75t_L g6247 ( 
.A(n_6171),
.B(n_700),
.Y(n_6247)
);

INVxp33_ASAP7_75t_L g6248 ( 
.A(n_6181),
.Y(n_6248)
);

NOR2xp33_ASAP7_75t_L g6249 ( 
.A(n_6201),
.B(n_700),
.Y(n_6249)
);

NAND2xp5_ASAP7_75t_L g6250 ( 
.A(n_6171),
.B(n_701),
.Y(n_6250)
);

O2A1O1Ixp33_ASAP7_75t_L g6251 ( 
.A1(n_6207),
.A2(n_703),
.B(n_701),
.C(n_702),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_6205),
.Y(n_6252)
);

XNOR2xp5_ASAP7_75t_L g6253 ( 
.A(n_6234),
.B(n_701),
.Y(n_6253)
);

NAND2xp5_ASAP7_75t_L g6254 ( 
.A(n_6245),
.B(n_702),
.Y(n_6254)
);

NAND2xp5_ASAP7_75t_SL g6255 ( 
.A(n_6212),
.B(n_4734),
.Y(n_6255)
);

BUFx2_ASAP7_75t_L g6256 ( 
.A(n_6235),
.Y(n_6256)
);

INVx1_ASAP7_75t_SL g6257 ( 
.A(n_6220),
.Y(n_6257)
);

NOR2xp33_ASAP7_75t_L g6258 ( 
.A(n_6231),
.B(n_702),
.Y(n_6258)
);

NAND2xp5_ASAP7_75t_L g6259 ( 
.A(n_6246),
.B(n_6249),
.Y(n_6259)
);

O2A1O1Ixp33_ASAP7_75t_L g6260 ( 
.A1(n_6247),
.A2(n_706),
.B(n_704),
.C(n_705),
.Y(n_6260)
);

NAND2xp5_ASAP7_75t_L g6261 ( 
.A(n_6225),
.B(n_704),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_6250),
.Y(n_6262)
);

NAND2xp5_ASAP7_75t_SL g6263 ( 
.A(n_6212),
.B(n_4734),
.Y(n_6263)
);

NOR2xp33_ASAP7_75t_L g6264 ( 
.A(n_6228),
.B(n_704),
.Y(n_6264)
);

OR2x2_ASAP7_75t_L g6265 ( 
.A(n_6243),
.B(n_706),
.Y(n_6265)
);

NOR4xp25_ASAP7_75t_L g6266 ( 
.A(n_6232),
.B(n_708),
.C(n_706),
.D(n_707),
.Y(n_6266)
);

AOI21xp5_ASAP7_75t_L g6267 ( 
.A1(n_6244),
.A2(n_707),
.B(n_708),
.Y(n_6267)
);

NAND2xp5_ASAP7_75t_SL g6268 ( 
.A(n_6206),
.B(n_4738),
.Y(n_6268)
);

NOR2xp33_ASAP7_75t_L g6269 ( 
.A(n_6248),
.B(n_708),
.Y(n_6269)
);

AND2x2_ASAP7_75t_L g6270 ( 
.A(n_6239),
.B(n_709),
.Y(n_6270)
);

AOI21xp5_ASAP7_75t_L g6271 ( 
.A1(n_6230),
.A2(n_709),
.B(n_710),
.Y(n_6271)
);

NAND4xp25_ASAP7_75t_L g6272 ( 
.A(n_6210),
.B(n_711),
.C(n_709),
.D(n_710),
.Y(n_6272)
);

NAND4xp75_ASAP7_75t_L g6273 ( 
.A(n_6233),
.B(n_6238),
.C(n_6215),
.D(n_6222),
.Y(n_6273)
);

NOR3x1_ASAP7_75t_L g6274 ( 
.A(n_6226),
.B(n_710),
.C(n_711),
.Y(n_6274)
);

NAND5xp2_ASAP7_75t_L g6275 ( 
.A(n_6227),
.B(n_713),
.C(n_711),
.D(n_712),
.E(n_714),
.Y(n_6275)
);

NOR3xp33_ASAP7_75t_SL g6276 ( 
.A(n_6216),
.B(n_712),
.C(n_713),
.Y(n_6276)
);

NOR2xp33_ASAP7_75t_L g6277 ( 
.A(n_6221),
.B(n_713),
.Y(n_6277)
);

NAND2xp5_ASAP7_75t_L g6278 ( 
.A(n_6208),
.B(n_714),
.Y(n_6278)
);

O2A1O1Ixp33_ASAP7_75t_L g6279 ( 
.A1(n_6219),
.A2(n_716),
.B(n_714),
.C(n_715),
.Y(n_6279)
);

AND2x2_ASAP7_75t_L g6280 ( 
.A(n_6240),
.B(n_715),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_6236),
.Y(n_6281)
);

NAND2xp5_ASAP7_75t_L g6282 ( 
.A(n_6242),
.B(n_6237),
.Y(n_6282)
);

NAND2xp5_ASAP7_75t_L g6283 ( 
.A(n_6211),
.B(n_715),
.Y(n_6283)
);

NOR2xp33_ASAP7_75t_L g6284 ( 
.A(n_6214),
.B(n_716),
.Y(n_6284)
);

AOI221xp5_ASAP7_75t_L g6285 ( 
.A1(n_6218),
.A2(n_718),
.B1(n_716),
.B2(n_717),
.C(n_719),
.Y(n_6285)
);

INVx1_ASAP7_75t_L g6286 ( 
.A(n_6223),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_6217),
.Y(n_6287)
);

OR2x2_ASAP7_75t_L g6288 ( 
.A(n_6213),
.B(n_717),
.Y(n_6288)
);

INVx2_ASAP7_75t_L g6289 ( 
.A(n_6224),
.Y(n_6289)
);

NAND4xp25_ASAP7_75t_L g6290 ( 
.A(n_6209),
.B(n_720),
.C(n_717),
.D(n_718),
.Y(n_6290)
);

NOR2xp33_ASAP7_75t_SL g6291 ( 
.A(n_6257),
.B(n_6241),
.Y(n_6291)
);

NAND2xp5_ASAP7_75t_SL g6292 ( 
.A(n_6266),
.B(n_6229),
.Y(n_6292)
);

AOI321xp33_ASAP7_75t_L g6293 ( 
.A1(n_6268),
.A2(n_6284),
.A3(n_6263),
.B1(n_6255),
.B2(n_6252),
.C(n_6282),
.Y(n_6293)
);

AOI222xp33_ASAP7_75t_L g6294 ( 
.A1(n_6280),
.A2(n_4806),
.B1(n_4821),
.B2(n_4804),
.C1(n_4776),
.C2(n_4743),
.Y(n_6294)
);

OAI221xp5_ASAP7_75t_L g6295 ( 
.A1(n_6285),
.A2(n_722),
.B1(n_720),
.B2(n_721),
.C(n_723),
.Y(n_6295)
);

AOI222xp33_ASAP7_75t_SL g6296 ( 
.A1(n_6287),
.A2(n_724),
.B1(n_726),
.B2(n_721),
.C1(n_722),
.C2(n_725),
.Y(n_6296)
);

AOI221xp5_ASAP7_75t_L g6297 ( 
.A1(n_6251),
.A2(n_725),
.B1(n_721),
.B2(n_724),
.C(n_726),
.Y(n_6297)
);

NAND2xp5_ASAP7_75t_L g6298 ( 
.A(n_6253),
.B(n_725),
.Y(n_6298)
);

NOR2xp33_ASAP7_75t_SL g6299 ( 
.A(n_6269),
.B(n_4738),
.Y(n_6299)
);

OAI221xp5_ASAP7_75t_L g6300 ( 
.A1(n_6290),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.C(n_729),
.Y(n_6300)
);

AOI211x1_ASAP7_75t_SL g6301 ( 
.A1(n_6259),
.A2(n_730),
.B(n_727),
.C(n_729),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_6254),
.Y(n_6302)
);

O2A1O1Ixp33_ASAP7_75t_L g6303 ( 
.A1(n_6260),
.A2(n_731),
.B(n_727),
.C(n_730),
.Y(n_6303)
);

OAI211xp5_ASAP7_75t_L g6304 ( 
.A1(n_6272),
.A2(n_733),
.B(n_730),
.C(n_732),
.Y(n_6304)
);

AOI21xp5_ASAP7_75t_L g6305 ( 
.A1(n_6267),
.A2(n_732),
.B(n_733),
.Y(n_6305)
);

OAI211xp5_ASAP7_75t_SL g6306 ( 
.A1(n_6276),
.A2(n_6278),
.B(n_6271),
.C(n_6279),
.Y(n_6306)
);

NOR3xp33_ASAP7_75t_L g6307 ( 
.A(n_6283),
.B(n_734),
.C(n_735),
.Y(n_6307)
);

NAND4xp75_ASAP7_75t_L g6308 ( 
.A(n_6274),
.B(n_736),
.C(n_734),
.D(n_735),
.Y(n_6308)
);

INVx2_ASAP7_75t_L g6309 ( 
.A(n_6265),
.Y(n_6309)
);

AOI222xp33_ASAP7_75t_L g6310 ( 
.A1(n_6277),
.A2(n_4814),
.B1(n_4753),
.B2(n_4819),
.C1(n_4807),
.C2(n_4743),
.Y(n_6310)
);

O2A1O1Ixp33_ASAP7_75t_L g6311 ( 
.A1(n_6281),
.A2(n_737),
.B(n_734),
.C(n_736),
.Y(n_6311)
);

A2O1A1Ixp33_ASAP7_75t_L g6312 ( 
.A1(n_6258),
.A2(n_5125),
.B(n_5142),
.C(n_5170),
.Y(n_6312)
);

OAI221xp5_ASAP7_75t_L g6313 ( 
.A1(n_6261),
.A2(n_738),
.B1(n_736),
.B2(n_737),
.C(n_739),
.Y(n_6313)
);

OAI222xp33_ASAP7_75t_L g6314 ( 
.A1(n_6288),
.A2(n_740),
.B1(n_742),
.B2(n_738),
.C1(n_739),
.C2(n_741),
.Y(n_6314)
);

NOR2xp33_ASAP7_75t_R g6315 ( 
.A(n_6256),
.B(n_738),
.Y(n_6315)
);

AOI211xp5_ASAP7_75t_SL g6316 ( 
.A1(n_6264),
.A2(n_741),
.B(n_739),
.C(n_740),
.Y(n_6316)
);

AOI22xp5_ASAP7_75t_L g6317 ( 
.A1(n_6270),
.A2(n_5197),
.B1(n_4807),
.B2(n_4814),
.Y(n_6317)
);

AOI211xp5_ASAP7_75t_L g6318 ( 
.A1(n_6275),
.A2(n_742),
.B(n_740),
.C(n_741),
.Y(n_6318)
);

INVx1_ASAP7_75t_L g6319 ( 
.A(n_6289),
.Y(n_6319)
);

O2A1O1Ixp33_ASAP7_75t_L g6320 ( 
.A1(n_6286),
.A2(n_745),
.B(n_743),
.C(n_744),
.Y(n_6320)
);

AOI211xp5_ASAP7_75t_L g6321 ( 
.A1(n_6262),
.A2(n_745),
.B(n_743),
.C(n_744),
.Y(n_6321)
);

AOI221xp5_ASAP7_75t_L g6322 ( 
.A1(n_6273),
.A2(n_746),
.B1(n_743),
.B2(n_744),
.C(n_747),
.Y(n_6322)
);

INVx1_ASAP7_75t_SL g6323 ( 
.A(n_6257),
.Y(n_6323)
);

O2A1O1Ixp33_ASAP7_75t_L g6324 ( 
.A1(n_6251),
.A2(n_748),
.B(n_746),
.C(n_747),
.Y(n_6324)
);

AOI22xp33_ASAP7_75t_L g6325 ( 
.A1(n_6319),
.A2(n_4913),
.B1(n_4922),
.B2(n_4909),
.Y(n_6325)
);

NOR2x1_ASAP7_75t_L g6326 ( 
.A(n_6308),
.B(n_747),
.Y(n_6326)
);

OAI211xp5_ASAP7_75t_SL g6327 ( 
.A1(n_6300),
.A2(n_750),
.B(n_748),
.C(n_749),
.Y(n_6327)
);

AOI221xp5_ASAP7_75t_L g6328 ( 
.A1(n_6311),
.A2(n_750),
.B1(n_748),
.B2(n_749),
.C(n_751),
.Y(n_6328)
);

OAI221xp5_ASAP7_75t_L g6329 ( 
.A1(n_6322),
.A2(n_751),
.B1(n_749),
.B2(n_750),
.C(n_752),
.Y(n_6329)
);

INVx2_ASAP7_75t_L g6330 ( 
.A(n_6323),
.Y(n_6330)
);

NAND4xp25_ASAP7_75t_SL g6331 ( 
.A(n_6318),
.B(n_755),
.C(n_753),
.D(n_754),
.Y(n_6331)
);

XOR2x2_ASAP7_75t_L g6332 ( 
.A(n_6316),
.B(n_753),
.Y(n_6332)
);

INVx2_ASAP7_75t_L g6333 ( 
.A(n_6309),
.Y(n_6333)
);

AOI221xp5_ASAP7_75t_L g6334 ( 
.A1(n_6314),
.A2(n_755),
.B1(n_753),
.B2(n_754),
.C(n_756),
.Y(n_6334)
);

AOI22xp5_ASAP7_75t_L g6335 ( 
.A1(n_6291),
.A2(n_4819),
.B1(n_4753),
.B2(n_4798),
.Y(n_6335)
);

NOR3xp33_ASAP7_75t_SL g6336 ( 
.A(n_6313),
.B(n_754),
.C(n_756),
.Y(n_6336)
);

AOI221xp5_ASAP7_75t_L g6337 ( 
.A1(n_6320),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.C(n_760),
.Y(n_6337)
);

AOI221xp5_ASAP7_75t_L g6338 ( 
.A1(n_6295),
.A2(n_6324),
.B1(n_6303),
.B2(n_6297),
.C(n_6304),
.Y(n_6338)
);

AOI21xp5_ASAP7_75t_L g6339 ( 
.A1(n_6292),
.A2(n_757),
.B(n_758),
.Y(n_6339)
);

A2O1A1Ixp33_ASAP7_75t_L g6340 ( 
.A1(n_6305),
.A2(n_759),
.B(n_757),
.C(n_758),
.Y(n_6340)
);

AOI21xp5_ASAP7_75t_L g6341 ( 
.A1(n_6298),
.A2(n_760),
.B(n_761),
.Y(n_6341)
);

NOR3xp33_ASAP7_75t_L g6342 ( 
.A(n_6306),
.B(n_760),
.C(n_761),
.Y(n_6342)
);

AOI221xp5_ASAP7_75t_L g6343 ( 
.A1(n_6307),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.C(n_765),
.Y(n_6343)
);

AOI22xp5_ASAP7_75t_L g6344 ( 
.A1(n_6296),
.A2(n_4798),
.B1(n_5141),
.B2(n_4913),
.Y(n_6344)
);

NOR3xp33_ASAP7_75t_L g6345 ( 
.A(n_6321),
.B(n_762),
.C(n_764),
.Y(n_6345)
);

AND4x1_ASAP7_75t_L g6346 ( 
.A(n_6301),
.B(n_6299),
.C(n_6302),
.D(n_6294),
.Y(n_6346)
);

XNOR2xp5_ASAP7_75t_L g6347 ( 
.A(n_6317),
.B(n_762),
.Y(n_6347)
);

NOR2xp33_ASAP7_75t_L g6348 ( 
.A(n_6330),
.B(n_6293),
.Y(n_6348)
);

AOI221x1_ASAP7_75t_L g6349 ( 
.A1(n_6342),
.A2(n_6315),
.B1(n_6312),
.B2(n_6310),
.C(n_766),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_6326),
.Y(n_6350)
);

INVx2_ASAP7_75t_L g6351 ( 
.A(n_6333),
.Y(n_6351)
);

NOR2xp33_ASAP7_75t_L g6352 ( 
.A(n_6327),
.B(n_764),
.Y(n_6352)
);

AOI22xp5_ASAP7_75t_L g6353 ( 
.A1(n_6331),
.A2(n_4798),
.B1(n_4922),
.B2(n_4909),
.Y(n_6353)
);

NAND2xp5_ASAP7_75t_L g6354 ( 
.A(n_6339),
.B(n_765),
.Y(n_6354)
);

NAND2xp5_ASAP7_75t_SL g6355 ( 
.A(n_6338),
.B(n_765),
.Y(n_6355)
);

OAI221xp5_ASAP7_75t_L g6356 ( 
.A1(n_6328),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.C(n_769),
.Y(n_6356)
);

AOI31xp33_ASAP7_75t_L g6357 ( 
.A1(n_6343),
.A2(n_768),
.A3(n_766),
.B(n_767),
.Y(n_6357)
);

AND2x4_ASAP7_75t_L g6358 ( 
.A(n_6346),
.B(n_768),
.Y(n_6358)
);

NAND2xp5_ASAP7_75t_SL g6359 ( 
.A(n_6334),
.B(n_770),
.Y(n_6359)
);

NOR3xp33_ASAP7_75t_L g6360 ( 
.A(n_6329),
.B(n_770),
.C(n_771),
.Y(n_6360)
);

OAI211xp5_ASAP7_75t_L g6361 ( 
.A1(n_6337),
.A2(n_772),
.B(n_770),
.C(n_771),
.Y(n_6361)
);

AOI22xp5_ASAP7_75t_SL g6362 ( 
.A1(n_6347),
.A2(n_773),
.B1(n_771),
.B2(n_772),
.Y(n_6362)
);

A2O1A1Ixp33_ASAP7_75t_L g6363 ( 
.A1(n_6341),
.A2(n_774),
.B(n_772),
.C(n_773),
.Y(n_6363)
);

OAI221xp5_ASAP7_75t_L g6364 ( 
.A1(n_6340),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.C(n_777),
.Y(n_6364)
);

NAND2xp5_ASAP7_75t_L g6365 ( 
.A(n_6345),
.B(n_6332),
.Y(n_6365)
);

OAI22xp5_ASAP7_75t_L g6366 ( 
.A1(n_6336),
.A2(n_778),
.B1(n_775),
.B2(n_777),
.Y(n_6366)
);

INVx1_ASAP7_75t_SL g6367 ( 
.A(n_6335),
.Y(n_6367)
);

NAND2xp5_ASAP7_75t_L g6368 ( 
.A(n_6325),
.B(n_775),
.Y(n_6368)
);

INVx1_ASAP7_75t_L g6369 ( 
.A(n_6344),
.Y(n_6369)
);

NOR4xp25_ASAP7_75t_L g6370 ( 
.A(n_6351),
.B(n_779),
.C(n_777),
.D(n_778),
.Y(n_6370)
);

NOR3xp33_ASAP7_75t_SL g6371 ( 
.A(n_6355),
.B(n_779),
.C(n_780),
.Y(n_6371)
);

NAND3xp33_ASAP7_75t_SL g6372 ( 
.A(n_6360),
.B(n_779),
.C(n_780),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_6354),
.Y(n_6373)
);

CKINVDCx8_ASAP7_75t_R g6374 ( 
.A(n_6358),
.Y(n_6374)
);

NAND2x1p5_ASAP7_75t_L g6375 ( 
.A(n_6367),
.B(n_780),
.Y(n_6375)
);

AOI221xp5_ASAP7_75t_L g6376 ( 
.A1(n_6357),
.A2(n_783),
.B1(n_781),
.B2(n_782),
.C(n_784),
.Y(n_6376)
);

INVx2_ASAP7_75t_SL g6377 ( 
.A(n_6358),
.Y(n_6377)
);

XNOR2x1_ASAP7_75t_L g6378 ( 
.A(n_6366),
.B(n_781),
.Y(n_6378)
);

NAND5xp2_ASAP7_75t_L g6379 ( 
.A(n_6348),
.B(n_784),
.C(n_782),
.D(n_783),
.E(n_785),
.Y(n_6379)
);

NOR2xp67_ASAP7_75t_L g6380 ( 
.A(n_6369),
.B(n_782),
.Y(n_6380)
);

NOR3xp33_ASAP7_75t_L g6381 ( 
.A(n_6361),
.B(n_785),
.C(n_786),
.Y(n_6381)
);

AND2x4_ASAP7_75t_L g6382 ( 
.A(n_6350),
.B(n_785),
.Y(n_6382)
);

NAND3xp33_ASAP7_75t_L g6383 ( 
.A(n_6352),
.B(n_786),
.C(n_787),
.Y(n_6383)
);

INVx1_ASAP7_75t_L g6384 ( 
.A(n_6368),
.Y(n_6384)
);

AND4x1_ASAP7_75t_L g6385 ( 
.A(n_6365),
.B(n_789),
.C(n_786),
.D(n_788),
.Y(n_6385)
);

NOR3xp33_ASAP7_75t_L g6386 ( 
.A(n_6364),
.B(n_6356),
.C(n_6359),
.Y(n_6386)
);

NOR2xp33_ASAP7_75t_L g6387 ( 
.A(n_6362),
.B(n_788),
.Y(n_6387)
);

NAND2x1p5_ASAP7_75t_L g6388 ( 
.A(n_6377),
.B(n_6349),
.Y(n_6388)
);

BUFx6f_ASAP7_75t_L g6389 ( 
.A(n_6374),
.Y(n_6389)
);

CKINVDCx5p33_ASAP7_75t_R g6390 ( 
.A(n_6371),
.Y(n_6390)
);

CKINVDCx5p33_ASAP7_75t_R g6391 ( 
.A(n_6382),
.Y(n_6391)
);

AOI21xp5_ASAP7_75t_L g6392 ( 
.A1(n_6378),
.A2(n_6363),
.B(n_6387),
.Y(n_6392)
);

INVx1_ASAP7_75t_L g6393 ( 
.A(n_6375),
.Y(n_6393)
);

NOR3xp33_ASAP7_75t_L g6394 ( 
.A(n_6372),
.B(n_6353),
.C(n_788),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_6380),
.Y(n_6395)
);

NAND3xp33_ASAP7_75t_SL g6396 ( 
.A(n_6376),
.B(n_789),
.C(n_790),
.Y(n_6396)
);

HB1xp67_ASAP7_75t_L g6397 ( 
.A(n_6385),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_6388),
.Y(n_6398)
);

INVx2_ASAP7_75t_L g6399 ( 
.A(n_6389),
.Y(n_6399)
);

AOI22xp5_ASAP7_75t_L g6400 ( 
.A1(n_6390),
.A2(n_6386),
.B1(n_6381),
.B2(n_6383),
.Y(n_6400)
);

XNOR2xp5_ASAP7_75t_L g6401 ( 
.A(n_6391),
.B(n_6370),
.Y(n_6401)
);

AND3x1_ASAP7_75t_L g6402 ( 
.A(n_6394),
.B(n_6379),
.C(n_6384),
.Y(n_6402)
);

AO21x2_ASAP7_75t_L g6403 ( 
.A1(n_6392),
.A2(n_6373),
.B(n_790),
.Y(n_6403)
);

AOI21xp5_ASAP7_75t_L g6404 ( 
.A1(n_6396),
.A2(n_790),
.B(n_791),
.Y(n_6404)
);

HB1xp67_ASAP7_75t_L g6405 ( 
.A(n_6389),
.Y(n_6405)
);

OAI22xp5_ASAP7_75t_L g6406 ( 
.A1(n_6393),
.A2(n_793),
.B1(n_791),
.B2(n_792),
.Y(n_6406)
);

INVx1_ASAP7_75t_L g6407 ( 
.A(n_6397),
.Y(n_6407)
);

OAI22xp33_ASAP7_75t_L g6408 ( 
.A1(n_6398),
.A2(n_6395),
.B1(n_793),
.B2(n_791),
.Y(n_6408)
);

OAI21xp5_ASAP7_75t_L g6409 ( 
.A1(n_6404),
.A2(n_792),
.B(n_793),
.Y(n_6409)
);

HB1xp67_ASAP7_75t_L g6410 ( 
.A(n_6403),
.Y(n_6410)
);

INVx1_ASAP7_75t_L g6411 ( 
.A(n_6406),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_6408),
.Y(n_6412)
);

AOI22x1_ASAP7_75t_L g6413 ( 
.A1(n_6412),
.A2(n_6401),
.B1(n_6407),
.B2(n_6405),
.Y(n_6413)
);

OAI21xp5_ASAP7_75t_L g6414 ( 
.A1(n_6413),
.A2(n_6399),
.B(n_6400),
.Y(n_6414)
);

OAI22xp5_ASAP7_75t_L g6415 ( 
.A1(n_6413),
.A2(n_6402),
.B1(n_6411),
.B2(n_6410),
.Y(n_6415)
);

OAI22xp5_ASAP7_75t_L g6416 ( 
.A1(n_6414),
.A2(n_6409),
.B1(n_795),
.B2(n_792),
.Y(n_6416)
);

INVx4_ASAP7_75t_L g6417 ( 
.A(n_6415),
.Y(n_6417)
);

NAND3xp33_ASAP7_75t_SL g6418 ( 
.A(n_6417),
.B(n_794),
.C(n_795),
.Y(n_6418)
);

AOI222xp33_ASAP7_75t_SL g6419 ( 
.A1(n_6416),
.A2(n_796),
.B1(n_798),
.B2(n_794),
.C1(n_795),
.C2(n_797),
.Y(n_6419)
);

OAI222xp33_ASAP7_75t_L g6420 ( 
.A1(n_6418),
.A2(n_798),
.B1(n_800),
.B2(n_796),
.C1(n_797),
.C2(n_799),
.Y(n_6420)
);

AOI22xp33_ASAP7_75t_L g6421 ( 
.A1(n_6419),
.A2(n_798),
.B1(n_796),
.B2(n_797),
.Y(n_6421)
);

AOI22xp33_ASAP7_75t_L g6422 ( 
.A1(n_6418),
.A2(n_801),
.B1(n_799),
.B2(n_800),
.Y(n_6422)
);

OAI21xp5_ASAP7_75t_L g6423 ( 
.A1(n_6422),
.A2(n_799),
.B(n_800),
.Y(n_6423)
);

OA21x2_ASAP7_75t_L g6424 ( 
.A1(n_6421),
.A2(n_801),
.B(n_802),
.Y(n_6424)
);

OR2x2_ASAP7_75t_L g6425 ( 
.A(n_6420),
.B(n_802),
.Y(n_6425)
);

AOI21xp5_ASAP7_75t_L g6426 ( 
.A1(n_6425),
.A2(n_6423),
.B(n_6424),
.Y(n_6426)
);

AOI211xp5_ASAP7_75t_L g6427 ( 
.A1(n_6426),
.A2(n_806),
.B(n_803),
.C(n_805),
.Y(n_6427)
);


endmodule