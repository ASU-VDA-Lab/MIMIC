module fake_jpeg_2184_n_247 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_247);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_2),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_20),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_62),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_64),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_69),
.B(n_71),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_72),
.B(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_32),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_81),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_92),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_30),
.B1(n_24),
.B2(n_36),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_44),
.A2(n_36),
.B1(n_35),
.B2(n_30),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_40),
.B1(n_38),
.B2(n_25),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_93),
.B1(n_55),
.B2(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_38),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_21),
.B1(n_1),
.B2(n_3),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_21),
.Y(n_97)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_127),
.Y(n_147)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_11),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_129),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_91),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_99),
.C(n_89),
.Y(n_134)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_126),
.Y(n_139)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_130),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_96),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_14),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_0),
.Y(n_146)
);

CKINVDCx12_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_132),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_121),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_83),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_140),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_111),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_84),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_150),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_85),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_95),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_155),
.B(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_95),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_96),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_168),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_130),
.B1(n_125),
.B2(n_116),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_176),
.B1(n_145),
.B2(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_108),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_103),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_173),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_163),
.C(n_174),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_173),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_148),
.B1(n_149),
.B2(n_151),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_194),
.A2(n_160),
.B1(n_158),
.B2(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_190),
.B(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_195),
.B(n_202),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_198),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_206),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_164),
.C(n_172),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_208),
.C(n_179),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_171),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_148),
.C(n_151),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_215),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_182),
.C(n_180),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_191),
.C(n_193),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_203),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_221),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_SL g222 ( 
.A(n_218),
.B(n_184),
.C(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_216),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_223),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_226),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_184),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_227),
.B1(n_211),
.B2(n_215),
.Y(n_229)
);

A2O1A1O1Ixp25_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_194),
.B(n_192),
.C(n_196),
.D(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_224),
.C(n_213),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_209),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_236),
.C(n_239),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_159),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_233),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_231),
.B1(n_237),
.B2(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_222),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_241),
.A2(n_7),
.B1(n_176),
.B2(n_240),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_176),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_244),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_246),
.Y(n_247)
);


endmodule