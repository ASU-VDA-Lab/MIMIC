module fake_jpeg_23470_n_325 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_25),
.Y(n_40)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_14),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_52),
.B(n_30),
.C(n_29),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_23),
.B1(n_13),
.B2(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_13),
.B1(n_23),
.B2(n_27),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_16),
.B(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_23),
.B1(n_14),
.B2(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_60),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_62),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_64),
.B(n_73),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_48),
.B1(n_32),
.B2(n_38),
.Y(n_96)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_14),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_38),
.B1(n_32),
.B2(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_34),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_54),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_34),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_87),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_97),
.B1(n_32),
.B2(n_47),
.Y(n_123)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_43),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_40),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_99),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_59),
.A2(n_57),
.B1(n_61),
.B2(n_66),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_37),
.C(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_86),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_71),
.Y(n_114)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_105),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_93),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_59),
.B1(n_49),
.B2(n_55),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_103),
.B(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_119),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_109),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_55),
.B1(n_69),
.B2(n_49),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_111),
.B1(n_118),
.B2(n_122),
.Y(n_125)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_68),
.B1(n_44),
.B2(n_29),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_44),
.B1(n_35),
.B2(n_37),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_95),
.B1(n_99),
.B2(n_80),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_94),
.B1(n_65),
.B2(n_82),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_126),
.A2(n_127),
.B(n_129),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_128),
.B(n_120),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_88),
.B(n_44),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_133),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_68),
.B1(n_92),
.B2(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_56),
.B1(n_51),
.B2(n_29),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_138),
.A2(n_103),
.B1(n_122),
.B2(n_108),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_30),
.Y(n_139)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_30),
.B1(n_51),
.B2(n_56),
.Y(n_141)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_106),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_150),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_109),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_118),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_117),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_155),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_113),
.C(n_121),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_137),
.C(n_138),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_22),
.B1(n_20),
.B2(n_26),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_116),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_113),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_122),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_113),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_105),
.B(n_93),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_28),
.B(n_21),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_141),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_105),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_174),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_111),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_111),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_51),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_178),
.Y(n_199)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_180),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_182),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_129),
.C(n_127),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_127),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_193),
.B1(n_198),
.B2(n_200),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_135),
.B1(n_131),
.B2(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_194),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_125),
.B1(n_130),
.B2(n_147),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_195),
.B1(n_197),
.B2(n_203),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_169),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_166),
.A2(n_130),
.B1(n_83),
.B2(n_26),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_79),
.B1(n_56),
.B2(n_63),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_170),
.B(n_28),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_172),
.B(n_165),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_171),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_79),
.B1(n_76),
.B2(n_15),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_208),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_163),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_204),
.B(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_152),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_160),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_220),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_153),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_223),
.C(n_225),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_193),
.B(n_160),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_222),
.B1(n_176),
.B2(n_168),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_153),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_151),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_158),
.B1(n_168),
.B2(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_192),
.C(n_175),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_24),
.B(n_21),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_182),
.C(n_183),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_233),
.C(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_181),
.C(n_198),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_185),
.B1(n_165),
.B2(n_161),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_246),
.B1(n_210),
.B2(n_215),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_176),
.B1(n_158),
.B2(n_200),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_202),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_247),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_177),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_162),
.C(n_173),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_228),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_178),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_218),
.B1(n_223),
.B2(n_219),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_205),
.A2(n_195),
.B1(n_203),
.B2(n_22),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_219),
.B(n_210),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_250),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_259),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_206),
.B1(n_216),
.B2(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_206),
.B(n_20),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_260),
.C(n_261),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_247),
.B(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_236),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_15),
.B1(n_21),
.B2(n_24),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_9),
.B(n_12),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_11),
.B1(n_21),
.B2(n_15),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_264),
.C(n_243),
.Y(n_275)
);

AO22x1_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_24),
.B1(n_15),
.B2(n_4),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_24),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_232),
.C(n_233),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_277),
.C(n_278),
.Y(n_282)
);

BUFx12_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_250),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_258),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_279),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_240),
.C(n_238),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_235),
.C(n_230),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_28),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_249),
.Y(n_286)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_251),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_285),
.B(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_263),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_293),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g287 ( 
.A(n_269),
.B(n_265),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_248),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_289),
.B(n_290),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_272),
.A2(n_261),
.B(n_254),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_28),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_268),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_4),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_280),
.C(n_271),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_297),
.C(n_5),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_292),
.A2(n_271),
.B(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_283),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_281),
.B(n_3),
.Y(n_300)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_0),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_303),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_19),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_5),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_312),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_5),
.B(n_6),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_19),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_299),
.B(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_297),
.C(n_311),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.C(n_316),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_301),
.C(n_307),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_313),
.B1(n_307),
.B2(n_8),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_6),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_6),
.C(n_7),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_7),
.B(n_8),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_7),
.B(n_8),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_7),
.B(n_19),
.Y(n_325)
);


endmodule