module real_aes_7138_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g116 ( .A(n_0), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_1), .A2(n_458), .B1(n_459), .B2(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_1), .Y(n_458) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_2), .A2(n_149), .B(n_154), .C(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_3), .A2(n_144), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g506 ( .A(n_4), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_5), .B(n_182), .Y(n_248) );
AOI21xp33_ASAP7_75t_L g513 ( .A1(n_6), .A2(n_144), .B(n_514), .Y(n_513) );
AND2x6_ASAP7_75t_L g149 ( .A(n_7), .B(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_8), .A2(n_279), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g161 ( .A(n_9), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_10), .B(n_43), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_11), .A2(n_33), .B1(n_461), .B2(n_462), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_11), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_12), .B(n_159), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_13), .B(n_206), .Y(n_485) );
INVx1_ASAP7_75t_L g518 ( .A(n_14), .Y(n_518) );
INVx1_ASAP7_75t_L g142 ( .A(n_15), .Y(n_142) );
INVx1_ASAP7_75t_L g497 ( .A(n_16), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_17), .A2(n_162), .B(n_176), .C(n_180), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_18), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_19), .B(n_476), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_20), .B(n_144), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_21), .B(n_288), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_22), .A2(n_206), .B(n_207), .C(n_209), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_23), .B(n_182), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_24), .B(n_159), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_25), .A2(n_178), .B(n_180), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_26), .B(n_159), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_27), .Y(n_230) );
INVx1_ASAP7_75t_L g218 ( .A(n_28), .Y(n_218) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_29), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_30), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_31), .B(n_159), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_32), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g461 ( .A(n_33), .Y(n_461) );
INVx1_ASAP7_75t_L g284 ( .A(n_34), .Y(n_284) );
INVx1_ASAP7_75t_L g526 ( .A(n_35), .Y(n_526) );
INVx2_ASAP7_75t_L g147 ( .A(n_36), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_37), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_38), .A2(n_206), .B(n_244), .C(n_246), .Y(n_243) );
INVxp67_ASAP7_75t_L g285 ( .A(n_39), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_40), .A2(n_154), .B(n_217), .C(n_223), .Y(n_216) );
CKINVDCx14_ASAP7_75t_R g242 ( .A(n_41), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_42), .A2(n_149), .B(n_154), .C(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g525 ( .A(n_44), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g157 ( .A1(n_45), .A2(n_158), .B(n_160), .C(n_163), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_46), .B(n_159), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_47), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_48), .Y(n_281) );
INVx1_ASAP7_75t_L g204 ( .A(n_49), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_50), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_51), .B(n_144), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_52), .A2(n_154), .B1(n_209), .B2(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_53), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_54), .Y(n_503) );
CKINVDCx14_ASAP7_75t_R g152 ( .A(n_55), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_56), .A2(n_158), .B(n_246), .C(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_57), .Y(n_563) );
INVx1_ASAP7_75t_L g515 ( .A(n_58), .Y(n_515) );
INVx1_ASAP7_75t_L g150 ( .A(n_59), .Y(n_150) );
INVx1_ASAP7_75t_L g141 ( .A(n_60), .Y(n_141) );
INVx1_ASAP7_75t_SL g245 ( .A(n_61), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_62), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_63), .B(n_182), .Y(n_211) );
INVx1_ASAP7_75t_L g233 ( .A(n_64), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_SL g534 ( .A1(n_65), .A2(n_246), .B(n_476), .C(n_535), .Y(n_534) );
INVxp67_ASAP7_75t_L g536 ( .A(n_66), .Y(n_536) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_68), .A2(n_144), .B(n_151), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_69), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_70), .A2(n_144), .B(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_71), .Y(n_529) );
INVx1_ASAP7_75t_L g557 ( .A(n_72), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_73), .A2(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g174 ( .A(n_74), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_75), .Y(n_215) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_76), .A2(n_77), .B1(n_445), .B2(n_446), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_76), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_77), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_78), .A2(n_149), .B(n_154), .C(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_SL g452 ( .A1(n_79), .A2(n_114), .B1(n_453), .B2(n_746), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_80), .A2(n_144), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g177 ( .A(n_81), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_82), .B(n_219), .Y(n_474) );
INVx2_ASAP7_75t_L g139 ( .A(n_83), .Y(n_139) );
INVx1_ASAP7_75t_L g193 ( .A(n_84), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_85), .B(n_476), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_86), .A2(n_149), .B(n_154), .C(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g125 ( .A(n_87), .B(n_114), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_88), .A2(n_154), .B(n_232), .C(n_235), .Y(n_231) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_89), .A2(n_91), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_89), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_90), .B(n_138), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_91), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_92), .A2(n_149), .B(n_154), .C(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_93), .Y(n_489) );
INVx1_ASAP7_75t_L g533 ( .A(n_94), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_95), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_96), .B(n_219), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_97), .A2(n_105), .B1(n_118), .B2(n_750), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_98), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_99), .B(n_167), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_100), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g208 ( .A(n_101), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_102), .A2(n_455), .B1(n_456), .B2(n_457), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_102), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_103), .A2(n_144), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g751 ( .A(n_108), .Y(n_751) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx3_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g747 ( .A(n_112), .Y(n_747) );
NOR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g744 ( .A(n_113), .Y(n_744) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B(n_451), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g749 ( .A(n_121), .Y(n_749) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_126), .B(n_448), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_125), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_130), .B1(n_131), .B2(n_447), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_127), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_128), .B(n_187), .Y(n_509) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
XOR2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_444), .Y(n_131) );
INVx2_ASAP7_75t_L g745 ( .A(n_132), .Y(n_745) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_374), .Y(n_132) );
NAND5xp2_ASAP7_75t_L g133 ( .A(n_134), .B(n_289), .C(n_321), .D(n_338), .E(n_361), .Y(n_133) );
AOI221xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_212), .B1(n_249), .B2(n_253), .C(n_257), .Y(n_134) );
INVx1_ASAP7_75t_L g401 ( .A(n_135), .Y(n_401) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_184), .Y(n_135) );
AND3x2_ASAP7_75t_L g376 ( .A(n_136), .B(n_186), .C(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_169), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_137), .B(n_255), .Y(n_254) );
BUFx3_ASAP7_75t_L g264 ( .A(n_137), .Y(n_264) );
AND2x2_ASAP7_75t_L g268 ( .A(n_137), .B(n_200), .Y(n_268) );
INVx2_ASAP7_75t_L g298 ( .A(n_137), .Y(n_298) );
OR2x2_ASAP7_75t_L g309 ( .A(n_137), .B(n_201), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_137), .B(n_185), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_137), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g388 ( .A(n_137), .B(n_201), .Y(n_388) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_143), .B(n_166), .Y(n_137) );
INVx1_ASAP7_75t_L g187 ( .A(n_138), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_138), .A2(n_190), .B(n_215), .C(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g238 ( .A(n_138), .Y(n_238) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_138), .A2(n_492), .B(n_498), .Y(n_491) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_L g168 ( .A(n_139), .B(n_140), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx2_ASAP7_75t_L g279 ( .A(n_144), .Y(n_279) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_145), .B(n_149), .Y(n_190) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g222 ( .A(n_146), .Y(n_222) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
INVx1_ASAP7_75t_L g210 ( .A(n_147), .Y(n_210) );
INVx1_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_148), .Y(n_162) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
INVx1_ASAP7_75t_L g476 ( .A(n_148), .Y(n_476) );
INVx4_ASAP7_75t_SL g165 ( .A(n_149), .Y(n_165) );
BUFx3_ASAP7_75t_L g223 ( .A(n_149), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_SL g151 ( .A1(n_152), .A2(n_153), .B(n_157), .C(n_165), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_153), .A2(n_165), .B(n_174), .C(n_175), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g203 ( .A1(n_153), .A2(n_165), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_153), .A2(n_165), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g280 ( .A1(n_153), .A2(n_165), .B(n_281), .C(n_282), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_153), .A2(n_165), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_153), .A2(n_165), .B(n_515), .C(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_153), .A2(n_165), .B(n_533), .C(n_534), .Y(n_532) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx3_ASAP7_75t_L g164 ( .A(n_155), .Y(n_164) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_155), .Y(n_247) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
INVx5_ASAP7_75t_L g219 ( .A(n_162), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_162), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_162), .B(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g180 ( .A(n_164), .Y(n_180) );
INVx1_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_165), .A2(n_190), .B1(n_523), .B2(n_527), .Y(n_522) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_167), .Y(n_171) );
INVx4_ASAP7_75t_L g183 ( .A(n_167), .Y(n_183) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_167), .A2(n_531), .B(n_537), .Y(n_530) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g276 ( .A(n_168), .Y(n_276) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_169), .Y(n_267) );
AND2x2_ASAP7_75t_L g329 ( .A(n_169), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_169), .B(n_185), .Y(n_348) );
INVx1_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
OR2x2_ASAP7_75t_L g256 ( .A(n_170), .B(n_185), .Y(n_256) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_170), .Y(n_263) );
AND2x2_ASAP7_75t_L g315 ( .A(n_170), .B(n_201), .Y(n_315) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_170), .B(n_184), .C(n_298), .Y(n_340) );
AND2x2_ASAP7_75t_L g405 ( .A(n_170), .B(n_186), .Y(n_405) );
AND2x2_ASAP7_75t_L g439 ( .A(n_170), .B(n_185), .Y(n_439) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_181), .Y(n_170) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_171), .A2(n_202), .B(n_211), .Y(n_201) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_171), .A2(n_240), .B(n_248), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_178), .B(n_208), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g283 ( .A1(n_178), .A2(n_219), .B1(n_284), .B2(n_285), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_178), .B(n_497), .Y(n_496) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g195 ( .A(n_179), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g524 ( .A1(n_179), .A2(n_195), .B1(n_525), .B2(n_526), .Y(n_524) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_182), .A2(n_513), .B(n_519), .Y(n_512) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_183), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_183), .B(n_225), .Y(n_224) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_183), .A2(n_229), .B(n_236), .Y(n_228) );
NOR2xp33_ASAP7_75t_SL g477 ( .A(n_183), .B(n_478), .Y(n_477) );
INVxp67_ASAP7_75t_L g265 ( .A(n_184), .Y(n_265) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_200), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_185), .B(n_298), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_185), .B(n_329), .Y(n_337) );
AND2x2_ASAP7_75t_L g387 ( .A(n_185), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g415 ( .A(n_185), .Y(n_415) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g322 ( .A(n_186), .B(n_315), .Y(n_322) );
BUFx3_ASAP7_75t_L g354 ( .A(n_186), .Y(n_354) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_198), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_187), .B(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_187), .B(n_563), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_190), .A2(n_230), .B(n_231), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_190), .A2(n_503), .B(n_504), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_190), .A2(n_557), .B(n_558), .Y(n_556) );
O2A1O1Ixp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_197), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_194), .A2(n_197), .B(n_233), .C(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_197), .A2(n_474), .B(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_197), .A2(n_560), .B(n_561), .Y(n_559) );
INVx2_ASAP7_75t_L g330 ( .A(n_200), .Y(n_330) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_201), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_206), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g508 ( .A(n_209), .Y(n_508) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_212), .A2(n_390), .B1(n_392), .B2(n_393), .Y(n_389) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
AND2x2_ASAP7_75t_L g249 ( .A(n_213), .B(n_250), .Y(n_249) );
INVx3_ASAP7_75t_SL g260 ( .A(n_213), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_213), .B(n_293), .Y(n_325) );
OR2x2_ASAP7_75t_L g344 ( .A(n_213), .B(n_227), .Y(n_344) );
AND2x2_ASAP7_75t_L g349 ( .A(n_213), .B(n_301), .Y(n_349) );
AND2x2_ASAP7_75t_L g352 ( .A(n_213), .B(n_294), .Y(n_352) );
AND2x2_ASAP7_75t_L g364 ( .A(n_213), .B(n_239), .Y(n_364) );
AND2x2_ASAP7_75t_L g380 ( .A(n_213), .B(n_228), .Y(n_380) );
AND2x4_ASAP7_75t_L g383 ( .A(n_213), .B(n_251), .Y(n_383) );
OR2x2_ASAP7_75t_L g400 ( .A(n_213), .B(n_336), .Y(n_400) );
OR2x2_ASAP7_75t_L g431 ( .A(n_213), .B(n_273), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_213), .B(n_359), .Y(n_433) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .C(n_221), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_219), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_222), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g307 ( .A(n_226), .B(n_271), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_226), .B(n_294), .Y(n_426) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_239), .Y(n_226) );
AND2x2_ASAP7_75t_L g259 ( .A(n_227), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g293 ( .A(n_227), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_227), .B(n_273), .Y(n_301) );
AND2x2_ASAP7_75t_L g319 ( .A(n_227), .B(n_251), .Y(n_319) );
OR2x2_ASAP7_75t_L g336 ( .A(n_227), .B(n_294), .Y(n_336) );
INVx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
BUFx2_ASAP7_75t_L g252 ( .A(n_228), .Y(n_252) );
AND2x2_ASAP7_75t_L g359 ( .A(n_228), .B(n_239), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g288 ( .A(n_238), .Y(n_288) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_238), .A2(n_481), .B(n_488), .Y(n_480) );
INVx2_ASAP7_75t_L g251 ( .A(n_239), .Y(n_251) );
INVx1_ASAP7_75t_L g371 ( .A(n_239), .Y(n_371) );
AND2x2_ASAP7_75t_L g421 ( .A(n_239), .B(n_260), .Y(n_421) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_247), .Y(n_486) );
AND2x2_ASAP7_75t_L g270 ( .A(n_250), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g305 ( .A(n_250), .B(n_260), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_250), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_L g292 ( .A(n_251), .B(n_260), .Y(n_292) );
OR2x2_ASAP7_75t_L g408 ( .A(n_252), .B(n_382), .Y(n_408) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_255), .B(n_388), .Y(n_394) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OAI32xp33_ASAP7_75t_L g350 ( .A1(n_256), .A2(n_351), .A3(n_353), .B1(n_355), .B2(n_356), .Y(n_350) );
OR2x2_ASAP7_75t_L g367 ( .A(n_256), .B(n_309), .Y(n_367) );
OAI21xp33_ASAP7_75t_SL g392 ( .A1(n_256), .A2(n_266), .B(n_297), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B1(n_266), .B2(n_269), .Y(n_257) );
INVxp33_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_259), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_260), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_260), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g418 ( .A(n_260), .B(n_359), .Y(n_418) );
OR2x2_ASAP7_75t_L g442 ( .A(n_260), .B(n_336), .Y(n_442) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_261), .A2(n_324), .B(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g302 ( .A(n_263), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_263), .B(n_268), .Y(n_320) );
AND2x2_ASAP7_75t_L g342 ( .A(n_264), .B(n_315), .Y(n_342) );
INVx1_ASAP7_75t_L g355 ( .A(n_264), .Y(n_355) );
OR2x2_ASAP7_75t_L g360 ( .A(n_264), .B(n_294), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_267), .B(n_309), .Y(n_308) );
OAI22xp33_ASAP7_75t_L g290 ( .A1(n_268), .A2(n_291), .B1(n_296), .B2(n_300), .Y(n_290) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_271), .A2(n_333), .B1(n_340), .B2(n_341), .Y(n_339) );
AND2x2_ASAP7_75t_L g417 ( .A(n_271), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_273), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g436 ( .A(n_273), .B(n_319), .Y(n_436) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B(n_286), .Y(n_273) );
INVx1_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_274), .A2(n_556), .B(n_562), .Y(n_555) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AOI21xp5_ASAP7_75t_SL g470 ( .A1(n_275), .A2(n_471), .B(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_276), .A2(n_502), .B(n_509), .Y(n_501) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_276), .A2(n_522), .B(n_528), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_276), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_278), .A2(n_287), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_302), .B1(n_303), .B2(n_308), .C(n_310), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_292), .B(n_294), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_292), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g311 ( .A(n_293), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g398 ( .A1(n_293), .A2(n_399), .B(n_400), .C(n_401), .Y(n_398) );
AND2x2_ASAP7_75t_L g403 ( .A(n_293), .B(n_383), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_SL g441 ( .A1(n_293), .A2(n_382), .B(n_442), .C(n_443), .Y(n_441) );
BUFx3_ASAP7_75t_L g333 ( .A(n_294), .Y(n_333) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_297), .B(n_354), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_297), .A2(n_417), .B(n_419), .C(n_425), .Y(n_416) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVxp67_ASAP7_75t_L g377 ( .A(n_299), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_301), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AOI211xp5_ASAP7_75t_L g321 ( .A1(n_305), .A2(n_322), .B(n_323), .C(n_331), .Y(n_321) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g406 ( .A(n_309), .Y(n_406) );
OR2x2_ASAP7_75t_L g423 ( .A(n_309), .B(n_353), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_317), .B2(n_320), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g323 ( .A1(n_312), .A2(n_324), .B1(n_325), .B2(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
OR2x2_ASAP7_75t_L g410 ( .A(n_314), .B(n_354), .Y(n_410) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g365 ( .A(n_315), .B(n_355), .Y(n_365) );
INVx1_ASAP7_75t_L g373 ( .A(n_316), .Y(n_373) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_319), .B(n_333), .Y(n_381) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_329), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g438 ( .A(n_330), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_337), .Y(n_331) );
INVx1_ASAP7_75t_L g368 ( .A(n_332), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_333), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_333), .B(n_364), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_333), .B(n_359), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_333), .B(n_380), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g395 ( .A1(n_333), .A2(n_343), .B(n_383), .C(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_343), .B1(n_345), .B2(n_349), .C(n_350), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_347), .B(n_355), .Y(n_429) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_349), .A2(n_364), .B(n_366), .C(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_352), .B(n_359), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_353), .B(n_406), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g353 ( .A(n_354), .Y(n_353) );
INVxp33_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
AOI21xp33_ASAP7_75t_SL g369 ( .A1(n_358), .A2(n_370), .B(n_372), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_358), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_359), .B(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_366), .B2(n_368), .C(n_369), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_365), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
NAND5xp2_ASAP7_75t_L g374 ( .A(n_375), .B(n_402), .C(n_416), .D(n_427), .E(n_440), .Y(n_374) );
AOI211xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .B(n_385), .C(n_398), .Y(n_375) );
INVx2_ASAP7_75t_SL g422 ( .A(n_376), .Y(n_422) );
NAND4xp25_ASAP7_75t_SL g378 ( .A(n_379), .B(n_381), .C(n_382), .D(n_384), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI211xp5_ASAP7_75t_SL g385 ( .A1(n_384), .A2(n_386), .B(n_389), .C(n_395), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_387), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_387), .A2(n_428), .B1(n_430), .B2(n_432), .C(n_434), .Y(n_427) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI221xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_404), .B1(n_407), .B2(n_409), .C(n_411), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_410), .A2(n_433), .B1(n_435), .B2(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_448), .B(n_452), .C(n_748), .Y(n_451) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
XOR2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_463), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_463) );
AND2x2_ASAP7_75t_SL g464 ( .A(n_465), .B(n_712), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_605), .C(n_678), .Y(n_465) );
OAI211xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_499), .B(n_538), .C(n_589), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
AND2x2_ASAP7_75t_L g554 ( .A(n_469), .B(n_555), .Y(n_554) );
INVx3_ASAP7_75t_L g572 ( .A(n_469), .Y(n_572) );
INVx2_ASAP7_75t_L g587 ( .A(n_469), .Y(n_587) );
INVx1_ASAP7_75t_L g617 ( .A(n_469), .Y(n_617) );
AND2x2_ASAP7_75t_L g667 ( .A(n_469), .B(n_588), .Y(n_667) );
AOI32xp33_ASAP7_75t_L g694 ( .A1(n_469), .A2(n_622), .A3(n_695), .B1(n_697), .B2(n_698), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_469), .B(n_544), .Y(n_700) );
AND2x2_ASAP7_75t_L g727 ( .A(n_469), .B(n_570), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_469), .B(n_736), .Y(n_735) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_477), .Y(n_469) );
AND2x2_ASAP7_75t_L g616 ( .A(n_479), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g638 ( .A(n_479), .Y(n_638) );
AND2x2_ASAP7_75t_L g723 ( .A(n_479), .B(n_554), .Y(n_723) );
AND2x2_ASAP7_75t_L g726 ( .A(n_479), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_490), .Y(n_479) );
INVx2_ASAP7_75t_L g546 ( .A(n_480), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_480), .B(n_570), .Y(n_576) );
AND2x2_ASAP7_75t_L g586 ( .A(n_480), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g622 ( .A(n_480), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_487), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B(n_486), .Y(n_483) );
AND2x2_ASAP7_75t_L g564 ( .A(n_490), .B(n_546), .Y(n_564) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g547 ( .A(n_491), .Y(n_547) );
AND2x2_ASAP7_75t_L g588 ( .A(n_491), .B(n_570), .Y(n_588) );
AND2x2_ASAP7_75t_L g657 ( .A(n_491), .B(n_555), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
OR2x2_ASAP7_75t_L g552 ( .A(n_500), .B(n_521), .Y(n_552) );
INVx1_ASAP7_75t_L g630 ( .A(n_500), .Y(n_630) );
AND2x2_ASAP7_75t_L g644 ( .A(n_500), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_500), .B(n_520), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_500), .B(n_642), .Y(n_696) );
AND2x2_ASAP7_75t_L g704 ( .A(n_500), .B(n_705), .Y(n_704) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g542 ( .A(n_501), .Y(n_542) );
AND2x2_ASAP7_75t_L g611 ( .A(n_501), .B(n_521), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_510), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g738 ( .A(n_510), .Y(n_738) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_511), .B(n_582), .Y(n_604) );
OR2x2_ASAP7_75t_L g633 ( .A(n_511), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g665 ( .A(n_511), .B(n_645), .Y(n_665) );
INVx1_ASAP7_75t_SL g685 ( .A(n_511), .Y(n_685) );
AND2x2_ASAP7_75t_L g689 ( .A(n_511), .B(n_551), .Y(n_689) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_512), .B(n_520), .Y(n_543) );
AND2x2_ASAP7_75t_L g550 ( .A(n_512), .B(n_530), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_512), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g592 ( .A(n_512), .B(n_574), .Y(n_592) );
INVx1_ASAP7_75t_SL g599 ( .A(n_512), .Y(n_599) );
BUFx2_ASAP7_75t_L g610 ( .A(n_512), .Y(n_610) );
AND2x2_ASAP7_75t_L g626 ( .A(n_512), .B(n_542), .Y(n_626) );
AND2x2_ASAP7_75t_L g641 ( .A(n_512), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g705 ( .A(n_512), .B(n_521), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_520), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g629 ( .A(n_520), .B(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_520), .A2(n_647), .B1(n_650), .B2(n_653), .C(n_658), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_520), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
INVx3_ASAP7_75t_L g574 ( .A(n_521), .Y(n_574) );
BUFx2_ASAP7_75t_L g584 ( .A(n_530), .Y(n_584) );
AND2x2_ASAP7_75t_L g598 ( .A(n_530), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g615 ( .A(n_530), .Y(n_615) );
OR2x2_ASAP7_75t_L g634 ( .A(n_530), .B(n_574), .Y(n_634) );
INVx3_ASAP7_75t_L g642 ( .A(n_530), .Y(n_642) );
AND2x2_ASAP7_75t_L g645 ( .A(n_530), .B(n_574), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_544), .B1(n_548), .B2(n_553), .C(n_565), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_541), .B(n_614), .Y(n_739) );
OR2x2_ASAP7_75t_L g742 ( .A(n_541), .B(n_573), .Y(n_742) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
OAI221xp5_ASAP7_75t_SL g565 ( .A1(n_542), .A2(n_566), .B1(n_573), .B2(n_575), .C(n_578), .Y(n_565) );
AND2x2_ASAP7_75t_L g582 ( .A(n_542), .B(n_574), .Y(n_582) );
AND2x2_ASAP7_75t_L g590 ( .A(n_542), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_542), .B(n_598), .Y(n_597) );
NAND2x1_ASAP7_75t_L g640 ( .A(n_542), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g692 ( .A(n_542), .B(n_634), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_544), .A2(n_652), .B1(n_681), .B2(n_683), .Y(n_680) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI322xp5_ASAP7_75t_L g589 ( .A1(n_545), .A2(n_554), .A3(n_590), .B1(n_593), .B2(n_596), .C1(n_600), .C2(n_603), .Y(n_589) );
OR2x2_ASAP7_75t_L g601 ( .A(n_545), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_546), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g580 ( .A(n_546), .B(n_555), .Y(n_580) );
INVx1_ASAP7_75t_L g595 ( .A(n_546), .Y(n_595) );
AND2x2_ASAP7_75t_L g661 ( .A(n_546), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g571 ( .A(n_547), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g662 ( .A(n_547), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_547), .B(n_570), .Y(n_736) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_551), .B(n_685), .Y(n_684) );
INVx3_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g636 ( .A(n_552), .B(n_583), .Y(n_636) );
OR2x2_ASAP7_75t_L g733 ( .A(n_552), .B(n_584), .Y(n_733) );
INVx1_ASAP7_75t_L g714 ( .A(n_553), .Y(n_714) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_564), .Y(n_553) );
INVx4_ASAP7_75t_L g602 ( .A(n_554), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_554), .B(n_621), .Y(n_627) );
INVx2_ASAP7_75t_L g570 ( .A(n_555), .Y(n_570) );
INVx1_ASAP7_75t_L g652 ( .A(n_564), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_564), .B(n_624), .Y(n_693) );
AOI21xp33_ASAP7_75t_L g639 ( .A1(n_566), .A2(n_640), .B(n_643), .Y(n_639) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g624 ( .A(n_570), .Y(n_624) );
INVx1_ASAP7_75t_L g651 ( .A(n_570), .Y(n_651) );
INVx1_ASAP7_75t_L g577 ( .A(n_571), .Y(n_577) );
AND2x2_ASAP7_75t_L g579 ( .A(n_571), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g675 ( .A(n_572), .B(n_661), .Y(n_675) );
AND2x2_ASAP7_75t_L g697 ( .A(n_572), .B(n_657), .Y(n_697) );
BUFx2_ASAP7_75t_L g649 ( .A(n_574), .Y(n_649) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AOI32xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .A3(n_582), .B1(n_583), .B2(n_585), .Y(n_578) );
INVx1_ASAP7_75t_L g659 ( .A(n_579), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_579), .A2(n_707), .B1(n_708), .B2(n_710), .Y(n_706) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_582), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_582), .B(n_641), .Y(n_682) );
AND2x2_ASAP7_75t_L g729 ( .A(n_582), .B(n_614), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_583), .B(n_630), .Y(n_677) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g730 ( .A(n_585), .Y(n_730) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g655 ( .A(n_586), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_588), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g702 ( .A(n_588), .B(n_622), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_588), .B(n_617), .Y(n_709) );
INVx1_ASAP7_75t_SL g691 ( .A(n_590), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_591), .B(n_642), .Y(n_669) );
NOR4xp25_ASAP7_75t_L g715 ( .A(n_591), .B(n_614), .C(n_716), .D(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_592), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVxp67_ASAP7_75t_L g672 ( .A(n_595), .Y(n_672) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI21xp33_ASAP7_75t_L g722 ( .A1(n_598), .A2(n_689), .B(n_723), .Y(n_722) );
AND2x4_ASAP7_75t_L g614 ( .A(n_599), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g663 ( .A(n_602), .Y(n_663) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND4xp25_ASAP7_75t_SL g605 ( .A(n_606), .B(n_631), .C(n_646), .D(n_666), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_612), .B(n_616), .C(n_618), .Y(n_606) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g698 ( .A(n_611), .B(n_641), .Y(n_698) );
AND2x2_ASAP7_75t_L g707 ( .A(n_611), .B(n_685), .Y(n_707) );
INVx3_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_614), .B(n_649), .Y(n_711) );
AND2x2_ASAP7_75t_L g623 ( .A(n_617), .B(n_624), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_625), .B1(n_627), .B2(n_628), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
AND2x2_ASAP7_75t_L g721 ( .A(n_621), .B(n_667), .Y(n_721) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_623), .B(n_672), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_624), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_635), .B(n_637), .C(n_639), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_632), .A2(n_667), .B1(n_668), .B2(n_670), .C(n_673), .Y(n_666) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_640), .A2(n_725), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_641), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_649), .B(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g679 ( .A(n_651), .Y(n_679) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_654), .A2(n_674), .B1(n_676), .B2(n_677), .Y(n_673) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI21xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B(n_664), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_663), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_674), .A2(n_700), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g719 ( .A(n_676), .Y(n_719) );
OAI211xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B(n_686), .C(n_706), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_690), .C(n_699), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B(n_693), .C(n_694), .Y(n_690) );
INVx1_ASAP7_75t_L g718 ( .A(n_696), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g740 ( .A1(n_697), .A2(n_723), .B(n_741), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI21xp5_ASAP7_75t_SL g732 ( .A1(n_709), .A2(n_733), .B(n_734), .Y(n_732) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_724), .C(n_737), .Y(n_712) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_720), .C(n_722), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
CKINVDCx14_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
endmodule