module real_aes_8629_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g484 ( .A1(n_0), .A2(n_145), .B(n_485), .C(n_488), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_1), .B(n_480), .Y(n_489) );
INVx1_ASAP7_75t_L g434 ( .A(n_2), .Y(n_434) );
INVx1_ASAP7_75t_L g143 ( .A(n_3), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_4), .B(n_146), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_5), .A2(n_448), .B(n_524), .Y(n_523) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_6), .A2(n_153), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_7), .A2(n_35), .B1(n_133), .B2(n_181), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_8), .B(n_153), .Y(n_161) );
AND2x6_ASAP7_75t_L g148 ( .A(n_9), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_10), .A2(n_148), .B(n_453), .C(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_11), .A2(n_39), .B1(n_728), .B2(n_729), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_11), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_12), .B(n_36), .Y(n_435) );
INVx1_ASAP7_75t_L g124 ( .A(n_13), .Y(n_124) );
INVx1_ASAP7_75t_L g127 ( .A(n_14), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_15), .B(n_129), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_16), .B(n_146), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_17), .B(n_120), .Y(n_227) );
AO32x2_ASAP7_75t_L g197 ( .A1(n_18), .A2(n_119), .A3(n_153), .B1(n_172), .B2(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_19), .B(n_133), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_20), .B(n_120), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_21), .A2(n_55), .B1(n_133), .B2(n_181), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g183 ( .A1(n_22), .A2(n_81), .B1(n_129), .B2(n_133), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_23), .B(n_133), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_24), .A2(n_172), .B(n_453), .C(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_25), .A2(n_172), .B(n_453), .C(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_26), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_27), .B(n_174), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_28), .A2(n_448), .B(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_29), .B(n_174), .Y(n_215) );
INVx2_ASAP7_75t_L g131 ( .A(n_30), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_31), .A2(n_451), .B(n_455), .C(n_461), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_32), .B(n_133), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_33), .B(n_174), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_34), .B(n_192), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_37), .B(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_38), .Y(n_501) );
INVx1_ASAP7_75t_L g729 ( .A(n_39), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_40), .B(n_146), .Y(n_518) );
AOI222xp33_ASAP7_75t_L g101 ( .A1(n_41), .A2(n_102), .B1(n_736), .B2(n_745), .C1(n_759), .C2(n_763), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_41), .A2(n_750), .B1(n_752), .B2(n_753), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_41), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_42), .B(n_448), .Y(n_504) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_43), .A2(n_107), .B1(n_108), .B2(n_429), .Y(n_106) );
INVx1_ASAP7_75t_L g429 ( .A(n_43), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_43), .A2(n_45), .B1(n_429), .B2(n_751), .Y(n_750) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_44), .A2(n_451), .B(n_461), .C(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_45), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_46), .B(n_133), .Y(n_156) );
INVx1_ASAP7_75t_L g486 ( .A(n_47), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_48), .A2(n_89), .B1(n_181), .B2(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g517 ( .A(n_49), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_50), .B(n_133), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_51), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_52), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_53), .B(n_448), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_54), .B(n_141), .Y(n_160) );
AOI22xp33_ASAP7_75t_SL g225 ( .A1(n_56), .A2(n_61), .B1(n_129), .B2(n_133), .Y(n_225) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_57), .A2(n_104), .B1(n_726), .B2(n_727), .C1(n_730), .C2(n_734), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_58), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_59), .B(n_133), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_60), .B(n_133), .Y(n_189) );
INVx1_ASAP7_75t_L g149 ( .A(n_62), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_63), .B(n_448), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_64), .B(n_480), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_65), .A2(n_135), .B(n_141), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_66), .B(n_133), .Y(n_144) );
INVx1_ASAP7_75t_L g123 ( .A(n_67), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_68), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_69), .B(n_146), .Y(n_459) );
AO32x2_ASAP7_75t_L g178 ( .A1(n_70), .A2(n_153), .A3(n_172), .B1(n_179), .B2(n_184), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_71), .B(n_147), .Y(n_498) );
INVx1_ASAP7_75t_L g168 ( .A(n_72), .Y(n_168) );
INVx1_ASAP7_75t_L g210 ( .A(n_73), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g483 ( .A(n_74), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_75), .B(n_458), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_76), .A2(n_453), .B(n_461), .C(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_77), .B(n_129), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_78), .Y(n_525) );
INVx1_ASAP7_75t_L g740 ( .A(n_79), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_80), .B(n_457), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_82), .B(n_181), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_83), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_84), .B(n_129), .Y(n_214) );
INVx2_ASAP7_75t_L g121 ( .A(n_85), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_86), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_87), .B(n_171), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_88), .B(n_129), .Y(n_157) );
OR2x2_ASAP7_75t_L g432 ( .A(n_90), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g439 ( .A(n_90), .Y(n_439) );
OR2x2_ASAP7_75t_L g744 ( .A(n_90), .B(n_733), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_91), .A2(n_100), .B1(n_129), .B2(n_130), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_92), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g456 ( .A(n_93), .Y(n_456) );
INVxp67_ASAP7_75t_L g528 ( .A(n_94), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_95), .B(n_129), .Y(n_166) );
INVx1_ASAP7_75t_L g494 ( .A(n_96), .Y(n_494) );
INVx1_ASAP7_75t_L g552 ( .A(n_97), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_98), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g519 ( .A(n_99), .B(n_174), .Y(n_519) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22x1_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_430), .B1(n_436), .B2(n_440), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_106), .A2(n_430), .B1(n_438), .B2(n_735), .Y(n_734) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_107), .A2(n_108), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_395), .Y(n_108) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_299), .C(n_383), .Y(n_109) );
NAND4xp25_ASAP7_75t_L g110 ( .A(n_111), .B(n_242), .C(n_264), .D(n_280), .Y(n_110) );
AOI221xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_175), .B1(n_201), .B2(n_220), .C(n_228), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_151), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_114), .B(n_220), .Y(n_254) );
NAND4xp25_ASAP7_75t_L g294 ( .A(n_114), .B(n_282), .C(n_295), .D(n_297), .Y(n_294) );
INVxp67_ASAP7_75t_L g411 ( .A(n_114), .Y(n_411) );
INVx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g293 ( .A(n_115), .B(n_231), .Y(n_293) );
AND2x2_ASAP7_75t_L g317 ( .A(n_115), .B(n_151), .Y(n_317) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g284 ( .A(n_116), .B(n_219), .Y(n_284) );
AND2x2_ASAP7_75t_L g324 ( .A(n_116), .B(n_305), .Y(n_324) );
AND2x2_ASAP7_75t_L g341 ( .A(n_116), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_116), .B(n_152), .Y(n_365) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g218 ( .A(n_117), .B(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g236 ( .A(n_117), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g248 ( .A(n_117), .B(n_152), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_117), .B(n_162), .Y(n_270) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_125), .B(n_150), .Y(n_117) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_118), .A2(n_163), .B(n_173), .Y(n_162) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_119), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_120), .Y(n_153) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_121), .B(n_122), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_139), .B(n_148), .Y(n_125) );
O2A1O1Ixp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B(n_132), .C(n_135), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_128), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_128), .A2(n_507), .B(n_508), .Y(n_506) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g134 ( .A(n_131), .Y(n_134) );
INVx1_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
INVx3_ASAP7_75t_L g209 ( .A(n_133), .Y(n_209) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_133), .Y(n_554) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g181 ( .A(n_134), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
AND2x6_ASAP7_75t_L g453 ( .A(n_134), .B(n_454), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_135), .A2(n_552), .B(n_553), .C(n_554), .Y(n_551) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_136), .A2(n_213), .B(n_214), .Y(n_212) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g458 ( .A(n_137), .Y(n_458) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx3_ASAP7_75t_L g147 ( .A(n_138), .Y(n_147) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
INVx1_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
AND2x2_ASAP7_75t_L g449 ( .A(n_138), .B(n_142), .Y(n_449) );
INVx1_ASAP7_75t_L g454 ( .A(n_138), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_143), .B(n_144), .C(n_145), .Y(n_139) );
O2A1O1Ixp5_ASAP7_75t_L g167 ( .A1(n_140), .A2(n_168), .B(n_169), .C(n_170), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_140), .A2(n_472), .B(n_473), .Y(n_471) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_145), .A2(n_159), .B(n_160), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_145), .A2(n_171), .B1(n_199), .B2(n_200), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_145), .A2(n_171), .B1(n_224), .B2(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_146), .A2(n_156), .B(n_157), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_146), .A2(n_165), .B(n_166), .Y(n_164) );
O2A1O1Ixp5_ASAP7_75t_SL g208 ( .A1(n_146), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_146), .B(n_528), .Y(n_527) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_147), .A2(n_171), .B1(n_180), .B2(n_183), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g154 ( .A1(n_148), .A2(n_155), .B(n_158), .Y(n_154) );
BUFx3_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_148), .A2(n_188), .B(n_193), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_148), .A2(n_208), .B(n_212), .Y(n_207) );
AND2x4_ASAP7_75t_L g448 ( .A(n_148), .B(n_449), .Y(n_448) );
INVx4_ASAP7_75t_SL g462 ( .A(n_148), .Y(n_462) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_148), .B(n_449), .Y(n_495) );
AND2x2_ASAP7_75t_L g251 ( .A(n_151), .B(n_252), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_151), .A2(n_301), .B1(n_304), .B2(n_306), .C(n_310), .Y(n_300) );
AND2x2_ASAP7_75t_L g359 ( .A(n_151), .B(n_324), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_151), .B(n_341), .Y(n_393) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_162), .Y(n_151) );
INVx3_ASAP7_75t_L g219 ( .A(n_152), .Y(n_219) );
AND2x2_ASAP7_75t_L g268 ( .A(n_152), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g322 ( .A(n_152), .B(n_237), .Y(n_322) );
AND2x2_ASAP7_75t_L g380 ( .A(n_152), .B(n_381), .Y(n_380) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_161), .Y(n_152) );
INVx4_ASAP7_75t_L g222 ( .A(n_153), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_153), .A2(n_504), .B(n_505), .Y(n_503) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_153), .Y(n_522) );
AND2x2_ASAP7_75t_L g220 ( .A(n_162), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g237 ( .A(n_162), .Y(n_237) );
INVx1_ASAP7_75t_L g292 ( .A(n_162), .Y(n_292) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_162), .Y(n_298) );
AND2x2_ASAP7_75t_L g343 ( .A(n_162), .B(n_219), .Y(n_343) );
OR2x2_ASAP7_75t_L g382 ( .A(n_162), .B(n_221), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_172), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_170), .A2(n_194), .B(n_195), .Y(n_193) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g487 ( .A(n_171), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g241 ( .A(n_172), .B(n_222), .C(n_223), .Y(n_241) );
INVx2_ASAP7_75t_L g184 ( .A(n_174), .Y(n_184) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_174), .A2(n_187), .B(n_196), .Y(n_186) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_174), .A2(n_207), .B(n_215), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_174), .A2(n_447), .B(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g477 ( .A(n_174), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_174), .A2(n_514), .B(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_175), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_185), .Y(n_175) );
AND2x2_ASAP7_75t_L g378 ( .A(n_176), .B(n_375), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_176), .B(n_360), .Y(n_410) );
BUFx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g309 ( .A(n_177), .B(n_233), .Y(n_309) );
AND2x2_ASAP7_75t_L g358 ( .A(n_177), .B(n_204), .Y(n_358) );
INVx1_ASAP7_75t_L g404 ( .A(n_177), .Y(n_404) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_178), .Y(n_217) );
AND2x2_ASAP7_75t_L g259 ( .A(n_178), .B(n_233), .Y(n_259) );
INVx1_ASAP7_75t_L g276 ( .A(n_178), .Y(n_276) );
AND2x2_ASAP7_75t_L g282 ( .A(n_178), .B(n_197), .Y(n_282) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_182), .Y(n_460) );
INVx2_ASAP7_75t_L g488 ( .A(n_182), .Y(n_488) );
INVx1_ASAP7_75t_L g474 ( .A(n_184), .Y(n_474) );
AND2x2_ASAP7_75t_L g350 ( .A(n_185), .B(n_258), .Y(n_350) );
INVx2_ASAP7_75t_L g415 ( .A(n_185), .Y(n_415) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_197), .Y(n_185) );
AND2x2_ASAP7_75t_L g232 ( .A(n_186), .B(n_233), .Y(n_232) );
OR2x2_ASAP7_75t_L g245 ( .A(n_186), .B(n_205), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_186), .B(n_204), .Y(n_273) );
INVx1_ASAP7_75t_L g279 ( .A(n_186), .Y(n_279) );
INVx1_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_186), .Y(n_308) );
INVx2_ASAP7_75t_L g376 ( .A(n_186), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g233 ( .A(n_197), .Y(n_233) );
BUFx2_ASAP7_75t_L g330 ( .A(n_197), .Y(n_330) );
AND2x2_ASAP7_75t_L g375 ( .A(n_197), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_216), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_203), .B(n_312), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_203), .A2(n_374), .B(n_388), .Y(n_398) );
AND2x2_ASAP7_75t_L g423 ( .A(n_203), .B(n_309), .Y(n_423) );
BUFx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g345 ( .A(n_205), .Y(n_345) );
AND2x2_ASAP7_75t_L g374 ( .A(n_205), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_206), .Y(n_258) );
INVx2_ASAP7_75t_L g277 ( .A(n_206), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_206), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g231 ( .A(n_217), .Y(n_231) );
OR2x2_ASAP7_75t_L g244 ( .A(n_217), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g312 ( .A(n_217), .B(n_308), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_217), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g413 ( .A(n_217), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_217), .B(n_350), .Y(n_425) );
AND2x2_ASAP7_75t_L g304 ( .A(n_218), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g327 ( .A(n_218), .B(n_220), .Y(n_327) );
INVx2_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
AND2x2_ASAP7_75t_L g267 ( .A(n_219), .B(n_240), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_219), .B(n_292), .Y(n_348) );
AND2x2_ASAP7_75t_L g262 ( .A(n_220), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g409 ( .A(n_220), .Y(n_409) );
AND2x2_ASAP7_75t_L g421 ( .A(n_220), .B(n_284), .Y(n_421) );
AND2x2_ASAP7_75t_L g247 ( .A(n_221), .B(n_237), .Y(n_247) );
INVx1_ASAP7_75t_L g342 ( .A(n_221), .Y(n_342) );
AO21x1_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_226), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_222), .B(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g480 ( .A(n_222), .Y(n_480) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_222), .A2(n_493), .B(n_500), .Y(n_492) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_222), .A2(n_549), .B(n_556), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_222), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x4_ASAP7_75t_L g240 ( .A(n_227), .B(n_241), .Y(n_240) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_234), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_231), .B(n_278), .Y(n_287) );
OR2x2_ASAP7_75t_L g419 ( .A(n_231), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g336 ( .A(n_232), .B(n_277), .Y(n_336) );
AND2x2_ASAP7_75t_L g344 ( .A(n_232), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g403 ( .A(n_232), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g427 ( .A(n_232), .B(n_274), .Y(n_427) );
NOR2xp67_ASAP7_75t_L g385 ( .A(n_233), .B(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g414 ( .A(n_233), .B(n_277), .Y(n_414) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2x1p5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
AND2x2_ASAP7_75t_L g266 ( .A(n_236), .B(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_L g428 ( .A(n_236), .Y(n_428) );
NOR2x1_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx1_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
AND2x2_ASAP7_75t_L g314 ( .A(n_239), .B(n_247), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_239), .B(n_382), .Y(n_408) );
INVx2_ASAP7_75t_L g253 ( .A(n_240), .Y(n_253) );
INVx3_ASAP7_75t_L g305 ( .A(n_240), .Y(n_305) );
OR2x2_ASAP7_75t_L g333 ( .A(n_240), .B(n_334), .Y(n_333) );
AOI311xp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_246), .A3(n_248), .B(n_249), .C(n_260), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g280 ( .A1(n_243), .A2(n_281), .B(n_283), .C(n_285), .Y(n_280) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_SL g265 ( .A(n_245), .Y(n_265) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g283 ( .A(n_247), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_247), .B(n_263), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_247), .B(n_248), .Y(n_416) );
AND2x2_ASAP7_75t_L g338 ( .A(n_248), .B(n_252), .Y(n_338) );
AOI21xp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_254), .B(n_255), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g396 ( .A(n_252), .B(n_284), .Y(n_396) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_253), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g290 ( .A(n_253), .Y(n_290) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
AND2x2_ASAP7_75t_L g281 ( .A(n_257), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g326 ( .A(n_259), .Y(n_326) );
AND2x4_ASAP7_75t_L g388 ( .A(n_259), .B(n_357), .Y(n_388) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AOI222xp33_ASAP7_75t_L g339 ( .A1(n_262), .A2(n_328), .B1(n_340), .B2(n_344), .C1(n_346), .C2(n_350), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_266), .B(n_268), .C(n_271), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_265), .B(n_309), .Y(n_332) );
INVx1_ASAP7_75t_L g354 ( .A(n_267), .Y(n_354) );
INVx1_ASAP7_75t_L g288 ( .A(n_269), .Y(n_288) );
OR2x2_ASAP7_75t_L g353 ( .A(n_270), .B(n_354), .Y(n_353) );
OAI21xp33_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_274), .B(n_278), .Y(n_271) );
NAND3xp33_ASAP7_75t_L g289 ( .A(n_272), .B(n_290), .C(n_291), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_272), .A2(n_309), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
AND2x2_ASAP7_75t_SL g295 ( .A(n_277), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g386 ( .A(n_277), .Y(n_386) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_277), .Y(n_402) );
INVx2_ASAP7_75t_L g360 ( .A(n_278), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_282), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g334 ( .A(n_284), .Y(n_334) );
OAI221xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B1(n_289), .B2(n_293), .C(n_294), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_288), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g422 ( .A(n_288), .Y(n_422) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g303 ( .A(n_295), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_295), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g361 ( .A(n_295), .B(n_309), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_295), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g394 ( .A(n_295), .B(n_329), .Y(n_394) );
BUFx3_ASAP7_75t_L g357 ( .A(n_296), .Y(n_357) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND5xp2_ASAP7_75t_L g299 ( .A(n_300), .B(n_318), .C(n_339), .D(n_351), .E(n_366), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AOI32xp33_ASAP7_75t_L g391 ( .A1(n_303), .A2(n_330), .A3(n_346), .B1(n_392), .B2(n_394), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_305), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g315 ( .A(n_309), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_313), .B1(n_315), .B2(n_316), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_325), .B1(n_327), .B2(n_328), .C(n_331), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g390 ( .A(n_322), .B(n_341), .Y(n_390) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_327), .A2(n_388), .B1(n_406), .B2(n_411), .C(n_412), .Y(n_405) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx2_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B1(n_335), .B2(n_337), .Y(n_331) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g349 ( .A(n_341), .Y(n_349) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AOI222xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B1(n_359), .B2(n_360), .C1(n_361), .C2(n_362), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_360), .A2(n_407), .B1(n_409), .B2(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_372), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_377), .B(n_379), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g420 ( .A(n_375), .Y(n_420) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
A2O1A1Ixp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B(n_389), .C(n_391), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_399), .C(n_424), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_396), .Y(n_400) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_405), .C(n_417), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B(n_416), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g438 ( .A(n_433), .B(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g733 ( .A(n_433), .Y(n_733) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2x2_ASAP7_75t_L g732 ( .A(n_439), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g735 ( .A(n_440), .Y(n_735) );
OR3x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_640), .C(n_683), .Y(n_440) );
NAND5xp2_ASAP7_75t_L g441 ( .A(n_442), .B(n_567), .C(n_597), .D(n_614), .E(n_629), .Y(n_441) );
AOI221xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_490), .B1(n_530), .B2(n_536), .C(n_540), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_465), .Y(n_443) );
OR2x2_ASAP7_75t_L g545 ( .A(n_444), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g584 ( .A(n_444), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g602 ( .A(n_444), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_444), .B(n_538), .Y(n_619) );
OR2x2_ASAP7_75t_L g631 ( .A(n_444), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_444), .B(n_590), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_444), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_444), .B(n_568), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_444), .B(n_576), .Y(n_682) );
AND2x2_ASAP7_75t_L g714 ( .A(n_444), .B(n_478), .Y(n_714) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_444), .Y(n_722) );
INVx5_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_445), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g542 ( .A(n_445), .B(n_520), .Y(n_542) );
BUFx2_ASAP7_75t_L g564 ( .A(n_445), .Y(n_564) );
AND2x2_ASAP7_75t_L g593 ( .A(n_445), .B(n_466), .Y(n_593) );
AND2x2_ASAP7_75t_L g648 ( .A(n_445), .B(n_546), .Y(n_648) );
OR2x6_ASAP7_75t_L g445 ( .A(n_446), .B(n_463), .Y(n_445) );
BUFx2_ASAP7_75t_L g469 ( .A(n_448), .Y(n_469) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_452), .A2(n_462), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_452), .A2(n_462), .B(n_525), .C(n_526), .Y(n_524) );
INVx5_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B(n_459), .C(n_460), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_457), .A2(n_460), .B(n_517), .C(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_465), .B(n_602), .Y(n_611) );
OAI32xp33_ASAP7_75t_L g625 ( .A1(n_465), .A2(n_561), .A3(n_626), .B1(n_627), .B2(n_628), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_465), .B(n_627), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_465), .B(n_545), .Y(n_668) );
INVx1_ASAP7_75t_SL g697 ( .A(n_465), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g706 ( .A(n_465), .B(n_492), .C(n_648), .D(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_478), .Y(n_465) );
INVx5_ASAP7_75t_L g539 ( .A(n_466), .Y(n_539) );
AND2x2_ASAP7_75t_L g568 ( .A(n_466), .B(n_479), .Y(n_568) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_466), .Y(n_647) );
AND2x2_ASAP7_75t_L g717 ( .A(n_466), .B(n_664), .Y(n_717) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
AOI21xp5_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_470), .B(n_474), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AND2x4_ASAP7_75t_L g590 ( .A(n_478), .B(n_539), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_478), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g624 ( .A(n_478), .B(n_546), .Y(n_624) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g538 ( .A(n_479), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g576 ( .A(n_479), .B(n_548), .Y(n_576) );
AND2x2_ASAP7_75t_L g585 ( .A(n_479), .B(n_547), .Y(n_585) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_489), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
AOI222xp33_ASAP7_75t_L g653 ( .A1(n_490), .A2(n_654), .B1(n_656), .B2(n_658), .C1(n_661), .C2(n_662), .Y(n_653) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_509), .Y(n_490) );
AND2x2_ASAP7_75t_L g586 ( .A(n_491), .B(n_587), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_491), .B(n_564), .C(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_502), .Y(n_491) );
INVx5_ASAP7_75t_SL g535 ( .A(n_492), .Y(n_535) );
OAI322xp33_ASAP7_75t_L g540 ( .A1(n_492), .A2(n_541), .A3(n_543), .B1(n_544), .B2(n_558), .C1(n_561), .C2(n_563), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_492), .B(n_533), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_492), .B(n_521), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_496), .Y(n_493) );
INVx2_ASAP7_75t_L g533 ( .A(n_502), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_502), .B(n_511), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_509), .B(n_571), .Y(n_626) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g605 ( .A(n_510), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
OR2x2_ASAP7_75t_L g534 ( .A(n_511), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_511), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g573 ( .A(n_511), .B(n_521), .Y(n_573) );
AND2x2_ASAP7_75t_L g596 ( .A(n_511), .B(n_533), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_511), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g612 ( .A(n_511), .B(n_571), .Y(n_612) );
AND2x2_ASAP7_75t_L g620 ( .A(n_511), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_511), .B(n_580), .Y(n_670) );
INVx5_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g560 ( .A(n_512), .B(n_535), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_512), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g587 ( .A(n_512), .B(n_521), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_512), .B(n_634), .Y(n_675) );
OR2x2_ASAP7_75t_L g691 ( .A(n_512), .B(n_635), .Y(n_691) );
AND2x2_ASAP7_75t_SL g698 ( .A(n_512), .B(n_652), .Y(n_698) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_512), .Y(n_705) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .Y(n_512) );
AND2x2_ASAP7_75t_L g559 ( .A(n_520), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g609 ( .A(n_520), .B(n_533), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_520), .B(n_535), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_520), .B(n_571), .Y(n_693) );
INVx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_521), .B(n_535), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_521), .B(n_533), .Y(n_581) );
OR2x2_ASAP7_75t_L g635 ( .A(n_521), .B(n_533), .Y(n_635) );
AND2x2_ASAP7_75t_L g652 ( .A(n_521), .B(n_532), .Y(n_652) );
INVxp67_ASAP7_75t_L g674 ( .A(n_521), .Y(n_674) );
AND2x2_ASAP7_75t_L g701 ( .A(n_521), .B(n_571), .Y(n_701) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_521), .Y(n_708) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_529), .Y(n_521) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_532), .B(n_582), .Y(n_655) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g571 ( .A(n_533), .B(n_535), .Y(n_571) );
OR2x2_ASAP7_75t_L g638 ( .A(n_533), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g582 ( .A(n_534), .Y(n_582) );
OR2x2_ASAP7_75t_L g643 ( .A(n_534), .B(n_635), .Y(n_643) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g543 ( .A(n_538), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_538), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g544 ( .A(n_539), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_539), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_539), .B(n_546), .Y(n_578) );
INVx2_ASAP7_75t_L g623 ( .A(n_539), .Y(n_623) );
AND2x2_ASAP7_75t_L g636 ( .A(n_539), .B(n_576), .Y(n_636) );
AND2x2_ASAP7_75t_L g661 ( .A(n_539), .B(n_585), .Y(n_661) );
INVx1_ASAP7_75t_L g613 ( .A(n_544), .Y(n_613) );
INVx2_ASAP7_75t_SL g600 ( .A(n_545), .Y(n_600) );
INVx1_ASAP7_75t_L g603 ( .A(n_546), .Y(n_603) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_547), .Y(n_566) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g664 ( .A(n_548), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .Y(n_549) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g633 ( .A(n_560), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g639 ( .A(n_560), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_560), .A2(n_642), .B1(n_644), .B2(n_649), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_560), .B(n_652), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_561), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g595 ( .A(n_562), .Y(n_595) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
OR2x2_ASAP7_75t_L g577 ( .A(n_564), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_564), .B(n_568), .Y(n_628) );
AND2x2_ASAP7_75t_L g651 ( .A(n_564), .B(n_652), .Y(n_651) );
BUFx2_ASAP7_75t_L g627 ( .A(n_566), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B(n_574), .C(n_588), .Y(n_567) );
INVx1_ASAP7_75t_L g591 ( .A(n_568), .Y(n_591) );
OAI221xp5_ASAP7_75t_SL g699 ( .A1(n_568), .A2(n_700), .B1(n_702), .B2(n_703), .C(n_706), .Y(n_699) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g718 ( .A(n_571), .Y(n_718) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g667 ( .A(n_573), .B(n_606), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_577), .B(n_579), .C(n_583), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OAI32xp33_ASAP7_75t_L g692 ( .A1(n_581), .A2(n_582), .A3(n_645), .B1(n_682), .B2(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
AND2x2_ASAP7_75t_L g724 ( .A(n_584), .B(n_623), .Y(n_724) );
AND2x2_ASAP7_75t_L g671 ( .A(n_585), .B(n_623), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_585), .B(n_593), .Y(n_689) );
AOI31xp33_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_591), .A3(n_592), .B(n_594), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_590), .B(n_602), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_590), .B(n_600), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_590), .A2(n_620), .B1(n_710), .B2(n_713), .C(n_715), .Y(n_709) );
CKINVDCx16_ASAP7_75t_R g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g615 ( .A(n_595), .B(n_616), .Y(n_615) );
AOI222xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_604), .B1(n_607), .B2(n_610), .C1(n_612), .C2(n_613), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g680 ( .A(n_599), .Y(n_680) );
INVx1_ASAP7_75t_L g702 ( .A(n_602), .Y(n_702) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_605), .A2(n_716), .B1(n_718), .B2(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g621 ( .A(n_606), .Y(n_621) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .B1(n_620), .B2(n_622), .C(n_625), .Y(n_614) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g659 ( .A(n_617), .B(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g711 ( .A(n_617), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g686 ( .A(n_622), .Y(n_686) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g650 ( .A(n_623), .Y(n_650) );
INVx1_ASAP7_75t_L g632 ( .A(n_624), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_627), .B(n_714), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_633), .B1(n_636), .B2(n_637), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g723 ( .A(n_636), .Y(n_723) );
INVxp33_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_638), .B(n_682), .Y(n_681) );
OAI32xp33_ASAP7_75t_L g672 ( .A1(n_639), .A2(n_673), .A3(n_674), .B1(n_675), .B2(n_676), .Y(n_672) );
NAND4xp25_ASAP7_75t_L g640 ( .A(n_641), .B(n_653), .C(n_665), .D(n_677), .Y(n_640) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
NAND2xp33_ASAP7_75t_SL g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_648), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
CKINVDCx16_ASAP7_75t_R g658 ( .A(n_659), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_662), .A2(n_678), .B1(n_695), .B2(n_698), .C(n_699), .Y(n_694) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g713 ( .A(n_664), .B(n_714), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B1(n_669), .B2(n_671), .C(n_672), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_674), .B(n_705), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g683 ( .A(n_684), .B(n_694), .C(n_709), .D(n_720), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B(n_690), .C(n_692), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g725 ( .A(n_712), .Y(n_725) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_724), .B(n_725), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
CKINVDCx14_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx3_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
NAND2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_742), .Y(n_737) );
NOR2xp33_ASAP7_75t_SL g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_SL g762 ( .A(n_739), .Y(n_762) );
INVx1_ASAP7_75t_L g761 ( .A(n_741), .Y(n_761) );
OA21x2_ASAP7_75t_L g764 ( .A1(n_741), .A2(n_762), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g755 ( .A(n_744), .Y(n_755) );
BUFx2_ASAP7_75t_L g765 ( .A(n_744), .Y(n_765) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_754), .B(n_756), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_750), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g758 ( .A(n_755), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
endmodule