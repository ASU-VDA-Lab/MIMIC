module real_aes_3877_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_932;
wire n_235;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_961;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_962;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_960;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_610;
wire n_581;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_968;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_0), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g963 ( .A1(n_0), .A2(n_16), .B1(n_140), .B2(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g593 ( .A(n_1), .Y(n_593) );
INVx1_ASAP7_75t_L g320 ( .A(n_2), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_3), .A2(n_21), .B1(n_227), .B2(n_270), .Y(n_290) );
AOI22x1_ASAP7_75t_SL g128 ( .A1(n_4), .A2(n_53), .B1(n_129), .B2(n_130), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_4), .Y(n_130) );
INVx2_ASAP7_75t_L g177 ( .A(n_5), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_6), .B(n_606), .Y(n_704) );
INVx1_ASAP7_75t_SL g239 ( .A(n_7), .Y(n_239) );
INVxp67_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
INVx1_ASAP7_75t_L g138 ( .A(n_8), .Y(n_138) );
INVx1_ASAP7_75t_L g936 ( .A(n_8), .Y(n_936) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_9), .B(n_216), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_10), .A2(n_43), .B1(n_605), .B2(n_656), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_11), .A2(n_49), .B1(n_268), .B2(n_585), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_12), .A2(n_69), .B1(n_567), .B2(n_568), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_13), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_14), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g588 ( .A(n_15), .Y(n_588) );
INVx1_ASAP7_75t_L g964 ( .A(n_16), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_17), .A2(n_58), .B1(n_215), .B2(n_216), .Y(n_214) );
INVx1_ASAP7_75t_L g591 ( .A(n_18), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g101 ( .A1(n_19), .A2(n_102), .B1(n_119), .B2(n_127), .C(n_950), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_19), .A2(n_962), .B1(n_963), .B2(n_965), .Y(n_961) );
CKINVDCx14_ASAP7_75t_R g965 ( .A(n_19), .Y(n_965) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_20), .A2(n_73), .B(n_157), .Y(n_156) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_20), .A2(n_73), .B(n_157), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_22), .A2(n_71), .B1(n_567), .B2(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_23), .B(n_173), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_24), .A2(n_83), .B1(n_160), .B2(n_163), .Y(n_159) );
INVx2_ASAP7_75t_L g274 ( .A(n_25), .Y(n_274) );
INVx1_ASAP7_75t_L g584 ( .A(n_26), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_27), .B(n_952), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_28), .A2(n_32), .B1(n_199), .B2(n_238), .Y(n_291) );
BUFx8_ASAP7_75t_SL g105 ( .A(n_29), .Y(n_105) );
BUFx3_ASAP7_75t_L g125 ( .A(n_29), .Y(n_125) );
O2A1O1Ixp5_ASAP7_75t_L g267 ( .A1(n_30), .A2(n_197), .B(n_268), .C(n_269), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_31), .A2(n_66), .B1(n_170), .B2(n_172), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_33), .Y(n_201) );
AO22x1_ASAP7_75t_L g701 ( .A1(n_34), .A2(n_81), .B1(n_244), .B2(n_702), .Y(n_701) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_35), .Y(n_609) );
AND2x2_ASAP7_75t_L g619 ( .A(n_36), .B(n_585), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_37), .B(n_244), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_38), .A2(n_84), .B1(n_224), .B2(n_226), .Y(n_223) );
INVx1_ASAP7_75t_L g116 ( .A(n_39), .Y(n_116) );
INVx1_ASAP7_75t_L g263 ( .A(n_40), .Y(n_263) );
AOI22x1_ASAP7_75t_L g641 ( .A1(n_41), .A2(n_98), .B1(n_567), .B2(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_42), .B(n_644), .Y(n_657) );
AND2x2_ASAP7_75t_L g117 ( .A(n_44), .B(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_45), .B(n_259), .Y(n_315) );
INVx2_ASAP7_75t_L g271 ( .A(n_46), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_47), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_48), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g279 ( .A(n_50), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_51), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g243 ( .A(n_52), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_53), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_54), .B(n_238), .Y(n_673) );
INVx1_ASAP7_75t_L g193 ( .A(n_55), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_56), .B(n_265), .Y(n_612) );
INVx1_ASAP7_75t_L g157 ( .A(n_57), .Y(n_157) );
AND2x4_ASAP7_75t_L g151 ( .A(n_59), .B(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g188 ( .A(n_59), .B(n_152), .Y(n_188) );
INVx1_ASAP7_75t_L g248 ( .A(n_60), .Y(n_248) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_61), .Y(n_168) );
INVx2_ASAP7_75t_L g570 ( .A(n_62), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_63), .A2(n_76), .B1(n_605), .B2(n_642), .Y(n_652) );
CKINVDCx14_ASAP7_75t_R g707 ( .A(n_64), .Y(n_707) );
AND2x2_ASAP7_75t_L g625 ( .A(n_65), .B(n_244), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_67), .B(n_241), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_68), .B(n_313), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_70), .B(n_307), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_72), .B(n_572), .Y(n_629) );
CKINVDCx14_ASAP7_75t_R g646 ( .A(n_74), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_75), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_77), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_78), .B(n_606), .Y(n_671) );
OR2x6_ASAP7_75t_L g113 ( .A(n_79), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_80), .B(n_164), .Y(n_245) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
INVx1_ASAP7_75t_L g118 ( .A(n_85), .Y(n_118) );
INVx1_ASAP7_75t_L g162 ( .A(n_86), .Y(n_162) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_86), .Y(n_165) );
BUFx5_ASAP7_75t_L g200 ( .A(n_86), .Y(n_200) );
INVx2_ASAP7_75t_L g595 ( .A(n_87), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_88), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g282 ( .A(n_89), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_90), .Y(n_946) );
INVx1_ASAP7_75t_L g286 ( .A(n_91), .Y(n_286) );
NAND2xp33_ASAP7_75t_L g621 ( .A(n_92), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g207 ( .A(n_93), .Y(n_207) );
INVx2_ASAP7_75t_SL g152 ( .A(n_94), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_95), .B(n_190), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_96), .B(n_628), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_97), .B(n_307), .Y(n_306) );
AO32x2_ASAP7_75t_L g288 ( .A1(n_99), .A2(n_272), .A3(n_289), .B1(n_293), .B2(n_294), .Y(n_288) );
AO22x2_ASAP7_75t_L g325 ( .A1(n_99), .A2(n_289), .B1(n_326), .B2(n_328), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_100), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_106), .B(n_117), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx5_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_SL g121 ( .A(n_109), .Y(n_121) );
BUFx8_ASAP7_75t_SL g953 ( .A(n_109), .Y(n_953) );
BUFx12f_ASAP7_75t_L g957 ( .A(n_109), .Y(n_957) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OR2x6_ASAP7_75t_L g935 ( .A(n_112), .B(n_936), .Y(n_935) );
INVx8_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g137 ( .A(n_113), .B(n_138), .Y(n_137) );
OR2x6_ASAP7_75t_L g949 ( .A(n_113), .B(n_138), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_117), .Y(n_126) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
CKINVDCx6p67_ASAP7_75t_R g970 ( .A(n_125), .Y(n_970) );
OR2x2_ASAP7_75t_SL g968 ( .A(n_126), .B(n_969), .Y(n_968) );
OAI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_131), .B(n_937), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g937 ( .A1(n_128), .A2(n_938), .B(n_945), .Y(n_937) );
INVxp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVxp67_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_139), .B(n_553), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx8_ASAP7_75t_L g940 ( .A(n_137), .Y(n_940) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_139), .A2(n_939), .B(n_941), .Y(n_938) );
XNOR2x1_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AOI22xp5_ASAP7_75t_SL g959 ( .A1(n_141), .A2(n_960), .B1(n_961), .B2(n_966), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_141), .Y(n_960) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_477), .Y(n_141) );
NOR2xp67_ASAP7_75t_L g142 ( .A(n_143), .B(n_399), .Y(n_142) );
NAND3xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_341), .C(n_378), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_249), .B(n_295), .Y(n_144) );
OAI31xp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_179), .A3(n_210), .B(n_230), .Y(n_145) );
INVx1_ASAP7_75t_L g536 ( .A(n_146), .Y(n_536) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g373 ( .A(n_147), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g405 ( .A(n_147), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_147), .B(n_332), .Y(n_419) );
AND2x2_ASAP7_75t_L g523 ( .A(n_147), .B(n_509), .Y(n_523) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g397 ( .A(n_148), .B(n_353), .Y(n_397) );
AND2x2_ASAP7_75t_L g436 ( .A(n_148), .B(n_333), .Y(n_436) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_148), .Y(n_470) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g350 ( .A(n_149), .Y(n_350) );
INVx1_ASAP7_75t_L g369 ( .A(n_149), .Y(n_369) );
AOI21x1_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_158), .B(n_176), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx3_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_151), .Y(n_293) );
AND2x2_ASAP7_75t_L g326 ( .A(n_151), .B(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g565 ( .A(n_151), .Y(n_565) );
INVx1_ASAP7_75t_L g580 ( .A(n_151), .Y(n_580) );
AOI21xp33_ASAP7_75t_SL g632 ( .A1(n_153), .A2(n_564), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_154), .B(n_219), .Y(n_235) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g572 ( .A(n_155), .Y(n_572) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
BUFx3_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_166), .B1(n_169), .B2(n_174), .Y(n_158) );
INVx2_ASAP7_75t_L g702 ( .A(n_160), .Y(n_702) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g185 ( .A(n_161), .Y(n_185) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g171 ( .A(n_162), .Y(n_171) );
INVx1_ASAP7_75t_L g568 ( .A(n_163), .Y(n_568) );
INVx1_ASAP7_75t_L g656 ( .A(n_163), .Y(n_656) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
INVx2_ASAP7_75t_L g238 ( .A(n_164), .Y(n_238) );
INVx1_ASAP7_75t_L g311 ( .A(n_164), .Y(n_311) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx6_ASAP7_75t_L g173 ( .A(n_165), .Y(n_173) );
INVx2_ASAP7_75t_L g191 ( .A(n_165), .Y(n_191) );
INVx2_ASAP7_75t_L g227 ( .A(n_165), .Y(n_227) );
AOI21x1_ASAP7_75t_L g700 ( .A1(n_166), .A2(n_701), .B(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_167), .B(n_218), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_167), .A2(n_237), .B(n_239), .C(n_240), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_167), .A2(n_185), .B(n_282), .C(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g292 ( .A(n_167), .Y(n_292) );
INVxp67_ASAP7_75t_L g614 ( .A(n_167), .Y(n_614) );
INVx2_ASAP7_75t_SL g631 ( .A(n_167), .Y(n_631) );
INVx1_ASAP7_75t_L g675 ( .A(n_167), .Y(n_675) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx3_ASAP7_75t_L g175 ( .A(n_168), .Y(n_175) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_168), .Y(n_197) );
INVx1_ASAP7_75t_L g229 ( .A(n_168), .Y(n_229) );
INVx4_ASAP7_75t_L g260 ( .A(n_168), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_168), .B(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_168), .B(n_588), .Y(n_587) );
INVxp67_ASAP7_75t_L g623 ( .A(n_168), .Y(n_623) );
INVx3_ASAP7_75t_L g268 ( .A(n_170), .Y(n_268) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
INVx1_ASAP7_75t_L g278 ( .A(n_172), .Y(n_278) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
INVx2_ASAP7_75t_L g257 ( .A(n_173), .Y(n_257) );
INVx2_ASAP7_75t_SL g270 ( .A(n_173), .Y(n_270) );
INVx1_ASAP7_75t_L g622 ( .A(n_173), .Y(n_622) );
INVx1_ASAP7_75t_L g628 ( .A(n_173), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_174), .B(n_187), .Y(n_186) );
NOR3xp33_ASAP7_75t_L g192 ( .A(n_174), .B(n_187), .C(n_193), .Y(n_192) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_174), .B(n_563), .C(n_564), .Y(n_574) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_175), .A2(n_243), .B(n_244), .C(n_245), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_175), .A2(n_278), .B(n_279), .C(n_280), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
BUFx3_ASAP7_75t_L g272 ( .A(n_178), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_178), .B(n_274), .Y(n_273) );
INVx3_ASAP7_75t_L g307 ( .A(n_178), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_178), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g360 ( .A(n_179), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_179), .B(n_361), .Y(n_453) );
BUFx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OR2x2_ASAP7_75t_L g233 ( .A(n_180), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g338 ( .A(n_180), .Y(n_338) );
AND2x2_ASAP7_75t_L g471 ( .A(n_180), .B(n_374), .Y(n_471) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_204), .B(n_206), .Y(n_180) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_181), .A2(n_206), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_194), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B1(n_189), .B2(n_192), .Y(n_182) );
NOR2xp67_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_187), .B(n_196), .Y(n_195) );
AOI221x1_ASAP7_75t_L g254 ( .A1(n_187), .A2(n_255), .B1(n_258), .B2(n_262), .C(n_264), .Y(n_254) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g225 ( .A(n_191), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_198), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_196), .B(n_608), .Y(n_607) );
OAI22x1_ASAP7_75t_L g638 ( .A1(n_196), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_638) );
INVx4_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_197), .A2(n_290), .B1(n_291), .B2(n_292), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_197), .A2(n_310), .B(n_312), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_197), .A2(n_605), .B1(n_607), .B2(n_610), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_197), .B(n_651), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_197), .A2(n_670), .B(n_671), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g215 ( .A(n_200), .Y(n_215) );
INVx2_ASAP7_75t_L g244 ( .A(n_200), .Y(n_244) );
INVx2_ASAP7_75t_L g313 ( .A(n_200), .Y(n_313) );
INVx1_ASAP7_75t_L g317 ( .A(n_200), .Y(n_317) );
INVx2_ASAP7_75t_L g606 ( .A(n_200), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_202), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g585 ( .A(n_202), .Y(n_585) );
NOR2xp67_ASAP7_75t_SL g645 ( .A(n_204), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g706 ( .A(n_204), .B(n_707), .Y(n_706) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OA21x2_ASAP7_75t_L g602 ( .A1(n_205), .A2(n_603), .B(n_615), .Y(n_602) );
OA21x2_ASAP7_75t_L g693 ( .A1(n_205), .A2(n_603), .B(n_615), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx1_ASAP7_75t_L g294 ( .A(n_208), .Y(n_294) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp67_ASAP7_75t_L g218 ( .A(n_209), .B(n_219), .Y(n_218) );
BUFx3_ASAP7_75t_L g221 ( .A(n_209), .Y(n_221) );
INVx1_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_209), .B(n_219), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_209), .B(n_219), .Y(n_321) );
INVx1_ASAP7_75t_L g327 ( .A(n_209), .Y(n_327) );
INVx2_ASAP7_75t_L g563 ( .A(n_209), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_209), .B(n_219), .Y(n_651) );
BUFx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g501 ( .A(n_211), .B(n_412), .Y(n_501) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g232 ( .A(n_212), .Y(n_232) );
INVx2_ASAP7_75t_L g337 ( .A(n_212), .Y(n_337) );
AND2x2_ASAP7_75t_L g356 ( .A(n_212), .B(n_305), .Y(n_356) );
AND2x2_ASAP7_75t_L g361 ( .A(n_212), .B(n_362), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g212 ( .A(n_213), .B(n_222), .Y(n_212) );
AND2x2_ASAP7_75t_SL g300 ( .A(n_213), .B(n_222), .Y(n_300) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_217), .B(n_220), .Y(n_213) );
INVx2_ASAP7_75t_L g567 ( .A(n_215), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_218), .B(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_228), .Y(n_222) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVxp67_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
INVx1_ASAP7_75t_L g640 ( .A(n_229), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_229), .B(n_651), .Y(n_654) );
INVx2_ASAP7_75t_L g515 ( .A(n_230), .Y(n_515) );
OR2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
AND2x4_ASAP7_75t_L g440 ( .A(n_231), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g455 ( .A(n_232), .B(n_339), .Y(n_455) );
INVx2_ASAP7_75t_L g417 ( .A(n_233), .Y(n_417) );
INVx1_ASAP7_75t_L g322 ( .A(n_234), .Y(n_322) );
INVx2_ASAP7_75t_L g340 ( .A(n_234), .Y(n_340) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_234), .Y(n_355) );
INVx2_ASAP7_75t_L g374 ( .A(n_234), .Y(n_374) );
AND2x2_ASAP7_75t_L g388 ( .A(n_234), .B(n_301), .Y(n_388) );
INVx1_ASAP7_75t_L g413 ( .A(n_234), .Y(n_413) );
AO31x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .A3(n_242), .B(n_246), .Y(n_234) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_244), .A2(n_265), .B1(n_590), .B2(n_592), .Y(n_589) );
NOR2xp33_ASAP7_75t_SL g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_247), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g644 ( .A(n_247), .Y(n_644) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_251), .B(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_287), .Y(n_251) );
AND2x2_ASAP7_75t_L g344 ( .A(n_252), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g372 ( .A(n_252), .Y(n_372) );
INVx2_ASAP7_75t_L g430 ( .A(n_252), .Y(n_430) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_275), .Y(n_252) );
INVx2_ASAP7_75t_L g333 ( .A(n_253), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_253), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g404 ( .A(n_253), .B(n_350), .Y(n_404) );
INVx1_ASAP7_75t_L g445 ( .A(n_253), .Y(n_445) );
AND2x2_ASAP7_75t_L g509 ( .A(n_253), .B(n_353), .Y(n_509) );
AO31x2_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_266), .A3(n_272), .B(n_273), .Y(n_253) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
AND2x2_ASAP7_75t_L g262 ( .A(n_259), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_260), .B(n_320), .Y(n_319) );
NAND3xp33_ASAP7_75t_SL g562 ( .A(n_260), .B(n_563), .C(n_564), .Y(n_562) );
NOR2xp33_ASAP7_75t_SL g590 ( .A(n_260), .B(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_260), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_265), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g328 ( .A(n_272), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
INVx2_ASAP7_75t_L g353 ( .A(n_275), .Y(n_353) );
AND2x4_ASAP7_75t_L g365 ( .A(n_275), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g407 ( .A(n_275), .Y(n_407) );
AND2x4_ASAP7_75t_L g444 ( .A(n_275), .B(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AO31x2_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .A3(n_284), .B(n_285), .Y(n_276) );
INVx1_ASAP7_75t_L g420 ( .A(n_287), .Y(n_420) );
INVx2_ASAP7_75t_L g422 ( .A(n_287), .Y(n_422) );
AND2x4_ASAP7_75t_L g451 ( .A(n_287), .B(n_436), .Y(n_451) );
AND2x2_ASAP7_75t_L g517 ( .A(n_287), .B(n_518), .Y(n_517) );
BUFx8_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g366 ( .A(n_288), .Y(n_366) );
AND2x2_ASAP7_75t_L g381 ( .A(n_288), .B(n_382), .Y(n_381) );
OAI21x1_ASAP7_75t_L g603 ( .A1(n_293), .A2(n_604), .B(n_611), .Y(n_603) );
AO31x2_ASAP7_75t_L g637 ( .A1(n_293), .A2(n_638), .A3(n_643), .B(n_645), .Y(n_637) );
AO31x2_ASAP7_75t_L g681 ( .A1(n_293), .A2(n_638), .A3(n_643), .B(n_645), .Y(n_681) );
INVxp67_ASAP7_75t_L g302 ( .A(n_294), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_323), .B1(n_330), .B2(n_334), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_296), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI211xp5_ASAP7_75t_L g496 ( .A1(n_297), .A2(n_379), .B(n_497), .C(n_503), .Y(n_496) );
AND2x4_ASAP7_75t_L g297 ( .A(n_298), .B(n_303), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NOR2xp67_ASAP7_75t_SL g490 ( .A(n_299), .B(n_392), .Y(n_490) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g425 ( .A(n_300), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g432 ( .A(n_300), .B(n_426), .Y(n_432) );
INVx1_ASAP7_75t_L g538 ( .A(n_300), .Y(n_538) );
OR2x2_ASAP7_75t_L g377 ( .A(n_301), .B(n_362), .Y(n_377) );
AND2x2_ASAP7_75t_L g384 ( .A(n_301), .B(n_337), .Y(n_384) );
AND2x2_ASAP7_75t_L g502 ( .A(n_301), .B(n_304), .Y(n_502) );
AND2x2_ASAP7_75t_L g461 ( .A(n_303), .B(n_384), .Y(n_461) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_322), .Y(n_303) );
OR2x2_ASAP7_75t_L g392 ( .A(n_304), .B(n_338), .Y(n_392) );
INVx1_ASAP7_75t_L g486 ( .A(n_304), .Y(n_486) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g339 ( .A(n_305), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g362 ( .A(n_305), .Y(n_362) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_305), .Y(n_414) );
INVx1_ASAP7_75t_L g426 ( .A(n_305), .Y(n_426) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_307), .B(n_565), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_314), .B(n_321), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B(n_318), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_L g398 ( .A(n_322), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_322), .B(n_512), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_323), .A2(n_418), .B(n_551), .C(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_329), .Y(n_324) );
INVx1_ASAP7_75t_L g345 ( .A(n_325), .Y(n_345) );
AND2x4_ASAP7_75t_L g352 ( .A(n_325), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g408 ( .A(n_325), .Y(n_408) );
AND2x2_ASAP7_75t_L g526 ( .A(n_325), .B(n_350), .Y(n_526) );
INVx2_ASAP7_75t_SL g402 ( .A(n_329), .Y(n_402) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_331), .B(n_402), .Y(n_474) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g393 ( .A(n_332), .B(n_366), .Y(n_393) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g380 ( .A(n_333), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_333), .B(n_366), .Y(n_395) );
BUFx3_ASAP7_75t_L g493 ( .A(n_333), .Y(n_493) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_336), .A2(n_391), .B1(n_393), .B2(n_394), .Y(n_390) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_337), .Y(n_465) );
BUFx2_ASAP7_75t_L g512 ( .A(n_337), .Y(n_512) );
AND2x4_ASAP7_75t_L g449 ( .A(n_338), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g383 ( .A(n_339), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g450 ( .A(n_340), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_354), .B(n_357), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_344), .B(n_536), .Y(n_541) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
OAI21xp33_ASAP7_75t_SL g385 ( .A1(n_348), .A2(n_351), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g481 ( .A(n_348), .Y(n_481) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g518 ( .A(n_349), .Y(n_518) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_350), .Y(n_549) );
INVx4_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_352), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x2_ASAP7_75t_L g387 ( .A(n_356), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g468 ( .A(n_356), .Y(n_468) );
AND2x2_ASAP7_75t_L g516 ( .A(n_356), .B(n_471), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_363), .B1(n_370), .B2(n_375), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_360), .B(n_543), .Y(n_542) );
NAND2xp67_ASAP7_75t_L g416 ( .A(n_361), .B(n_417), .Y(n_416) );
BUFx3_ASAP7_75t_L g438 ( .A(n_361), .Y(n_438) );
AND2x2_ASAP7_75t_L g546 ( .A(n_361), .B(n_449), .Y(n_546) );
AND2x2_ASAP7_75t_L g552 ( .A(n_361), .B(n_388), .Y(n_552) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_365), .B(n_368), .Y(n_386) );
INVx2_ASAP7_75t_L g498 ( .A(n_365), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_366), .B(n_382), .Y(n_460) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_SL g433 ( .A(n_368), .Y(n_433) );
AND2x2_ASAP7_75t_L g534 ( .A(n_368), .B(n_444), .Y(n_534) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g382 ( .A(n_369), .Y(n_382) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NOR2xp67_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_374), .Y(n_476) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g521 ( .A(n_376), .B(n_501), .Y(n_521) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g441 ( .A(n_377), .Y(n_441) );
OR2x6_ASAP7_75t_L g475 ( .A(n_377), .B(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_377), .Y(n_495) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_383), .B1(n_385), .B2(n_387), .C(n_389), .Y(n_378) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g505 ( .A(n_381), .Y(n_505) );
AND2x4_ASAP7_75t_L g410 ( .A(n_384), .B(n_411), .Y(n_410) );
NOR3xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_396), .C(n_398), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g548 ( .A(n_395), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g492 ( .A(n_397), .B(n_493), .Y(n_492) );
NAND4xp25_ASAP7_75t_L g399 ( .A(n_400), .B(n_427), .C(n_443), .D(n_456), .Y(n_399) );
O2A1O1Ixp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_405), .B(n_409), .C(n_415), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g467 ( .A(n_402), .Y(n_467) );
OAI32xp33_ASAP7_75t_L g535 ( .A1(n_402), .A2(n_423), .A3(n_504), .B1(n_536), .B2(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g421 ( .A(n_404), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g530 ( .A(n_404), .Y(n_530) );
INVx1_ASAP7_75t_L g466 ( .A(n_406), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_406), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g551 ( .A(n_406), .B(n_493), .Y(n_551) );
AND2x4_ASAP7_75t_SL g406 ( .A(n_407), .B(n_408), .Y(n_406) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_412), .Y(n_424) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI32xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .A3(n_420), .B1(n_421), .B2(n_423), .Y(n_415) );
AND2x2_ASAP7_75t_L g431 ( .A(n_417), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g482 ( .A(n_421), .Y(n_482) );
AND2x2_ASAP7_75t_L g508 ( .A(n_422), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g543 ( .A(n_425), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_433), .B(n_434), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_430), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_430), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g448 ( .A(n_432), .B(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B1(n_439), .B2(n_442), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g473 ( .A(n_436), .B(n_459), .Y(n_473) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_442), .A2(n_498), .B(n_499), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .B1(n_451), .B2(n_452), .Y(n_443) );
INVx2_ASAP7_75t_L g506 ( .A(n_444), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_444), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g485 ( .A(n_449), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g511 ( .A(n_449), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AOI221xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_461), .B1(n_462), .B2(n_469), .C(n_472), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_464), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g494 ( .A(n_465), .B(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g533 ( .A(n_471), .Y(n_533) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_471), .B(n_538), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_475), .Y(n_472) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_513), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_487), .C(n_496), .Y(n_478) );
OAI21xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_482), .B(n_483), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVxp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_490), .A2(n_528), .B1(n_531), .B2(n_534), .C(n_535), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_507), .B(n_510), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g532 ( .A(n_512), .Y(n_532) );
NAND3xp33_ASAP7_75t_SL g513 ( .A(n_514), .B(n_527), .C(n_539), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .C(n_519), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_522), .B1(n_524), .B2(n_525), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NOR2x1p5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_542), .B(n_544), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B(n_550), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_932), .Y(n_553) );
INVx2_ASAP7_75t_L g944 ( .A(n_554), .Y(n_944) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_555), .B(n_806), .Y(n_554) );
NOR4xp75_ASAP7_75t_L g555 ( .A(n_556), .B(n_719), .C(n_737), .D(n_763), .Y(n_555) );
AO21x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_596), .B(n_687), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_559), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g727 ( .A(n_559), .B(n_697), .Y(n_727) );
INVx2_ASAP7_75t_L g789 ( .A(n_559), .Y(n_789) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_576), .Y(n_559) );
INVx1_ASAP7_75t_L g661 ( .A(n_560), .Y(n_661) );
INVx1_ASAP7_75t_L g686 ( .A(n_560), .Y(n_686) );
AND2x2_ASAP7_75t_L g709 ( .A(n_560), .B(n_577), .Y(n_709) );
INVx1_ASAP7_75t_L g740 ( .A(n_560), .Y(n_740) );
INVx2_ASAP7_75t_L g772 ( .A(n_560), .Y(n_772) );
NOR2x1_ASAP7_75t_L g814 ( .A(n_560), .B(n_815), .Y(n_814) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_560), .Y(n_829) );
AND2x2_ASAP7_75t_L g878 ( .A(n_560), .B(n_665), .Y(n_878) );
OR2x6_ASAP7_75t_L g560 ( .A(n_561), .B(n_573), .Y(n_560) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_566), .B(n_569), .Y(n_561) );
INVx1_ASAP7_75t_L g579 ( .A(n_563), .Y(n_579) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g616 ( .A(n_571), .Y(n_616) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g771 ( .A(n_576), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g776 ( .A(n_577), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g796 ( .A(n_577), .Y(n_796) );
INVx1_ASAP7_75t_L g815 ( .A(n_577), .Y(n_815) );
AND2x2_ASAP7_75t_L g877 ( .A(n_577), .B(n_742), .Y(n_877) );
INVxp67_ASAP7_75t_L g907 ( .A(n_577), .Y(n_907) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_594), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OR2x2_ASAP7_75t_L g699 ( .A(n_580), .B(n_616), .Y(n_699) );
NAND3xp33_ASAP7_75t_SL g581 ( .A(n_582), .B(n_586), .C(n_589), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_658), .B1(n_677), .B2(n_684), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_634), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g848 ( .A(n_600), .Y(n_848) );
OR2x2_ASAP7_75t_L g930 ( .A(n_600), .B(n_762), .Y(n_930) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g761 ( .A(n_601), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_617), .Y(n_601) );
AND2x2_ASAP7_75t_L g678 ( .A(n_602), .B(n_679), .Y(n_678) );
NAND2x1_ASAP7_75t_L g723 ( .A(n_602), .B(n_636), .Y(n_723) );
AND2x2_ASAP7_75t_L g858 ( .A(n_602), .B(n_648), .Y(n_858) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_613), .B(n_614), .Y(n_611) );
AND2x2_ASAP7_75t_L g688 ( .A(n_617), .B(n_681), .Y(n_688) );
AND2x4_ASAP7_75t_L g712 ( .A(n_617), .B(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g831 ( .A(n_617), .B(n_681), .Y(n_831) );
AO21x2_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_624), .B(n_632), .Y(n_617) );
AO21x2_ASAP7_75t_L g683 ( .A1(n_618), .A2(n_624), .B(n_632), .Y(n_683) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_623), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g642 ( .A(n_622), .Y(n_642) );
OAI21x1_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B(n_630), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_629), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g633 ( .A(n_629), .Y(n_633) );
AOI21x1_ASAP7_75t_L g703 ( .A1(n_631), .A2(n_704), .B(n_705), .Y(n_703) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_647), .Y(n_634) );
INVx2_ASAP7_75t_L g714 ( .A(n_635), .Y(n_714) );
INVx1_ASAP7_75t_L g746 ( .A(n_635), .Y(n_746) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g736 ( .A(n_636), .B(n_683), .Y(n_736) );
INVx1_ASAP7_75t_L g750 ( .A(n_636), .Y(n_750) );
AND2x2_ASAP7_75t_L g890 ( .A(n_636), .B(n_694), .Y(n_890) );
INVx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g762 ( .A(n_647), .Y(n_762) );
OR2x2_ASAP7_75t_L g874 ( .A(n_647), .B(n_723), .Y(n_874) );
INVx2_ASAP7_75t_L g882 ( .A(n_647), .Y(n_882) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g679 ( .A(n_649), .B(n_653), .Y(n_679) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
OA21x2_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B(n_657), .Y(n_653) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g797 ( .A(n_661), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g822 ( .A(n_663), .B(n_782), .Y(n_822) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g756 ( .A(n_664), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g697 ( .A(n_665), .B(n_698), .Y(n_697) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g718 ( .A(n_666), .Y(n_718) );
AND2x2_ASAP7_75t_L g741 ( .A(n_666), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g753 ( .A(n_666), .B(n_698), .Y(n_753) );
AND2x4_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OAI21x1_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B(n_676), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B(n_675), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
AND2x2_ASAP7_75t_L g778 ( .A(n_678), .B(n_722), .Y(n_778) );
INVx1_ASAP7_75t_L g891 ( .A(n_678), .Y(n_891) );
AND2x2_ASAP7_75t_L g923 ( .A(n_678), .B(n_750), .Y(n_923) );
INVx2_ASAP7_75t_L g694 ( .A(n_679), .Y(n_694) );
AND2x2_ASAP7_75t_L g733 ( .A(n_679), .B(n_692), .Y(n_733) );
INVx1_ASAP7_75t_L g783 ( .A(n_679), .Y(n_783) );
INVx1_ASAP7_75t_L g835 ( .A(n_679), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_679), .B(n_802), .Y(n_843) );
BUFx3_ASAP7_75t_L g730 ( .A(n_680), .Y(n_730) );
NOR2xp67_ASAP7_75t_L g850 ( .A(n_680), .B(n_732), .Y(n_850) );
AND2x4_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g760 ( .A(n_681), .Y(n_760) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_L g722 ( .A(n_683), .Y(n_722) );
INVx1_ASAP7_75t_L g802 ( .A(n_683), .Y(n_802) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g752 ( .A(n_685), .B(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g755 ( .A(n_685), .B(n_756), .Y(n_755) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_685), .Y(n_784) );
OR2x2_ASAP7_75t_L g911 ( .A(n_685), .B(n_788), .Y(n_911) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g774 ( .A(n_686), .B(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_686), .B(n_840), .Y(n_839) );
OAI32xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .A3(n_695), .B1(n_710), .B2(n_715), .Y(n_687) );
INVx2_ASAP7_75t_L g846 ( .A(n_688), .Y(n_846) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g873 ( .A(n_690), .Y(n_873) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g793 ( .A(n_691), .Y(n_793) );
OR2x2_ASAP7_75t_L g800 ( .A(n_691), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g885 ( .A(n_692), .Y(n_885) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g713 ( .A(n_693), .Y(n_713) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_693), .Y(n_841) );
INVx1_ASAP7_75t_L g735 ( .A(n_694), .Y(n_735) );
INVx2_ASAP7_75t_L g725 ( .A(n_695), .Y(n_725) );
OR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_708), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_L g813 ( .A(n_697), .B(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g900 ( .A(n_697), .B(n_771), .Y(n_900) );
INVx2_ASAP7_75t_SL g742 ( .A(n_698), .Y(n_742) );
OAI21x1_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B(n_706), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_699), .A2(n_700), .B(n_706), .Y(n_777) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g849 ( .A(n_709), .B(n_753), .Y(n_849) );
NAND2x1_ASAP7_75t_SL g871 ( .A(n_709), .B(n_741), .Y(n_871) );
AND2x2_ASAP7_75t_L g880 ( .A(n_709), .B(n_769), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_709), .B(n_922), .Y(n_921) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g924 ( .A(n_711), .B(n_782), .Y(n_924) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
AND2x4_ASAP7_75t_SL g749 ( .A(n_712), .B(n_750), .Y(n_749) );
BUFx3_ASAP7_75t_L g825 ( .A(n_712), .Y(n_825) );
INVxp67_ASAP7_75t_SL g818 ( .A(n_713), .Y(n_818) );
INVx1_ASAP7_75t_L g851 ( .A(n_715), .Y(n_851) );
AOI211xp5_ASAP7_75t_SL g838 ( .A1(n_716), .A2(n_750), .B(n_839), .C(n_841), .Y(n_838) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g795 ( .A(n_717), .B(n_796), .Y(n_795) );
OR2x2_ASAP7_75t_L g853 ( .A(n_717), .B(n_854), .Y(n_853) );
AND2x2_ASAP7_75t_L g920 ( .A(n_717), .B(n_771), .Y(n_920) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g804 ( .A(n_718), .B(n_740), .Y(n_804) );
OR2x2_ASAP7_75t_L g819 ( .A(n_718), .B(n_776), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_718), .B(n_907), .Y(n_906) );
OAI22xp5_ASAP7_75t_SL g719 ( .A1(n_720), .A2(n_724), .B1(n_726), .B2(n_728), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_722), .Y(n_817) );
AND3x2_ASAP7_75t_L g897 ( .A(n_722), .B(n_882), .C(n_885), .Y(n_897) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OA21x2_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B(n_734), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g916 ( .A(n_731), .Y(n_916) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g747 ( .A(n_733), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
BUFx3_ASAP7_75t_L g811 ( .A(n_736), .Y(n_811) );
AND2x2_ASAP7_75t_L g881 ( .A(n_736), .B(n_882), .Y(n_881) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_743), .B(n_751), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
AND2x2_ASAP7_75t_L g861 ( .A(n_741), .B(n_771), .Y(n_861) );
INVx2_ASAP7_75t_L g869 ( .A(n_741), .Y(n_869) );
INVx1_ASAP7_75t_L g757 ( .A(n_742), .Y(n_757) );
INVx1_ASAP7_75t_L g786 ( .A(n_742), .Y(n_786) );
INVxp67_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_745), .B(n_748), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_745), .A2(n_766), .B1(n_781), .B2(n_787), .Y(n_780) );
OR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
OR2x2_ASAP7_75t_L g856 ( .A(n_746), .B(n_857), .Y(n_856) );
INVx2_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g766 ( .A(n_749), .Y(n_766) );
OAI21xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .B(n_758), .Y(n_751) );
INVx2_ASAP7_75t_L g788 ( .A(n_753), .Y(n_788) );
AND2x2_ASAP7_75t_L g833 ( .A(n_753), .B(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_755), .A2(n_856), .B1(n_884), .B2(n_886), .Y(n_883) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_757), .Y(n_769) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_759), .B(n_793), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_759), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND3x1_ASAP7_75t_L g763 ( .A(n_764), .B(n_779), .C(n_790), .Y(n_763) );
AOI21x1_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_767), .B(n_773), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_768), .A2(n_853), .B1(n_930), .B2(n_931), .Y(n_929) );
OR2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_778), .Y(n_773) );
INVx1_ASAP7_75t_L g823 ( .A(n_775), .Y(n_823) );
AND2x2_ASAP7_75t_L g903 ( .A(n_775), .B(n_829), .Y(n_903) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g805 ( .A(n_776), .Y(n_805) );
BUFx2_ASAP7_75t_L g798 ( .A(n_777), .Y(n_798) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .C(n_785), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g837 ( .A(n_786), .B(n_796), .Y(n_837) );
OR2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVxp67_ASAP7_75t_L g827 ( .A(n_789), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_794), .B1(n_799), .B2(n_803), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND3xp33_ASAP7_75t_SL g845 ( .A(n_792), .B(n_846), .C(n_847), .Y(n_845) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
AND2x2_ASAP7_75t_L g905 ( .A(n_797), .B(n_906), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_797), .B(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g840 ( .A(n_798), .Y(n_840) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_801), .B(n_835), .Y(n_931) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_802), .A2(n_827), .B1(n_828), .B2(n_830), .Y(n_826) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
NAND2x2_ASAP7_75t_L g914 ( .A(n_804), .B(n_915), .Y(n_914) );
NOR2x1_ASAP7_75t_L g806 ( .A(n_807), .B(n_892), .Y(n_806) );
NAND4xp25_ASAP7_75t_L g807 ( .A(n_808), .B(n_844), .C(n_859), .D(n_879), .Y(n_807) );
NOR2xp67_ASAP7_75t_L g808 ( .A(n_809), .B(n_820), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_812), .B1(n_816), .B2(n_819), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AOI21xp33_ASAP7_75t_L g901 ( .A1(n_812), .A2(n_824), .B(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g854 ( .A(n_814), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
OAI211xp5_ASAP7_75t_SL g836 ( .A1(n_818), .A2(n_837), .B(n_838), .C(n_842), .Y(n_836) );
INVx1_ASAP7_75t_L g863 ( .A(n_818), .Y(n_863) );
AOI21xp33_ASAP7_75t_L g888 ( .A1(n_819), .A2(n_889), .B(n_891), .Y(n_888) );
OAI321xp33_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .A3(n_824), .B1(n_826), .B2(n_832), .C(n_836), .Y(n_820) );
INVx2_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
OR2x2_ASAP7_75t_L g886 ( .A(n_823), .B(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_825), .B(n_866), .Y(n_865) );
NOR2x1_ASAP7_75t_R g908 ( .A(n_825), .B(n_889), .Y(n_908) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AND2x2_ASAP7_75t_L g909 ( .A(n_830), .B(n_858), .Y(n_909) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
OR2x2_ASAP7_75t_L g884 ( .A(n_831), .B(n_885), .Y(n_884) );
INVx2_ASAP7_75t_L g896 ( .A(n_831), .Y(n_896) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g866 ( .A(n_835), .Y(n_866) );
INVxp67_ASAP7_75t_L g922 ( .A(n_840), .Y(n_922) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
AOI222xp33_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_849), .B1(n_850), .B2(n_851), .C1(n_852), .C2(n_855), .Y(n_844) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g913 ( .A(n_848), .Y(n_913) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
OR2x2_ASAP7_75t_L g868 ( .A(n_854), .B(n_869), .Y(n_868) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
AOI221x1_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_862), .B1(n_864), .B2(n_867), .C(n_870), .Y(n_859) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OAI22xp33_ASAP7_75t_SL g870 ( .A1(n_871), .A2(n_872), .B1(n_874), .B2(n_875), .Y(n_870) );
INVx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AND2x4_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
BUFx3_ASAP7_75t_L g915 ( .A(n_877), .Y(n_915) );
INVx2_ASAP7_75t_L g887 ( .A(n_878), .Y(n_887) );
AOI211xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B(n_883), .C(n_888), .Y(n_879) );
NAND2x1_ASAP7_75t_L g895 ( .A(n_882), .B(n_896), .Y(n_895) );
OAI22xp5_ASAP7_75t_SL g912 ( .A1(n_886), .A2(n_913), .B1(n_914), .B2(n_916), .Y(n_912) );
INVx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
NAND3xp33_ASAP7_75t_SL g892 ( .A(n_893), .B(n_904), .C(n_917), .Y(n_892) );
O2A1O1Ixp33_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_897), .B(n_898), .C(n_901), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_908), .B1(n_909), .B2(n_910), .C(n_912), .Y(n_904) );
HB1xp67_ASAP7_75t_L g928 ( .A(n_907), .Y(n_928) );
INVxp67_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_923), .B1(n_924), .B2(n_925), .C(n_929), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_919), .B(n_921), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
BUFx12f_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
CKINVDCx11_ASAP7_75t_R g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g942 ( .A(n_935), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_940), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .Y(n_941) );
INVx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
AOI21xp33_ASAP7_75t_SL g950 ( .A1(n_951), .A2(n_954), .B(n_967), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g952 ( .A(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_955), .B(n_958), .Y(n_954) );
INVx2_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVxp33_ASAP7_75t_SL g966 ( .A(n_961), .Y(n_966) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
BUFx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
endmodule