module fake_jpeg_25536_n_82 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_42),
.Y(n_44)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_22),
.B(n_26),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_43),
.B(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_1),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_32),
.B1(n_35),
.B2(n_34),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_46),
.B(n_53),
.Y(n_59)
);

NOR4xp25_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_18),
.C(n_27),
.D(n_25),
.Y(n_46)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_29),
.B1(n_12),
.B2(n_24),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_30),
.B1(n_10),
.B2(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_4),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_60),
.Y(n_71)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_2),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_3),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_66),
.B1(n_5),
.B2(n_6),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_66),
.B(n_65),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_74),
.B(n_71),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_59),
.B(n_8),
.C(n_9),
.D(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_70),
.Y(n_79)
);

AO21x2_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_68),
.B(n_72),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_57),
.C(n_5),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_20),
.Y(n_82)
);


endmodule