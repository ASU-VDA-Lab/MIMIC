module real_jpeg_27217_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_287, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_287;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_256;
wire n_274;
wire n_101;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_18),
.B1(n_19),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_SL g88 ( 
.A1(n_0),
.A2(n_24),
.B(n_26),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_0),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_0),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_0),
.B(n_25),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_0),
.A2(n_42),
.B(n_47),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_0),
.A2(n_8),
.B(n_65),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_0),
.B(n_41),
.Y(n_165)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_1),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_5),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_5),
.A2(n_20),
.B1(n_64),
.B2(n_65),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_5),
.A2(n_20),
.B1(n_42),
.B2(n_44),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_7),
.A2(n_42),
.B1(n_44),
.B2(n_53),
.Y(n_111)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_8),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_11),
.A2(n_18),
.B1(n_19),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_11),
.A2(n_29),
.B1(n_42),
.B2(n_44),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_11),
.A2(n_29),
.B1(n_64),
.B2(n_65),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_279),
.B(n_283),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_68),
.B(n_278),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_30),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_15),
.B(n_30),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_15),
.B(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_21),
.B1(n_25),
.B2(n_28),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_17),
.A2(n_33),
.B(n_34),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_19),
.A2(n_23),
.B(n_36),
.C(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_21),
.A2(n_25),
.B1(n_35),
.B2(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_21),
.B(n_25),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_27),
.B1(n_43),
.B2(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_26),
.A2(n_36),
.B(n_48),
.C(n_140),
.Y(n_139)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_28),
.B(n_282),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_31),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_31),
.B(n_276),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_37),
.CI(n_49),
.CON(n_31),
.SN(n_31)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_33),
.A2(n_34),
.B(n_52),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_35),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_36),
.A2(n_42),
.B(n_62),
.C(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_36),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_36),
.B(n_63),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_41),
.B1(n_45),
.B2(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_40),
.B(n_80),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_41),
.A2(n_55),
.B(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_44),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_81),
.Y(n_100)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.C(n_56),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_77),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_50),
.B(n_84),
.C(n_85),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_50),
.A2(n_83),
.B1(n_99),
.B2(n_124),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_50),
.B(n_124),
.C(n_218),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_50),
.A2(n_83),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_54),
.A2(n_56),
.B1(n_257),
.B2(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_54),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_56),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_56),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_67),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_59),
.A2(n_63),
.B1(n_104),
.B2(n_111),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_59),
.A2(n_63),
.B1(n_67),
.B2(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_63),
.A2(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_64),
.B(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_92),
.Y(n_91)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_275),
.B(n_277),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_249),
.A3(n_268),
.B1(n_273),
.B2(n_274),
.C(n_287),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_231),
.B(n_248),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_212),
.B(n_230),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_133),
.B(n_195),
.C(n_211),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_121),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_74),
.B(n_121),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_96),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_75),
.B(n_97),
.C(n_107),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_85),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_130),
.C(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_77),
.A2(n_84),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_77),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_77),
.B(n_237),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_82),
.B(n_100),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_89),
.A2(n_128),
.B1(n_164),
.B2(n_167),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_89),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_89),
.B(n_179),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_89),
.B(n_154),
.C(n_166),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_95),
.B(n_118),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_91),
.B(n_92),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_91),
.A2(n_95),
.B1(n_116),
.B2(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_106),
.B2(n_107),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.C(n_105),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_99),
.A2(n_108),
.B1(n_109),
.B2(n_124),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_100),
.Y(n_256)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_105),
.A2(n_125),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_105),
.A2(n_125),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_105),
.A2(n_125),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_105),
.B(n_255),
.C(n_257),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_105),
.B(n_262),
.C(n_267),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_108),
.A2(n_109),
.B1(n_161),
.B2(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_115),
.Y(n_205)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_124),
.C(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_109),
.B(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B(n_113),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_113),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.C(n_129),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_125),
.B(n_205),
.C(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_129),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_130),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_194),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_189),
.B(n_193),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_157),
.B(n_188),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_145),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_144),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_154),
.C(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_153),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_156),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_156),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_201),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_183),
.B(n_187),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_168),
.B(n_182),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_163),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_161),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_164),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_172),
.B(n_181),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_178),
.B(n_180),
.Y(n_172)
);

INVx5_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_209),
.B2(n_210),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_204),
.C(n_210),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_201),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_209),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_214),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_229),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_221),
.C(n_229),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_226),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_226),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_226),
.A2(n_240),
.B(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_233),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_246),
.B2(n_247),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_239),
.C(n_247),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_251),
.C(n_258),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_251),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_245),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_260),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_260),
.Y(n_274)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_259),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);


endmodule