module fake_jpeg_21451_n_212 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

OR2x4_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_22),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_35),
.B1(n_42),
.B2(n_45),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_31),
.B1(n_32),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_43),
.B1(n_44),
.B2(n_37),
.Y(n_82)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_41),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_30),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_0),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_28),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_25),
.C(n_1),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_22),
.B1(n_20),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_15),
.B1(n_29),
.B2(n_21),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_36),
.A3(n_41),
.B1(n_24),
.B2(n_25),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_23),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_23),
.B(n_28),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_23),
.B(n_1),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_34),
.B1(n_39),
.B2(n_27),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_67),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_46),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_84),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_76),
.B1(n_82),
.B2(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_16),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_78),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_111)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_92),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_35),
.B1(n_43),
.B2(n_15),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_16),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_121)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_87),
.Y(n_109)
);

OR2x2_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_28),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_95),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_21),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_27),
.B1(n_23),
.B2(n_18),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_68),
.Y(n_116)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_97),
.B1(n_2),
.B2(n_6),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_99),
.C(n_1),
.Y(n_101)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_44),
.A3(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_37),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_96),
.Y(n_110)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_36),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_47),
.C(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_99),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_83),
.C(n_98),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_120),
.B1(n_121),
.B2(n_89),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_7),
.B(n_8),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_92),
.Y(n_137)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_140),
.C(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_104),
.B(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_79),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_119),
.B1(n_102),
.B2(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_73),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_84),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_84),
.B(n_96),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_102),
.B(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_77),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_139),
.B1(n_117),
.B2(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

XOR2x2_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_93),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_142),
.B1(n_111),
.B2(n_102),
.C(n_103),
.Y(n_150)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_85),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_108),
.B1(n_107),
.B2(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_147),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_117),
.B1(n_114),
.B2(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_131),
.B1(n_138),
.B2(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_158),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_134),
.A2(n_90),
.B1(n_97),
.B2(n_94),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_159),
.B1(n_155),
.B2(n_144),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_128),
.B(n_140),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_167),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_169),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_159),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_173),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_157),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_185),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_170),
.B1(n_160),
.B2(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_177),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_146),
.C(n_126),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_144),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_184),
.B(n_164),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_171),
.B(n_164),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_155),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_194),
.B(n_158),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_170),
.B1(n_143),
.B2(n_172),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_149),
.B1(n_123),
.B2(n_148),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_174),
.B(n_152),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_183),
.A2(n_123),
.B1(n_162),
.B2(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_197),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_179),
.B1(n_182),
.B2(n_181),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_189),
.B1(n_127),
.B2(n_139),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_199),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_185),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_175),
.Y(n_200)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_192),
.B(n_187),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_197),
.B(n_196),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_204),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_207),
.B(n_203),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_200),
.B(n_123),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_209),
.B1(n_12),
.B2(n_10),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_202),
.C(n_12),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_11),
.B(n_131),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_211),
.Y(n_212)
);


endmodule