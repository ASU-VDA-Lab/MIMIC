module fake_jpeg_4558_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

OR2x2_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_17),
.B1(n_19),
.B2(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_44),
.B1(n_25),
.B2(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_53),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_59),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_17),
.B1(n_15),
.B2(n_19),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_73),
.B1(n_23),
.B2(n_52),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

NAND2x1_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_34),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_64),
.B(n_52),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_23),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_53),
.B1(n_20),
.B2(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_48),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_23),
.B1(n_24),
.B2(n_22),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_16),
.B(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_42),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_89),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_63),
.B(n_64),
.Y(n_97)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_74),
.B1(n_72),
.B2(n_30),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_61),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_41),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_95),
.B1(n_64),
.B2(n_58),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_41),
.B1(n_30),
.B2(n_28),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_35),
.B(n_55),
.C(n_29),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_76),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22x1_ASAP7_75t_L g95 ( 
.A1(n_63),
.A2(n_35),
.B1(n_30),
.B2(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_108),
.B(n_113),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_58),
.C(n_75),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_101),
.C(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_88),
.C(n_89),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_81),
.B1(n_66),
.B2(n_28),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_75),
.C(n_74),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_68),
.C(n_47),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_62),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_119),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_90),
.B1(n_92),
.B2(n_95),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_109),
.B1(n_110),
.B2(n_104),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_128),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_103),
.B1(n_99),
.B2(n_94),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_103),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_1),
.B(n_2),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_142),
.B1(n_119),
.B2(n_118),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_98),
.B1(n_107),
.B2(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_120),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_125),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_123),
.C(n_126),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_77),
.B1(n_4),
.B2(n_5),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_134),
.B(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_150),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_129),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_123),
.C(n_114),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_139),
.C(n_137),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_138),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_127),
.C(n_118),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_146),
.B(n_150),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_136),
.B(n_139),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_150),
.B1(n_143),
.B2(n_6),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_161),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_133),
.B1(n_128),
.B2(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_133),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_163),
.B(n_164),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_13),
.B(n_12),
.Y(n_164)
);

OAI31xp33_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_11),
.A3(n_5),
.B(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_11),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_156),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_171),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_172),
.B(n_161),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_157),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_170),
.A2(n_160),
.B1(n_8),
.B2(n_9),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_3),
.C(n_8),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_9),
.B(n_168),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_177),
.B(n_9),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_173),
.Y(n_180)
);


endmodule