module real_jpeg_29751_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_339, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_339;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_0),
.B(n_56),
.Y(n_117)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_0),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_1),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_95),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_1),
.A2(n_61),
.B1(n_62),
.B2(n_95),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_1),
.A2(n_56),
.B1(n_58),
.B2(n_95),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_37),
.B1(n_61),
.B2(n_62),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_37),
.B1(n_56),
.B2(n_58),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_4),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_97),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_4),
.A2(n_56),
.B1(n_58),
.B2(n_97),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_97),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_5),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_7),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_7),
.A2(n_56),
.B1(n_58),
.B2(n_105),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_105),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_105),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_8),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_112),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_112),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_8),
.A2(n_56),
.B1(n_58),
.B2(n_112),
.Y(n_205)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_10),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_102),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_10),
.A2(n_56),
.B1(n_58),
.B2(n_102),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_102),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_11),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_29),
.B(n_33),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_11),
.B(n_31),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_11),
.A2(n_61),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_61),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_11),
.B(n_75),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_11),
.A2(n_137),
.B1(n_139),
.B2(n_205),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_11),
.A2(n_32),
.B(n_220),
.Y(n_219)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_12),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_13),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_13),
.A2(n_27),
.B1(n_56),
.B2(n_58),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_13),
.A2(n_27),
.B1(n_61),
.B2(n_62),
.Y(n_269)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_15),
.A2(n_61),
.B1(n_62),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_16),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_17),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_17),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_49),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_22),
.B(n_43),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_24),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_26),
.A2(n_35),
.B(n_109),
.C(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_31),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_31),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_28),
.A2(n_31),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_28),
.A2(n_31),
.B1(n_146),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_28),
.A2(n_31),
.B1(n_165),
.B2(n_260),
.Y(n_259)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_32),
.A2(n_69),
.B(n_71),
.C(n_72),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_32),
.B(n_69),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g228 ( 
.A1(n_32),
.A2(n_62),
.A3(n_69),
.B1(n_221),
.B2(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_33),
.B(n_109),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_83),
.B(n_336),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_76),
.C(n_78),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_44),
.A2(n_45),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_65),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_46),
.B(n_319),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_48),
.A2(n_80),
.B1(n_82),
.B2(n_287),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_52),
.A2(n_310),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_52),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_52),
.A2(n_65),
.B1(n_313),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_64),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_53),
.A2(n_59),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_53),
.A2(n_59),
.B1(n_135),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_53),
.A2(n_59),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_53),
.A2(n_59),
.B1(n_179),
.B2(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_53),
.B(n_109),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_53),
.A2(n_59),
.B1(n_101),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_53),
.A2(n_59),
.B1(n_64),
.B2(n_269),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_54),
.A2(n_58),
.A3(n_61),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_55),
.B(n_56),
.Y(n_183)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_56),
.B(n_210),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_61),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_65),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_74),
.B2(n_75),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_66),
.A2(n_67),
.B1(n_75),
.B2(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_67),
.A2(n_75),
.B1(n_94),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_67),
.A2(n_75),
.B1(n_149),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_67),
.A2(n_75),
.B1(n_167),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_72),
.B(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_72),
.B1(n_93),
.B2(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_68),
.A2(n_72),
.B1(n_96),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_68),
.A2(n_72),
.B1(n_126),
.B2(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_68),
.A2(n_72),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_69),
.Y(n_230)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_76),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_80),
.A2(n_82),
.B1(n_111),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_80),
.A2(n_82),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_329),
.B(n_335),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_304),
.A3(n_323),
.B1(n_327),
.B2(n_328),
.C(n_339),
.Y(n_84)
);

AOI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_256),
.A3(n_293),
.B1(n_298),
.B2(n_303),
.C(n_340),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_151),
.C(n_169),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_130),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_88),
.B(n_130),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_113),
.C(n_122),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_89),
.B(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_107),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_98),
.B2(n_99),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_99),
.C(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_103),
.A2(n_106),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_103),
.A2(n_106),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_109),
.B(n_139),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_113),
.A2(n_122),
.B1(n_123),
.B2(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_113),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_116),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_117),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_129),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_124),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_127),
.B(n_129),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_128),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_142),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_141),
.C(n_142),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_139),
.B1(n_140),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_137),
.A2(n_139),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_137),
.A2(n_139),
.B1(n_198),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_137),
.A2(n_139),
.B1(n_193),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_137),
.A2(n_139),
.B(n_158),
.Y(n_271)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_147),
.C(n_150),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_152),
.A2(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_153),
.B(n_154),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_168),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_156),
.B(n_161),
.C(n_168),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_157),
.B(n_159),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_160),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_250),
.B(n_255),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_236),
.B(n_249),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_214),
.B(n_235),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_194),
.B(n_213),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_184),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_174),
.B(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_176),
.B1(n_180),
.B2(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_192),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_202),
.B(n_212),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_196),
.B(n_201),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_207),
.B(n_211),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_218),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_226),
.C(n_234),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_231),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_238),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_245),
.C(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_273),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_273),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_264),
.C(n_272),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_264),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_258),
.Y(n_337)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.CI(n_263),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_261),
.C(n_263),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_260),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_262),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_270),
.B2(n_271),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_271),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_270),
.A2(n_285),
.B(n_288),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_291),
.B2(n_292),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_282),
.C(n_292),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_280),
.B(n_281),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_280),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_279),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_306),
.C(n_315),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_306),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_282)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_299),
.B(n_302),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_295),
.B(n_296),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_316),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_316),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_314),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_308),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_310),
.C(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_321),
.C(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_309),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_325),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule