module fake_jpeg_19968_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_9),
.B(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_85),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_89),
.Y(n_91)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_52),
.B1(n_59),
.B2(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_100),
.B1(n_76),
.B2(n_69),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_82),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_81),
.C(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_76),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_77),
.B1(n_54),
.B2(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_104),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_69),
.B1(n_64),
.B2(n_61),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_112),
.B1(n_73),
.B2(n_78),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_111),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_100),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_93),
.B1(n_60),
.B2(n_101),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_82),
.B1(n_62),
.B2(n_56),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_62),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_0),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_64),
.B(n_68),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_120),
.B(n_22),
.Y(n_146)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_58),
.B(n_63),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_126),
.B1(n_129),
.B2(n_67),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_55),
.B1(n_101),
.B2(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_79),
.B1(n_75),
.B2(n_74),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_127),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_135),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_141),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_66),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_145),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_33),
.B1(n_50),
.B2(n_46),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_12),
.B1(n_15),
.B2(n_20),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_24),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_154),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_159),
.Y(n_163)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_139),
.B(n_141),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_160),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_143),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_143),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_161),
.C(n_162),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_163),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_156),
.B1(n_151),
.B2(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_168),
.B(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_158),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_25),
.B(n_34),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_38),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_174),
.A2(n_132),
.B(n_41),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_51),
.Y(n_177)
);


endmodule