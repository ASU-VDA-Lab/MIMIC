module real_jpeg_23659_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_0),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_0),
.A2(n_52),
.B1(n_56),
.B2(n_60),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_0),
.A2(n_37),
.B1(n_41),
.B2(n_60),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_60),
.Y(n_186)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_5),
.A2(n_26),
.B1(n_37),
.B2(n_41),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_7),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_32),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_7),
.A2(n_32),
.B1(n_52),
.B2(n_56),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_8),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_44),
.B1(n_52),
.B2(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_44),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_8),
.A2(n_55),
.B(n_67),
.C(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_8),
.A2(n_44),
.B1(n_59),
.B2(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_51),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_8),
.A2(n_56),
.B(n_75),
.C(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_8),
.B(n_25),
.C(n_40),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_8),
.B(n_131),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_8),
.B(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_8),
.B(n_42),
.Y(n_202)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_134),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_132),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_110),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_110),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_96),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_82),
.B2(n_83),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_21),
.B(n_33),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_29),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_22),
.A2(n_91),
.B(n_95),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_23),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_25),
.B(n_198),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_31),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_27),
.B(n_94),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_27),
.A2(n_92),
.B(n_94),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_27),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_28),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_30),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_30),
.B(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_45),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_34),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_43),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_35),
.B(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_35),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_36)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_37),
.A2(n_41),
.B1(n_75),
.B2(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_37),
.B(n_174),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_41),
.A2(n_44),
.B(n_77),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_42),
.B(n_154),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_43),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_44),
.A2(n_54),
.B(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_45),
.B(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_71),
.B1(n_72),
.B2(n_81),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_63),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_68),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_56),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_64),
.Y(n_100)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_121),
.Y(n_120)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_78),
.B(n_79),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_73),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_73),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_73),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_78),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_80),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_85),
.B(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_87),
.B(n_171),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_89),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_95),
.B(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_106),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_109),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_116),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_111),
.A2(n_112),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_115),
.Y(n_230)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_126),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_119),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_130),
.B(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_231),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_225),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_165),
.B(n_224),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_155),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_138),
.B(n_155),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_146),
.C(n_150),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_139),
.B(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_142),
.C(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_146),
.B(n_150),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_147),
.A2(n_149),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_147),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_149),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_158),
.B(n_159),
.C(n_160),
.Y(n_226)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_219),
.B(n_223),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_207),
.B(n_218),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_188),
.B(n_206),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_169),
.B(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_172),
.B1(n_173),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_182),
.B2(n_187),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_181),
.C(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_186),
.B(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_195),
.B(n_205),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_190),
.B(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_201),
.B(n_204),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);


endmodule