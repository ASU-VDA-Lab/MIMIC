module real_jpeg_6854_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_1),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_1),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_1),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_1),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_1),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_2),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_2),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_2),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_2),
.B(n_36),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_2),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_3),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_3),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_3),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_3),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_3),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_3),
.B(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_4),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_5),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_5),
.B(n_68),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_5),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_5),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_5),
.B(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_5),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_5),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_5),
.B(n_443),
.Y(n_442)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_7),
.Y(n_135)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_7),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_7),
.Y(n_255)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_7),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_8),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_8),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_8),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_8),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_8),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_8),
.B(n_426),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_10),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_10),
.B(n_129),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_10),
.B(n_327),
.Y(n_364)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_12),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_12),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_12),
.Y(n_327)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_13),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_13),
.Y(n_247)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_13),
.Y(n_428)
);

BUFx5_ASAP7_75t_L g443 ( 
.A(n_13),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_14),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_14),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_14),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_14),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_14),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_14),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_15),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_15),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_15),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_15),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_15),
.B(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_115),
.B(n_364),
.C(n_526),
.D(n_528),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_20),
.B(n_73),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_56),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_44),
.C(n_48),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_22),
.A2(n_23),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_43),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_26),
.A2(n_27),
.B1(n_65),
.B2(n_69),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_26),
.A2(n_27),
.B1(n_241),
.B2(n_248),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_26),
.B(n_60),
.C(n_65),
.Y(n_528)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_33),
.C(n_39),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_27),
.B(n_330),
.C(n_331),
.Y(n_329)
);

OR2x2_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_30),
.Y(n_232)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_31),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_31),
.Y(n_342)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_32),
.B(n_108),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_32),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_49),
.C(n_53),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_33),
.A2(n_34),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_34),
.B(n_161),
.C(n_166),
.Y(n_263)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_37),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_37),
.Y(n_289)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_38),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_38),
.Y(n_397)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_39),
.A2(n_43),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_39),
.B(n_349),
.C(n_353),
.Y(n_501)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_101),
.C(n_106),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_49),
.A2(n_114),
.B1(n_187),
.B2(n_198),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_49),
.B(n_188),
.C(n_194),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_49),
.A2(n_106),
.B1(n_107),
.B2(n_114),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_51),
.Y(n_225)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_51),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_51),
.Y(n_384)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_51),
.Y(n_401)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_52),
.Y(n_143)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_64),
.B2(n_70),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_59),
.A2(n_60),
.B1(n_493),
.B2(n_494),
.Y(n_492)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_86),
.C(n_90),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_65),
.A2(n_69),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_65),
.B(n_253),
.C(n_290),
.Y(n_361)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_68),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_71),
.B(n_527),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.C(n_95),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_79),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.C(n_92),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_81),
.B1(n_92),
.B2(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_86),
.A2(n_90),
.B1(n_257),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_86),
.Y(n_495)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_90),
.A2(n_250),
.B1(n_251),
.B2(n_257),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_90),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_90),
.B(n_144),
.C(n_253),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_92),
.A2(n_99),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_92),
.B(n_328),
.C(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_92),
.A2(n_99),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_94),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_95),
.B(n_522),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_112),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_96),
.A2(n_97),
.B1(n_504),
.B2(n_505),
.Y(n_503)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_99),
.B(n_361),
.C(n_364),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_100),
.B(n_112),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_101),
.B(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_106),
.A2(n_107),
.B1(n_144),
.B2(n_252),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_106),
.A2(n_107),
.B1(n_290),
.B2(n_317),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_139),
.C(n_144),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_107),
.B(n_290),
.C(n_340),
.Y(n_502)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_110),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_111),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_520),
.B(n_525),
.Y(n_115)
);

AOI21x1_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_486),
.B(n_517),
.Y(n_116)
);

AO21x2_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_334),
.B(n_366),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_298),
.B(n_333),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_272),
.B(n_297),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_120),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_234),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_121),
.B(n_234),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_185),
.C(n_219),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_122),
.B(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_157),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_123),
.B(n_158),
.C(n_169),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_138),
.C(n_147),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_124),
.B(n_293),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_124),
.Y(n_529)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_132),
.CI(n_136),
.CON(n_124),
.SN(n_124)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_125),
.B(n_132),
.C(n_136),
.Y(n_233)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_129),
.Y(n_418)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_130),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_138),
.A2(n_147),
.B1(n_148),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_138),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_139),
.B(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_144),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_154),
.Y(n_291)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_152),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_152),
.Y(n_437)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_161),
.A2(n_168),
.B1(n_204),
.B2(n_205),
.Y(n_402)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_171),
.B(n_172),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_170),
.B(n_178),
.C(n_180),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_176),
.B(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_181),
.B(n_386),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_181),
.B(n_400),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_181),
.B(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_185),
.B(n_219),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_199),
.C(n_201),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_186),
.A2(n_199),
.B1(n_200),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_186),
.Y(n_277)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_193),
.B1(n_194),
.B2(n_197),
.Y(n_187)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_193),
.A2(n_194),
.B1(n_306),
.B2(n_312),
.Y(n_305)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_194),
.B(n_307),
.C(n_308),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_201),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.C(n_215),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_202),
.A2(n_203),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_216),
.Y(n_474)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_214),
.Y(n_351)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_233),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_222),
.C(n_233),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_226),
.C(n_229),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_224),
.A2(n_349),
.B1(n_352),
.B2(n_353),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_224),
.Y(n_353)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_235),
.B(n_237),
.C(n_271),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_258),
.B1(n_270),
.B2(n_271),
.Y(n_236)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_249),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_239),
.B(n_240),
.C(n_249),
.Y(n_320)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_242),
.Y(n_330)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_246),
.Y(n_331)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_253),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_253),
.A2(n_256),
.B1(n_290),
.B2(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_253),
.A2(n_256),
.B1(n_394),
.B2(n_395),
.Y(n_412)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_256),
.B(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_259),
.B(n_261),
.C(n_262),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_265),
.B(n_267),
.C(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_295),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_273),
.B(n_295),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.C(n_292),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_274),
.A2(n_275),
.B1(n_479),
.B2(n_480),
.Y(n_478)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_278),
.B(n_292),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.C(n_291),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_279),
.B(n_466),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_281),
.B(n_291),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.C(n_290),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_282),
.A2(n_283),
.B1(n_287),
.B2(n_288),
.Y(n_391)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_290),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_290),
.A2(n_317),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_299),
.B(n_334),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_301),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_335),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_301),
.B(n_335),
.Y(n_485)
);

FAx1_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_319),
.CI(n_332),
.CON(n_301),
.SN(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_315),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_313),
.B2(n_314),
.Y(n_303)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_304),
.B(n_314),
.C(n_315),
.Y(n_356)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_311),
.Y(n_411)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_322),
.C(n_324),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_329),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_336),
.B(n_338),
.C(n_354),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_354),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_344),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_339),
.B(n_345),
.C(n_346),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

INVx6_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_349),
.Y(n_352)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_365),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_355),
.B(n_358),
.C(n_360),
.Y(n_513)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_357),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_364),
.Y(n_363)
);

OAI31xp33_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_482),
.A3(n_483),
.B(n_485),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_476),
.B(n_481),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_369),
.A2(n_461),
.B(n_475),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_413),
.B(n_460),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_403),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_371),
.B(n_403),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_392),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_389),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_373),
.B(n_389),
.C(n_392),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_380),
.C(n_385),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_374),
.A2(n_375),
.B1(n_380),
.B2(n_381),
.Y(n_405)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx8_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_385),
.B(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_398),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_393),
.B(n_470),
.C(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_402),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_406),
.C(n_412),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_404),
.B(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_406),
.A2(n_412),
.B1(n_452),
.B2(n_458),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_410),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_407),
.Y(n_450)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_412),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_454),
.B(n_459),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_439),
.B(n_453),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_423),
.B(n_438),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_434),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_434),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_429),
.B(n_433),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_429),
.Y(n_433)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_433),
.A2(n_441),
.B1(n_447),
.B2(n_448),
.Y(n_440)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_433),
.Y(n_447)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_449),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_449),
.Y(n_453)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_441),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_442),
.A2(n_444),
.B(n_447),
.Y(n_455)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_450),
.A2(n_451),
.B(n_452),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_455),
.B(n_456),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_463),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_464),
.A2(n_465),
.B1(n_467),
.B2(n_468),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_469),
.C(n_472),
.Y(n_477)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.Y(n_468)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_478),
.Y(n_481)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_479),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_514),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_487),
.A2(n_518),
.B(n_519),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_506),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_506),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_488),
.Y(n_531)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_497),
.CI(n_503),
.CON(n_488),
.SN(n_488)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_489),
.B(n_497),
.C(n_503),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.C(n_496),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_491),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_496),
.Y(n_508)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_501),
.C(n_502),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_498),
.A2(n_499),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_502),
.Y(n_512)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_504),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_510),
.C(n_513),
.Y(n_506)
);

FAx1_ASAP7_75t_SL g516 ( 
.A(n_507),
.B(n_510),
.CI(n_513),
.CON(n_516),
.SN(n_516)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_508),
.Y(n_509)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_516),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_516),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_524),
.Y(n_525)
);


endmodule