module fake_jpeg_23406_n_52 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_52);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_17;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_11),
.B1(n_30),
.B2(n_27),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_36),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_33),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_19),
.A2(n_20),
.B1(n_17),
.B2(n_22),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_SL g39 ( 
.A1(n_21),
.A2(n_27),
.B(n_28),
.C(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_42),
.B1(n_38),
.B2(n_39),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.C(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_40),
.C(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_48),
.Y(n_50)
);

AO21x1_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_39),
.B(n_25),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_26),
.B(n_32),
.Y(n_52)
);


endmodule