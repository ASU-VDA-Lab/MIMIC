module fake_jpeg_30237_n_302 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_302);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_25),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_8),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_20),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_62),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_24),
.B1(n_30),
.B2(n_37),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_75),
.A2(n_77),
.B1(n_98),
.B2(n_0),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_24),
.B1(n_30),
.B2(n_37),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_23),
.B1(n_42),
.B2(n_19),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_84),
.A2(n_45),
.B1(n_60),
.B2(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_37),
.B1(n_24),
.B2(n_30),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_105),
.B1(n_106),
.B2(n_33),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_38),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_97),
.Y(n_121)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_30),
.B1(n_37),
.B2(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_40),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_19),
.B1(n_23),
.B2(n_31),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_23),
.B1(n_21),
.B2(n_36),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_57),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_107),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_113),
.A2(n_123),
.B1(n_133),
.B2(n_134),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_36),
.B1(n_21),
.B2(n_35),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_122),
.B1(n_132),
.B2(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_26),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_119),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_131),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_35),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_42),
.B1(n_29),
.B2(n_27),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_43),
.B1(n_42),
.B2(n_29),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_99),
.A3(n_72),
.B1(n_76),
.B2(n_83),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_102),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_27),
.B1(n_8),
.B2(n_11),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_0),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_7),
.B1(n_16),
.B2(n_14),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_7),
.B1(n_16),
.B2(n_14),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_11),
.B1(n_16),
.B2(n_14),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_0),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_145),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_6),
.C(n_13),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_79),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_1),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_78),
.B(n_86),
.C(n_4),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_94),
.B(n_112),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_92),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_78),
.B(n_74),
.C(n_110),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_116),
.B(n_142),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_118),
.B(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_118),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_168),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_144),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_94),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_117),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_171),
.B(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_78),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_82),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_135),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_113),
.B1(n_116),
.B2(n_126),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_181),
.A2(n_186),
.B1(n_193),
.B2(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_182),
.B(n_198),
.Y(n_222)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_121),
.B(n_138),
.C(n_115),
.D(n_119),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_183),
.A2(n_174),
.B(n_176),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_197),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_132),
.B1(n_134),
.B2(n_125),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_140),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_195),
.C(n_166),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_139),
.C(n_82),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_192),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_117),
.A3(n_147),
.B1(n_136),
.B2(n_131),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_131),
.B1(n_145),
.B2(n_146),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_156),
.C(n_169),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_153),
.A2(n_145),
.B1(n_129),
.B2(n_135),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_144),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_92),
.B1(n_112),
.B2(n_96),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_203),
.B1(n_207),
.B2(n_150),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_161),
.B1(n_166),
.B2(n_154),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_175),
.A2(n_153),
.B1(n_155),
.B2(n_163),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_156),
.B(n_12),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_135),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_194),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_155),
.A2(n_102),
.B1(n_4),
.B2(n_17),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_225),
.B1(n_181),
.B2(n_197),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_207),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_230),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_220),
.C(n_221),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_224),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_151),
.C(n_149),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_151),
.C(n_149),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_161),
.B(n_170),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_164),
.B1(n_172),
.B2(n_152),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_226),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_152),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_229),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_196),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_228),
.A2(n_202),
.B1(n_203),
.B2(n_189),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_225),
.B1(n_230),
.B2(n_192),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_220),
.C(n_221),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_246),
.C(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_204),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_188),
.C(n_193),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_185),
.B(n_188),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_228),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_254),
.C(n_262),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_222),
.A3(n_211),
.B1(n_215),
.B2(n_216),
.C1(n_224),
.C2(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_251),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_237),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_243),
.A2(n_186),
.B1(n_211),
.B2(n_209),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_255),
.B1(n_236),
.B2(n_243),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_189),
.C(n_218),
.Y(n_254)
);

AOI321xp33_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_183),
.A3(n_226),
.B1(n_200),
.B2(n_196),
.C(n_208),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_258),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_240),
.Y(n_258)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_208),
.A3(n_200),
.B1(n_184),
.B2(n_179),
.C1(n_162),
.C2(n_172),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_242),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_178),
.C(n_184),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_238),
.B(n_235),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_231),
.B(n_178),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_272),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_268),
.B1(n_273),
.B2(n_162),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_247),
.B(n_232),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_257),
.B(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_245),
.C(n_232),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_249),
.C(n_239),
.Y(n_277)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_256),
.B1(n_260),
.B2(n_261),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_278),
.B(n_279),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_281),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_269),
.Y(n_288)
);

OAI31xp33_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_231),
.A3(n_177),
.B(n_179),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_162),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_R g281 ( 
.A(n_270),
.B(n_17),
.C(n_2),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_265),
.Y(n_289)
);

NAND4xp25_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_273),
.C(n_266),
.D(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_267),
.C(n_269),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_267),
.C(n_275),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_274),
.B(n_279),
.C(n_278),
.D(n_17),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.C(n_286),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_294),
.B(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_287),
.C(n_284),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_292),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_298),
.A2(n_293),
.B1(n_102),
.B2(n_3),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_299),
.B(n_1),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_1),
.Y(n_302)
);


endmodule