module fake_jpeg_29679_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_58),
.Y(n_61)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_71),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_76),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_21),
.B1(n_35),
.B2(n_28),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_96),
.B1(n_26),
.B2(n_1),
.Y(n_126)
);

OR2x4_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_22),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_39),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_31),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_20),
.B1(n_22),
.B2(n_15),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_84),
.B1(n_89),
.B2(n_91),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_25),
.B1(n_32),
.B2(n_31),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_110),
.C(n_26),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_40),
.A2(n_20),
.B1(n_15),
.B2(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_32),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_0),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_20),
.B1(n_15),
.B2(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_36),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_90),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_28),
.B1(n_35),
.B2(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_93),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_35),
.B1(n_28),
.B2(n_30),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_46),
.B1(n_37),
.B2(n_26),
.Y(n_123)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_36),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_100),
.C(n_106),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_34),
.B(n_30),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_34),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_102),
.Y(n_136)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_23),
.B1(n_33),
.B2(n_60),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_107),
.B1(n_109),
.B2(n_37),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_55),
.B(n_24),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_60),
.B1(n_48),
.B2(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_41),
.A2(n_37),
.B1(n_29),
.B2(n_9),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_37),
.Y(n_110)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_122),
.A2(n_128),
.B1(n_108),
.B2(n_78),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_132),
.B1(n_138),
.B2(n_14),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_63),
.A2(n_37),
.B1(n_26),
.B2(n_8),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_139),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_69),
.B1(n_87),
.B2(n_94),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_65),
.B(n_7),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_10),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_26),
.B1(n_6),
.B2(n_10),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_1),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_76),
.A2(n_6),
.B1(n_13),
.B2(n_10),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_68),
.A2(n_83),
.B1(n_110),
.B2(n_73),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_SL g143 ( 
.A(n_117),
.B(n_88),
.C(n_61),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_158),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_82),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_145),
.B(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_82),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_82),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_157),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_137),
.B(n_138),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_111),
.B(n_112),
.C(n_64),
.D(n_95),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_168),
.B1(n_112),
.B2(n_104),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_75),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_127),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_110),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_170),
.C(n_173),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_93),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_118),
.A2(n_94),
.B1(n_87),
.B2(n_69),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_95),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_139),
.B(n_72),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_135),
.B1(n_3),
.B2(n_4),
.Y(n_208)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_103),
.C(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_124),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_187),
.Y(n_216)
);

NAND2x1p5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_134),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_193),
.Y(n_230)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_132),
.B1(n_123),
.B2(n_108),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_190),
.A2(n_206),
.B1(n_152),
.B2(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_195),
.B1(n_201),
.B2(n_208),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_129),
.B1(n_98),
.B2(n_75),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_197),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_154),
.A2(n_141),
.B(n_125),
.C(n_64),
.D(n_72),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_125),
.B(n_141),
.C(n_86),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_174),
.B(n_153),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_130),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_157),
.C(n_172),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_104),
.B1(n_86),
.B2(n_115),
.Y(n_201)
);

NAND2x1_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_119),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_205),
.A2(n_193),
.B(n_202),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_175),
.A2(n_144),
.B1(n_147),
.B2(n_164),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_173),
.B(n_171),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_223),
.B(n_182),
.C(n_192),
.D(n_183),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_214),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_147),
.B(n_150),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_199),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_163),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_229),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_153),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_226),
.C(n_201),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_222),
.A2(n_228),
.B1(n_207),
.B2(n_204),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_167),
.B(n_165),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_195),
.C(n_180),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_162),
.B1(n_159),
.B2(n_150),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_177),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_152),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_184),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_231),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_234),
.Y(n_256)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_191),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_248),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_197),
.B1(n_194),
.B2(n_196),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_181),
.C(n_188),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_223),
.C(n_210),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_250),
.B1(n_211),
.B2(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_179),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_203),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_182),
.B1(n_178),
.B2(n_185),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_239),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_245),
.A2(n_230),
.B1(n_218),
.B2(n_224),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_230),
.B1(n_218),
.B2(n_224),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_214),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_259),
.B(n_234),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_230),
.C(n_215),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_247),
.C(n_249),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_228),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_211),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_250),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_276),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_243),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_269),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_233),
.Y(n_269)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_274),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_232),
.B1(n_241),
.B2(n_237),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_271),
.A2(n_262),
.B1(n_261),
.B2(n_260),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_238),
.B(n_242),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_256),
.B(n_257),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_275),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_240),
.C(n_248),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_244),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_277),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_239),
.C(n_229),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_278),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_198),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_265),
.Y(n_284)
);

NOR2x1_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_268),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_286),
.A2(n_268),
.B1(n_270),
.B2(n_219),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_213),
.B(n_151),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_289),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_278),
.B(n_276),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_266),
.B1(n_273),
.B2(n_275),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_286),
.B1(n_293),
.B2(n_279),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_295),
.C(n_280),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_283),
.B(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_296),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_213),
.C(n_3),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_1),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_279),
.B(n_4),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_281),
.B(n_287),
.C(n_280),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_5),
.B(n_299),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_295),
.B(n_291),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_303),
.B(n_304),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_306),
.A2(n_305),
.B(n_5),
.Y(n_308)
);

NOR3xp33_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_307),
.C(n_5),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_5),
.Y(n_310)
);


endmodule