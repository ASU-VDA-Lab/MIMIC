module fake_jpeg_7580_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_20),
.B(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_57),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_2),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_20),
.B(n_42),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_23),
.B1(n_22),
.B2(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_60),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_43),
.B1(n_39),
.B2(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_3),
.Y(n_79)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_68),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_85),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_16),
.C(n_21),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_45),
.C(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_79),
.B(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_21),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_78),
.Y(n_92)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_16),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_38),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_84),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_4),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_14),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_51),
.B1(n_48),
.B2(n_38),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_51),
.B1(n_48),
.B2(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_64),
.C(n_69),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_52),
.B(n_55),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_71),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_106),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_4),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_105),
.B(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_95),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_38),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_113),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_80),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_91),
.B1(n_96),
.B2(n_98),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_65),
.C(n_66),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_122),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_105),
.B(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_99),
.B(n_113),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_100),
.B(n_88),
.C(n_94),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_98),
.C(n_110),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_100),
.B1(n_77),
.B2(n_120),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_51),
.B1(n_86),
.B2(n_35),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_96),
.B1(n_83),
.B2(n_84),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_99),
.B1(n_117),
.B2(n_108),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_139),
.C(n_123),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_121),
.C(n_109),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_148),
.C(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_111),
.B(n_105),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_111),
.C(n_75),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_22),
.C(n_28),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_132),
.C(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_158),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_157),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_131),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_154),
.A2(n_127),
.B(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_162),
.B(n_6),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_127),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_165),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_127),
.C(n_129),
.Y(n_165)
);

AOI31xp67_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_6),
.A3(n_7),
.B(n_28),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_159),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_171),
.C(n_9),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_152),
.B1(n_156),
.B2(n_8),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_160),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_165),
.B(n_161),
.C(n_9),
.D(n_13),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_175),
.B1(n_171),
.B2(n_14),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_174),
.B1(n_15),
.B2(n_7),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_177),
.Y(n_179)
);


endmodule