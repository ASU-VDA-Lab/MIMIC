module real_jpeg_28149_n_18 (n_17, n_8, n_0, n_2, n_341, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_341;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_0),
.B(n_49),
.Y(n_89)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_2),
.A2(n_27),
.B1(n_49),
.B2(n_51),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_2),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_4),
.A2(n_44),
.B1(n_55),
.B2(n_56),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_4),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_5),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_115),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_115),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_5),
.A2(n_49),
.B1(n_51),
.B2(n_115),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_6),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_6),
.A2(n_29),
.B(n_33),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_119),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_6),
.B(n_31),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_6),
.A2(n_55),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_6),
.B(n_55),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_6),
.B(n_71),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_6),
.A2(n_88),
.B1(n_243),
.B2(n_247),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_6),
.A2(n_32),
.B(n_259),
.Y(n_258)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_8),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_109),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_109),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_8),
.A2(n_49),
.B1(n_51),
.B2(n_109),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_9),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_9),
.A2(n_46),
.B1(n_55),
.B2(n_56),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_46),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_10),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_104),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_104),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_10),
.A2(n_49),
.B1(n_51),
.B2(n_104),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_12),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_106),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_12),
.A2(n_49),
.B1(n_51),
.B2(n_106),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_12),
.A2(n_55),
.B1(n_56),
.B2(n_106),
.Y(n_263)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_15),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_15),
.A2(n_37),
.B1(n_49),
.B2(n_51),
.Y(n_128)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_17),
.A2(n_55),
.B1(n_56),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_17),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_99),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_99),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_17),
.A2(n_49),
.B1(n_51),
.B2(n_99),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_332),
.B(n_335),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_79),
.B(n_331),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_21),
.B(n_38),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_21),
.B(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_21),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_23),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_25),
.A2(n_35),
.B(n_119),
.C(n_120),
.Y(n_118)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_31),
.B1(n_42),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_28),
.A2(n_31),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_28),
.A2(n_31),
.B1(n_105),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_28),
.A2(n_31),
.B1(n_114),
.B2(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_28),
.A2(n_31),
.B(n_36),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_31),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_63),
.B(n_65),
.C(n_66),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_63),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g267 ( 
.A1(n_32),
.A2(n_56),
.A3(n_67),
.B1(n_260),
.B2(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_33),
.B(n_119),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_72),
.C(n_74),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_39),
.A2(n_40),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.C(n_60),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_41),
.B(n_316),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_43),
.A2(n_76),
.B1(n_78),
.B2(n_166),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_47),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_47),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_47),
.A2(n_60),
.B1(n_310),
.B2(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_53),
.B(n_59),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_53),
.B1(n_97),
.B2(n_100),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_48),
.A2(n_53),
.B1(n_100),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_48),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_48),
.A2(n_53),
.B1(n_59),
.B2(n_139),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_48),
.A2(n_53),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_48),
.A2(n_53),
.B1(n_217),
.B2(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_48),
.B(n_119),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_48),
.A2(n_53),
.B1(n_184),
.B2(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_49),
.B(n_52),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_49),
.B(n_249),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_51),
.A2(n_55),
.A3(n_58),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_54)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_55),
.B(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_60),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_61),
.A2(n_71),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_61),
.A2(n_71),
.B1(n_110),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_61),
.A2(n_71),
.B1(n_180),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_61),
.A2(n_69),
.B1(n_71),
.B2(n_308),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_66),
.B(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_62),
.A2(n_66),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_62),
.A2(n_66),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_62),
.A2(n_66),
.B1(n_124),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_62),
.A2(n_66),
.B1(n_192),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_67),
.Y(n_269)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_72),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_78),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_76),
.A2(n_78),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_324),
.B(n_330),
.Y(n_79)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_301),
.A3(n_320),
.B1(n_322),
.B2(n_323),
.C(n_340),
.Y(n_80)
);

AOI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_150),
.A3(n_172),
.B1(n_295),
.B2(n_300),
.C(n_341),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_83),
.A2(n_296),
.B(n_299),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_131),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_84),
.B(n_131),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_111),
.C(n_126),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_85),
.B(n_126),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_101),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_102),
.C(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_96),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_87),
.B(n_96),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_90),
.B1(n_92),
.B2(n_95),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_92),
.B1(n_95),
.B2(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_92),
.B(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_88),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_88),
.A2(n_94),
.B1(n_237),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_88),
.A2(n_231),
.B1(n_232),
.B2(n_271),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_89),
.A2(n_93),
.B1(n_122),
.B2(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_89),
.A2(n_93),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g232 ( 
.A(n_93),
.Y(n_232)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_94),
.B(n_119),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_98),
.A2(n_137),
.B1(n_140),
.B2(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_123),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_112),
.B(n_123),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_117),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_121),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_129),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_149),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_143),
.C(n_149),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_141),
.B2(n_142),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_137),
.A2(n_140),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_142),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_141),
.A2(n_164),
.B(n_167),
.Y(n_312)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_143),
.Y(n_338)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_146),
.CI(n_148),
.CON(n_143),
.SN(n_143)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_146),
.C(n_148),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_151),
.B(n_152),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_170),
.B2(n_171),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_155),
.B(n_161),
.C(n_171),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B(n_160),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_159),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_158),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_160),
.B(n_303),
.CI(n_312),
.CON(n_302),
.SN(n_302)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_161)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_170),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_202),
.C(n_207),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_196),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_174),
.B(n_196),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_187),
.C(n_188),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_175),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_185),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_182),
.C(n_185),
.Y(n_199)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_187),
.Y(n_293)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_190),
.B(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_193),
.B(n_195),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_194),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_203),
.A2(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_204),
.B(n_205),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_289),
.B(n_294),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_275),
.B(n_288),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_253),
.B(n_274),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_233),
.B(n_252),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_222),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_212),
.B(n_222),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_218),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_214),
.B1(n_218),
.B2(n_219),
.Y(n_239)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_227),
.C(n_229),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_230),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_240),
.B(n_251),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_239),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_245),
.B(n_250),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_254),
.B(n_255),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_266),
.B1(n_272),
.B2(n_273),
.Y(n_255)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_261),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_265),
.C(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_277),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_284),
.C(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_313),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_302),
.B(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_313),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_306),
.B2(n_311),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_305),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_307),
.C(n_310),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_318),
.C(n_319),
.Y(n_325)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.Y(n_313)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_336),
.Y(n_335)
);


endmodule