module fake_jpeg_19938_n_66 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_66);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_66;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx11_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_22),
.Y(n_25)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_15),
.B1(n_18),
.B2(n_8),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_21),
.B(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_17),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_16),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_14),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

OR2x4_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_39),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_13),
.B1(n_10),
.B2(n_16),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_13),
.B1(n_18),
.B2(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_52),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_23),
.C(n_34),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_40),
.C(n_23),
.Y(n_55)
);

XOR2x2_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_41),
.B2(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_53),
.C(n_55),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_53),
.B(n_56),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_51),
.C(n_41),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_62),
.B1(n_4),
.B2(n_7),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_3),
.Y(n_66)
);


endmodule