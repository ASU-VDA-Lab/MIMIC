module fake_ariane_1385_n_219 (n_8, n_24, n_7, n_22, n_43, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_219);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_219;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_179;
wire n_64;
wire n_180;
wire n_160;
wire n_124;
wire n_119;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_205;
wire n_71;
wire n_109;
wire n_208;
wire n_96;
wire n_156;
wire n_209;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_200;
wire n_51;
wire n_166;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_217;
wire n_44;
wire n_82;
wire n_178;
wire n_57;
wire n_131;
wire n_201;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_214;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_188;
wire n_185;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_198;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_206;
wire n_207;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_211;
wire n_194;
wire n_97;
wire n_154;
wire n_215;
wire n_142;
wire n_161;
wire n_163;
wire n_186;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_63;
wire n_59;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_54;

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVxp33_ASAP7_75t_SL g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g58 ( 
.A(n_11),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

INVxp67_ASAP7_75t_SL g64 ( 
.A(n_7),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_0),
.Y(n_67)
);

INVxp33_ASAP7_75t_SL g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_31),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_22),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_1),
.B(n_2),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_1),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_2),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_3),
.B(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_60),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_5),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_53),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_62),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_53),
.B1(n_68),
.B2(n_65),
.Y(n_104)
);

OR2x6_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_70),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_61),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_74),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_85),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_113),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AO221x1_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_78),
.B1(n_90),
.B2(n_89),
.C(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

OR2x6_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_83),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NAND2x1p5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_89),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_104),
.C(n_101),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_106),
.Y(n_136)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_102),
.B(n_98),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_127),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

OAI21x1_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_111),
.B(n_107),
.Y(n_140)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_90),
.B(n_80),
.C(n_78),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_80),
.B(n_58),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_86),
.B(n_76),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_121),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_73),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_128),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

OAI21x1_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_115),
.B(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_136),
.B1(n_135),
.B2(n_138),
.Y(n_155)
);

OAI21x1_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_120),
.B(n_130),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_124),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_76),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_94),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_142),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_158),
.B1(n_154),
.B2(n_161),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_141),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_150),
.B1(n_159),
.B2(n_151),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_157),
.Y(n_175)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_148),
.B(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_6),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_6),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_179),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_172),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_176),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_181),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_165),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_88),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_163),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_160),
.B(n_163),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_144),
.B1(n_137),
.B2(n_73),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

OAI31xp33_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_199),
.A3(n_195),
.B(n_196),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_204),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_193),
.B1(n_198),
.B2(n_200),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_193),
.Y(n_209)
);

NAND4xp25_ASAP7_75t_SL g210 ( 
.A(n_208),
.B(n_8),
.C(n_9),
.D(n_12),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_25),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_210),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_27),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_213),
.A2(n_33),
.B(n_35),
.Y(n_216)
);

NAND2x1_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_43),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_216),
.B(n_214),
.Y(n_219)
);


endmodule