module fake_jpeg_11708_n_165 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx8_ASAP7_75t_SL g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_6),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_74),
.Y(n_80)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_18),
.B1(n_43),
.B2(n_40),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_66),
.B1(n_59),
.B2(n_63),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_73),
.A2(n_50),
.B1(n_67),
.B2(n_52),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_0),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_91),
.B1(n_63),
.B2(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_95),
.Y(n_103)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_49),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_67),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_64),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_76),
.B(n_64),
.C(n_53),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_98),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_57),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_105),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_82),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_114),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_62),
.B(n_61),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_7),
.C(n_9),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_81),
.B1(n_56),
.B2(n_23),
.Y(n_118)
);

AOI22x1_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_56),
.B1(n_60),
.B2(n_55),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_123),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_130),
.B1(n_30),
.B2(n_33),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_3),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_4),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_4),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_26),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_13),
.C(n_17),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_5),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_6),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_124),
.B1(n_133),
.B2(n_120),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_97),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_129),
.C(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_142),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_108),
.B1(n_107),
.B2(n_105),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_145),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_148),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_122),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_152),
.C(n_155),
.Y(n_156)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_116),
.B1(n_115),
.B2(n_125),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_153),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_34),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_147),
.C(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_141),
.C(n_146),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_155),
.B1(n_142),
.B2(n_149),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_160),
.B1(n_156),
.B2(n_161),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_35),
.B(n_37),
.C(n_39),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_45),
.Y(n_165)
);


endmodule