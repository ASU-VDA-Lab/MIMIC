module fake_jpeg_23744_n_306 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_284;
wire n_288;
wire n_272;
wire n_265;
wire n_234;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_24),
.B1(n_33),
.B2(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_21),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_58),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_63),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_78),
.B(n_50),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_1),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_28),
.B1(n_26),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_70),
.B1(n_72),
.B2(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_68),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_18),
.B1(n_26),
.B2(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_44),
.B(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_75),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_23),
.B1(n_18),
.B2(n_27),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_39),
.B(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_47),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_28),
.B1(n_34),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_48),
.B1(n_39),
.B2(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_82),
.Y(n_120)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_47),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_43),
.B1(n_41),
.B2(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_94),
.B1(n_100),
.B2(n_116),
.Y(n_129)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_43),
.B1(n_34),
.B2(n_29),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_92),
.B(n_4),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_72),
.B1(n_56),
.B2(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_67),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_45),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_3),
.C(n_4),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_63),
.B(n_64),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_38),
.B1(n_31),
.B2(n_30),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_57),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_114),
.Y(n_141)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_76),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_55),
.A2(n_47),
.B1(n_31),
.B2(n_38),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_104),
.B(n_95),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_119),
.B(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_98),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_86),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_143),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_16),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_144),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_45),
.B(n_35),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_30),
.B(n_22),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_22),
.B(n_20),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_88),
.B1(n_87),
.B2(n_115),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_101),
.B1(n_89),
.B2(n_83),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_20),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_140),
.B(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_92),
.B(n_2),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_2),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_3),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_84),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_3),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_149),
.A2(n_83),
.B1(n_5),
.B2(n_6),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_82),
.B1(n_109),
.B2(n_80),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_140),
.B1(n_135),
.B2(n_126),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_133),
.A2(n_80),
.B1(n_110),
.B2(n_93),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_155),
.B1(n_130),
.B2(n_147),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_110),
.B1(n_93),
.B2(n_106),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_81),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_167),
.B1(n_172),
.B2(n_149),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_178),
.B(n_143),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_129),
.Y(n_183)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_137),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_179),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_15),
.Y(n_171)
);

NAND2x1_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_175),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_15),
.Y(n_175)
);

BUFx24_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_9),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_123),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_166),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_209),
.B1(n_205),
.B2(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_186),
.B(n_171),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_171),
.B(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_127),
.B1(n_126),
.B2(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_154),
.B1(n_155),
.B2(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_144),
.B1(n_122),
.B2(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_143),
.B(n_145),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_200),
.B(n_205),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_139),
.B(n_131),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_138),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_147),
.Y(n_202)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_206),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_147),
.Y(n_204)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_128),
.B(n_12),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_128),
.C(n_125),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_223),
.B1(n_209),
.B2(n_167),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_151),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_215),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_164),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_218),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_185),
.B(n_187),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_204),
.B(n_202),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_199),
.B1(n_182),
.B2(n_178),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_165),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_231),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_166),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_227),
.C(n_183),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_194),
.B(n_158),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_190),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_196),
.B(n_191),
.Y(n_227)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_153),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_238),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_237),
.A2(n_246),
.B1(n_232),
.B2(n_229),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_198),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_212),
.B1(n_221),
.B2(n_231),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_216),
.C(n_213),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_201),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_180),
.C(n_189),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_228),
.C(n_227),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_245),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_199),
.B(n_178),
.Y(n_247)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_178),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_158),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_161),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_253),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_211),
.C(n_219),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_211),
.C(n_219),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_224),
.C(n_225),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_260),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_216),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_214),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_261),
.B(n_263),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_242),
.C(n_232),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_247),
.B(n_248),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_264),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_235),
.B(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_268),
.Y(n_283)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_273),
.Y(n_282)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_245),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_277),
.B(n_268),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_275),
.C(n_251),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_284),
.Y(n_293)
);

AOI321xp33_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_258),
.A3(n_253),
.B1(n_250),
.B2(n_254),
.C(n_260),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_265),
.B(n_256),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_236),
.C(n_241),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_236),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_291),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_246),
.CI(n_239),
.CON(n_295),
.SN(n_295)
);

NOR2xp67_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_283),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_234),
.B(n_220),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_278),
.B(n_269),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_282),
.C(n_241),
.Y(n_294)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_295),
.A3(n_296),
.B1(n_234),
.B2(n_220),
.C1(n_230),
.C2(n_293),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_300),
.A3(n_301),
.B1(n_295),
.B2(n_176),
.C1(n_124),
.C2(n_165),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_274),
.A3(n_161),
.B1(n_184),
.B2(n_195),
.C1(n_163),
.C2(n_247),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_274),
.B(n_174),
.Y(n_301)
);

NOR3xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_303),
.C(n_14),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_11),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_14),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_15),
.Y(n_306)
);


endmodule