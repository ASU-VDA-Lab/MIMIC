module real_aes_10460_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_914, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_914;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_884;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_889;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_892;
wire n_372;
wire n_528;
wire n_202;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_298;
wire n_860;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g205 ( .A(n_0), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g610 ( .A(n_1), .Y(n_610) );
OAI22xp5_ASAP7_75t_SL g891 ( .A1(n_2), .A2(n_85), .B1(n_892), .B2(n_893), .Y(n_891) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_2), .Y(n_893) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_3), .B(n_543), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_4), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_5), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_6), .B(n_169), .Y(n_203) );
AOI22xp5_ASAP7_75t_SL g489 ( .A1(n_7), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_7), .Y(n_492) );
OAI22x1_ASAP7_75t_SL g486 ( .A1(n_8), .A2(n_101), .B1(n_487), .B2(n_488), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_8), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_9), .B(n_211), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_10), .Y(n_200) );
NOR2xp67_ASAP7_75t_L g115 ( .A(n_11), .B(n_93), .Y(n_115) );
INVx1_ASAP7_75t_L g909 ( .A(n_11), .Y(n_909) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_12), .B(n_164), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_13), .B(n_184), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_14), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_15), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_16), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_17), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_18), .B(n_187), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_19), .B(n_226), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_20), .B(n_164), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_21), .Y(n_603) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_22), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_23), .B(n_184), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_24), .B(n_211), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_25), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_26), .B(n_146), .Y(n_588) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_27), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_28), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_29), .B(n_146), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_30), .B(n_226), .Y(n_577) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_31), .Y(n_138) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_32), .A2(n_204), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_33), .B(n_184), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_34), .B(n_182), .Y(n_181) );
NAND2xp33_ASAP7_75t_SL g144 ( .A(n_35), .B(n_140), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_36), .B(n_184), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_37), .B(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_38), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_39), .A2(n_105), .B1(n_900), .B2(n_910), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_40), .B(n_137), .Y(n_255) );
INVx1_ASAP7_75t_L g114 ( .A(n_41), .Y(n_114) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_42), .A2(n_74), .B(n_132), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_43), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_44), .B(n_184), .Y(n_587) );
OAI22x1_ASAP7_75t_R g876 ( .A1(n_45), .A2(n_49), .B1(n_877), .B2(n_878), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_45), .Y(n_877) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_46), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_47), .B(n_173), .Y(n_243) );
AND2x6_ASAP7_75t_L g151 ( .A(n_48), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g878 ( .A(n_49), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_50), .B(n_128), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_51), .A2(n_89), .B1(n_543), .B2(n_561), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_52), .B(n_128), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_53), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_54), .B(n_158), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_55), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_56), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_57), .Y(n_626) );
INVx1_ASAP7_75t_L g152 ( .A(n_58), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_59), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_60), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_61), .B(n_561), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_62), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_63), .B(n_561), .Y(n_560) );
NAND2xp33_ASAP7_75t_L g139 ( .A(n_64), .B(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_65), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_65), .B(n_173), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_66), .B(n_158), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_67), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_68), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g905 ( .A(n_69), .B(n_906), .Y(n_905) );
INVx2_ASAP7_75t_L g619 ( .A(n_70), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_71), .B(n_146), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_72), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_73), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_75), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_76), .B(n_164), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_77), .B(n_226), .Y(n_239) );
INVx1_ASAP7_75t_L g613 ( .A(n_78), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_79), .B(n_173), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_80), .Y(n_533) );
BUFx10_ASAP7_75t_L g107 ( .A(n_81), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_82), .Y(n_501) );
INVx1_ASAP7_75t_L g527 ( .A(n_83), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_84), .B(n_164), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_85), .Y(n_892) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_86), .B(n_184), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_87), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_88), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_90), .B(n_158), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_91), .B(n_164), .Y(n_238) );
INVx1_ASAP7_75t_L g621 ( .A(n_92), .Y(n_621) );
AND2x2_ASAP7_75t_L g908 ( .A(n_93), .B(n_909), .Y(n_908) );
INVx2_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
OR2x2_ASAP7_75t_L g111 ( .A(n_95), .B(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_95), .B(n_113), .Y(n_505) );
BUFx2_ASAP7_75t_L g883 ( .A(n_95), .Y(n_883) );
INVx1_ASAP7_75t_L g907 ( .A(n_95), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_96), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_97), .B(n_182), .Y(n_253) );
INVx1_ASAP7_75t_L g906 ( .A(n_98), .Y(n_906) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_99), .B(n_211), .Y(n_218) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_100), .B(n_597), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_101), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_102), .Y(n_167) );
NAND2xp33_ASAP7_75t_L g539 ( .A(n_103), .B(n_158), .Y(n_539) );
AO211x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_108), .B(n_500), .C(n_506), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g504 ( .A(n_107), .Y(n_504) );
BUFx12f_ASAP7_75t_L g899 ( .A(n_107), .Y(n_899) );
AO21x1_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_116), .B(n_493), .Y(n_108) );
BUFx12f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_111), .Y(n_499) );
AND2x2_ASAP7_75t_L g882 ( .A(n_112), .B(n_883), .Y(n_882) );
AND2x4_ASAP7_75t_L g888 ( .A(n_112), .B(n_889), .Y(n_888) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g903 ( .A(n_114), .B(n_904), .C(n_907), .Y(n_903) );
XNOR2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_489), .Y(n_116) );
XNOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_486), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g884 ( .A1(n_118), .A2(n_879), .B(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_118), .B(n_886), .Y(n_885) );
NAND4xp75_ASAP7_75t_L g118 ( .A(n_119), .B(n_390), .C(n_432), .D(n_454), .Y(n_118) );
NOR2x1_ASAP7_75t_L g119 ( .A(n_120), .B(n_334), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_278), .C(n_310), .Y(n_120) );
AOI222xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_192), .B1(n_244), .B2(n_259), .C1(n_268), .C2(n_274), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI21xp33_ASAP7_75t_L g301 ( .A1(n_123), .A2(n_302), .B(n_306), .Y(n_301) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_154), .Y(n_123) );
OR2x2_ASAP7_75t_L g351 ( .A(n_124), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g389 ( .A(n_124), .Y(n_389) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_125), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g344 ( .A(n_125), .B(n_246), .Y(n_344) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g258 ( .A(n_126), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_126), .B(n_273), .Y(n_290) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_126), .Y(n_396) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_127), .Y(n_322) );
AND2x2_ASAP7_75t_L g375 ( .A(n_127), .B(n_247), .Y(n_375) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_133), .B(n_153), .Y(n_127) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_128), .A2(n_236), .B(n_243), .Y(n_235) );
INVx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g220 ( .A(n_129), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_129), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx5_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_130), .Y(n_191) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_143), .B(n_149), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_139), .C(n_141), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_136), .A2(n_627), .B1(n_633), .B2(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g187 ( .A(n_137), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_137), .A2(n_184), .B1(n_199), .B2(n_200), .Y(n_198) );
INVx2_ASAP7_75t_L g543 ( .A(n_137), .Y(n_543) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_138), .Y(n_140) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_138), .Y(n_147) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_138), .Y(n_164) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx1_ASAP7_75t_L g212 ( .A(n_138), .Y(n_212) );
INVx2_ASAP7_75t_L g217 ( .A(n_140), .Y(n_217) );
INVx2_ASAP7_75t_L g561 ( .A(n_140), .Y(n_561) );
INVx2_ASAP7_75t_L g598 ( .A(n_140), .Y(n_598) );
INVx2_ASAP7_75t_L g600 ( .A(n_140), .Y(n_600) );
INVx2_ASAP7_75t_SL g148 ( .A(n_141), .Y(n_148) );
INVx2_ASAP7_75t_SL g165 ( .A(n_141), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_141), .A2(n_181), .B(n_183), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_141), .A2(n_225), .B(n_227), .Y(n_224) );
CKINVDCx6p67_ASAP7_75t_R g541 ( .A(n_141), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_141), .A2(n_587), .B(n_588), .Y(n_586) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx5_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
BUFx12f_ASAP7_75t_L g204 ( .A(n_142), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_148), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_146), .B(n_533), .Y(n_532) );
INVxp67_ASAP7_75t_L g548 ( .A(n_146), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_146), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
INVx2_ASAP7_75t_L g169 ( .A(n_147), .Y(n_169) );
INVx2_ASAP7_75t_L g182 ( .A(n_147), .Y(n_182) );
INVx2_ASAP7_75t_L g627 ( .A(n_147), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_148), .A2(n_186), .B(n_188), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_148), .A2(n_151), .B(n_198), .C(n_201), .Y(n_197) );
AOI21x1_ASAP7_75t_L g228 ( .A1(n_148), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_148), .A2(n_590), .B(n_591), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_149), .A2(n_160), .B(n_166), .Y(n_159) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_149), .A2(n_224), .B(n_228), .Y(n_223) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_149), .A2(n_586), .B(n_589), .Y(n_585) );
INVx2_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
INVx8_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_150), .A2(n_173), .B(n_535), .Y(n_534) );
INVx8_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI21x1_ASAP7_75t_SL g208 ( .A1(n_151), .A2(n_209), .B(n_215), .Y(n_208) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_151), .A2(n_237), .B(n_240), .Y(n_236) );
INVx1_ASAP7_75t_L g551 ( .A(n_151), .Y(n_551) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_151), .A2(n_174), .B(n_620), .Y(n_622) );
INVx1_ASAP7_75t_L g630 ( .A(n_151), .Y(n_630) );
INVx1_ASAP7_75t_L g373 ( .A(n_154), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_176), .Y(n_154) );
INVx1_ASAP7_75t_L g347 ( .A(n_155), .Y(n_347) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g269 ( .A(n_156), .B(n_248), .Y(n_269) );
INVx2_ASAP7_75t_L g288 ( .A(n_156), .Y(n_288) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g353 ( .A(n_157), .Y(n_353) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_172), .Y(n_157) );
OAI21x1_ASAP7_75t_L g178 ( .A1(n_158), .A2(n_179), .B(n_190), .Y(n_178) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_158), .A2(n_197), .B(n_205), .Y(n_196) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_158), .A2(n_250), .B(n_257), .Y(n_249) );
NOR2x1p5_ASAP7_75t_SL g550 ( .A(n_158), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g594 ( .A(n_158), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_165), .Y(n_160) );
INVx5_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
OR2x2_ASAP7_75t_L g529 ( .A(n_164), .B(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_165), .A2(n_241), .B(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_165), .A2(n_252), .B(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_165), .A2(n_547), .B(n_548), .C(n_549), .Y(n_546) );
O2A1O1Ixp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_170), .C(n_171), .Y(n_166) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_171), .A2(n_210), .B(n_211), .C(n_213), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_171), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_171), .A2(n_255), .B(n_256), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_171), .A2(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g579 ( .A(n_171), .Y(n_579) );
OAI21xp33_ASAP7_75t_L g624 ( .A1(n_171), .A2(n_625), .B(n_629), .Y(n_624) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_174), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_174), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_175), .Y(n_206) );
AND2x2_ASAP7_75t_L g313 ( .A(n_176), .B(n_262), .Y(n_313) );
BUFx2_ASAP7_75t_L g443 ( .A(n_176), .Y(n_443) );
AND2x2_ASAP7_75t_L g479 ( .A(n_176), .B(n_195), .Y(n_479) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx3_ASAP7_75t_L g343 ( .A(n_177), .Y(n_343) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g273 ( .A(n_178), .Y(n_273) );
OAI21x1_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_185), .B(n_189), .Y(n_179) );
INVx2_ASAP7_75t_L g523 ( .A(n_184), .Y(n_523) );
INVx2_ASAP7_75t_L g574 ( .A(n_184), .Y(n_574) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_189), .A2(n_251), .B(n_254), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_189), .A2(n_558), .B(n_562), .Y(n_557) );
OAI21x1_ASAP7_75t_SL g570 ( .A1(n_189), .A2(n_571), .B(n_576), .Y(n_570) );
AO31x2_ASAP7_75t_L g593 ( .A1(n_189), .A2(n_594), .A3(n_595), .B(n_602), .Y(n_593) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_221), .Y(n_194) );
INVx1_ASAP7_75t_L g473 ( .A(n_195), .Y(n_473) );
AND2x2_ASAP7_75t_L g480 ( .A(n_195), .B(n_294), .Y(n_480) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_207), .Y(n_195) );
INVx3_ASAP7_75t_L g262 ( .A(n_196), .Y(n_262) );
AND2x2_ASAP7_75t_L g275 ( .A(n_196), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g293 ( .A(n_196), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_204), .A2(n_216), .B(n_218), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_204), .Y(n_525) );
INVx3_ASAP7_75t_L g575 ( .A(n_204), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_204), .A2(n_596), .B1(n_599), .B2(n_601), .Y(n_595) );
BUFx2_ASAP7_75t_L g614 ( .A(n_204), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_204), .B(n_632), .Y(n_631) );
OAI21x1_ASAP7_75t_L g207 ( .A1(n_206), .A2(n_208), .B(n_219), .Y(n_207) );
BUFx4f_ASAP7_75t_L g232 ( .A(n_206), .Y(n_232) );
INVx3_ASAP7_75t_L g556 ( .A(n_206), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_206), .B(n_630), .Y(n_629) );
INVx3_ASAP7_75t_L g267 ( .A(n_207), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_211), .A2(n_522), .B1(n_523), .B2(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g214 ( .A(n_212), .Y(n_214) );
INVx2_ASAP7_75t_L g231 ( .A(n_214), .Y(n_231) );
INVx2_ASAP7_75t_L g617 ( .A(n_217), .Y(n_617) );
INVx1_ASAP7_75t_L g371 ( .A(n_221), .Y(n_371) );
INVx2_ASAP7_75t_L g415 ( .A(n_221), .Y(n_415) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_234), .Y(n_221) );
BUFx2_ASAP7_75t_L g265 ( .A(n_222), .Y(n_265) );
AND2x2_ASAP7_75t_L g325 ( .A(n_222), .B(n_235), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_232), .B(n_233), .Y(n_222) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_223), .A2(n_232), .B(n_233), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_226), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_226), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_616) );
OAI21x1_ASAP7_75t_SL g569 ( .A1(n_232), .A2(n_570), .B(n_580), .Y(n_569) );
OAI21x1_ASAP7_75t_L g584 ( .A1(n_232), .A2(n_585), .B(n_592), .Y(n_584) );
INVx1_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
NOR2xp67_ASAP7_75t_L g282 ( .A(n_234), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g300 ( .A(n_234), .B(n_267), .Y(n_300) );
AND2x2_ASAP7_75t_L g338 ( .A(n_234), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_234), .Y(n_357) );
INVx1_ASAP7_75t_L g364 ( .A(n_234), .Y(n_364) );
INVx1_ASAP7_75t_L g485 ( .A(n_234), .Y(n_485) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
BUFx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g466 ( .A(n_245), .Y(n_466) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_258), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g298 ( .A(n_248), .B(n_288), .Y(n_298) );
INVx1_ASAP7_75t_L g321 ( .A(n_248), .Y(n_321) );
INVx1_ASAP7_75t_L g349 ( .A(n_248), .Y(n_349) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g305 ( .A(n_258), .Y(n_305) );
AND2x2_ASAP7_75t_L g399 ( .A(n_258), .B(n_273), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_259), .A2(n_269), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_264), .Y(n_259) );
AND2x4_ASAP7_75t_L g330 ( .A(n_260), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_260), .B(n_264), .Y(n_424) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
AND2x2_ASAP7_75t_L g309 ( .A(n_261), .B(n_267), .Y(n_309) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g337 ( .A(n_262), .B(n_276), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_262), .B(n_267), .Y(n_405) );
AND2x2_ASAP7_75t_L g417 ( .A(n_262), .B(n_339), .Y(n_417) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g308 ( .A(n_265), .Y(n_308) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_265), .Y(n_472) );
INVx1_ASAP7_75t_L g381 ( .A(n_266), .Y(n_381) );
AND2x2_ASAP7_75t_L g455 ( .A(n_266), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g283 ( .A(n_267), .Y(n_283) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_267), .Y(n_324) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_267), .Y(n_332) );
INVx2_ASAP7_75t_SL g339 ( .A(n_267), .Y(n_339) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x2_ASAP7_75t_L g398 ( .A(n_269), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g463 ( .A(n_269), .B(n_443), .Y(n_463) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g318 ( .A(n_272), .Y(n_318) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_272), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2x1_ASAP7_75t_L g356 ( .A(n_275), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g462 ( .A(n_275), .B(n_338), .Y(n_462) );
INVx2_ASAP7_75t_SL g294 ( .A(n_276), .Y(n_294) );
AND2x4_ASAP7_75t_L g363 ( .A(n_276), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_R g333 ( .A(n_277), .Y(n_333) );
NOR2xp33_ASAP7_75t_SL g278 ( .A(n_279), .B(n_301), .Y(n_278) );
OAI31xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .A3(n_291), .B(n_295), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g460 ( .A(n_282), .B(n_337), .Y(n_460) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_283), .Y(n_393) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g379 ( .A(n_288), .Y(n_379) );
AND2x2_ASAP7_75t_L g401 ( .A(n_288), .B(n_349), .Y(n_401) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g328 ( .A(n_290), .Y(n_328) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_293), .B(n_363), .Y(n_362) );
INVx4_ASAP7_75t_L g370 ( .A(n_293), .Y(n_370) );
AND2x4_ASAP7_75t_L g299 ( .A(n_294), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g403 ( .A(n_294), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_296), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g329 ( .A(n_297), .Y(n_329) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g303 ( .A(n_298), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g395 ( .A(n_298), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g439 ( .A(n_299), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g315 ( .A(n_300), .Y(n_315) );
AND2x2_ASAP7_75t_L g410 ( .A(n_300), .B(n_333), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_300), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g451 ( .A(n_300), .B(n_370), .Y(n_451) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_303), .B(n_408), .Y(n_407) );
AOI31xp33_ASAP7_75t_L g433 ( .A1(n_303), .A2(n_381), .A3(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g366 ( .A(n_305), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g469 ( .A(n_305), .Y(n_469) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_308), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g408 ( .A(n_308), .B(n_338), .Y(n_408) );
INVx1_ASAP7_75t_L g434 ( .A(n_308), .Y(n_434) );
AND2x2_ASAP7_75t_L g385 ( .A(n_309), .B(n_325), .Y(n_385) );
AND2x2_ASAP7_75t_L g436 ( .A(n_309), .B(n_363), .Y(n_436) );
AOI222xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B1(n_316), .B2(n_323), .C1(n_326), .C2(n_330), .Y(n_310) );
BUFx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OR2x2_ASAP7_75t_L g421 ( .A(n_318), .B(n_320), .Y(n_421) );
OA211x2_ASAP7_75t_L g432 ( .A1(n_318), .A2(n_433), .B(n_437), .C(n_441), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g481 ( .A1(n_319), .A2(n_329), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_324), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_325), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g446 ( .A(n_325), .Y(n_446) );
AND2x2_ASAP7_75t_L g465 ( .A(n_325), .B(n_417), .Y(n_465) );
NOR2xp67_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g448 ( .A(n_327), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g435 ( .A(n_329), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_332), .B(n_485), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_360), .C(n_376), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B1(n_350), .B2(n_354), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx2_ASAP7_75t_L g431 ( .A(n_337), .Y(n_431) );
INVx1_ASAP7_75t_L g382 ( .A(n_338), .Y(n_382) );
NAND2xp33_ASAP7_75t_SL g340 ( .A(n_341), .B(n_345), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
AND2x4_ASAP7_75t_SL g383 ( .A(n_342), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g427 ( .A(n_342), .Y(n_427) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g346 ( .A(n_343), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g387 ( .A(n_343), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
OAI22xp33_ASAP7_75t_R g477 ( .A1(n_344), .A2(n_371), .B1(n_403), .B2(n_478), .Y(n_477) );
NAND2x1_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g367 ( .A(n_346), .Y(n_367) );
AND2x2_ASAP7_75t_L g475 ( .A(n_346), .B(n_384), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_347), .B(n_349), .Y(n_452) );
AND2x4_ASAP7_75t_L g411 ( .A(n_348), .B(n_412), .Y(n_411) );
OAI32xp33_ASAP7_75t_L g442 ( .A1(n_348), .A2(n_362), .A3(n_443), .B1(n_444), .B2(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g478 ( .A(n_348), .Y(n_478) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g412 ( .A(n_352), .Y(n_412) );
INVx1_ASAP7_75t_L g445 ( .A(n_352), .Y(n_445) );
OAI22xp33_ASAP7_75t_SL g377 ( .A1(n_353), .A2(n_378), .B1(n_380), .B2(n_382), .Y(n_377) );
INVx2_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
OR2x2_ASAP7_75t_L g392 ( .A(n_356), .B(n_393), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_365), .B1(n_368), .B2(n_372), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_363), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g437 ( .A1(n_365), .A2(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_369), .A2(n_388), .B1(n_392), .B2(n_394), .C(n_397), .Y(n_391) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AOI33xp33_ASAP7_75t_L g376 ( .A1(n_370), .A2(n_377), .A3(n_383), .B1(n_385), .B2(n_386), .B3(n_389), .Y(n_376) );
INVx1_ASAP7_75t_L g440 ( .A(n_370), .Y(n_440) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx2_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_375), .A2(n_419), .B(n_420), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_375), .B(n_445), .Y(n_444) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AOI32xp33_ASAP7_75t_L g464 ( .A1(n_387), .A2(n_465), .A3(n_466), .B1(n_467), .B2(n_914), .Y(n_464) );
AND2x4_ASAP7_75t_SL g423 ( .A(n_388), .B(n_399), .Y(n_423) );
NOR3x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_406), .C(n_413), .Y(n_390) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g457 ( .A(n_395), .B(n_443), .Y(n_457) );
AND2x2_ASAP7_75t_L g400 ( .A(n_396), .B(n_401), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_402), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_398), .A2(n_477), .B1(n_479), .B2(n_480), .Y(n_476) );
AND2x2_ASAP7_75t_L g426 ( .A(n_401), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_408), .A2(n_423), .B1(n_462), .B2(n_463), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g449 ( .A(n_412), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_418), .B1(n_422), .B2(n_424), .C(n_425), .Y(n_413) );
OR2x6_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g438 ( .A(n_419), .Y(n_438) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x6_ASAP7_75t_L g483 ( .A(n_431), .B(n_484), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_447), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B1(n_452), .B2(n_453), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp33_ASAP7_75t_L g453 ( .A(n_451), .Y(n_453) );
OR2x2_ASAP7_75t_L g468 ( .A(n_452), .B(n_469), .Y(n_468) );
AOI211x1_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_457), .B(n_458), .C(n_470), .Y(n_454) );
NAND3xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_461), .C(n_464), .Y(n_458) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
OAI211xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_474), .B(n_476), .C(n_481), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g897 ( .A(n_493), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx6_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx5_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_R g500 ( .A(n_501), .B(n_502), .Y(n_500) );
BUFx12f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AOI31xp67_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_894), .A3(n_897), .B(n_898), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_508), .B(n_890), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_881), .B1(n_884), .B2(n_887), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_510), .A2(n_881), .B1(n_887), .B2(n_896), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_876), .B1(n_879), .B2(n_880), .Y(n_510) );
INVx3_ASAP7_75t_L g880 ( .A(n_511), .Y(n_880) );
AND3x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_754), .C(n_825), .Y(n_511) );
NOR2x1_ASAP7_75t_L g512 ( .A(n_513), .B(n_704), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_652), .C(n_691), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_566), .B(n_581), .C(n_636), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NOR2xp67_ASAP7_75t_L g809 ( .A(n_516), .B(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_536), .Y(n_516) );
INVx1_ASAP7_75t_L g729 ( .A(n_517), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_517), .B(n_686), .Y(n_821) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_518), .B(n_538), .Y(n_688) );
AND2x2_ASAP7_75t_L g725 ( .A(n_518), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g753 ( .A(n_518), .B(n_568), .Y(n_753) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g641 ( .A(n_519), .Y(n_641) );
BUFx3_ASAP7_75t_L g690 ( .A(n_519), .Y(n_690) );
OAI21x1_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_528), .B(n_534), .Y(n_519) );
AO21x1_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_525), .B(n_526), .Y(n_520) );
INVx2_ASAP7_75t_L g611 ( .A(n_523), .Y(n_611) );
AOI21x1_ASAP7_75t_L g528 ( .A1(n_525), .A2(n_529), .B(n_531), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_525), .A2(n_616), .B(n_620), .Y(n_615) );
INVxp67_ASAP7_75t_L g535 ( .A(n_526), .Y(n_535) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_552), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_537), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_537), .Y(n_643) );
AND2x2_ASAP7_75t_L g846 ( .A(n_537), .B(n_568), .Y(n_846) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g658 ( .A(n_538), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_538), .B(n_645), .Y(n_671) );
INVx1_ASAP7_75t_L g684 ( .A(n_538), .Y(n_684) );
INVx1_ASAP7_75t_L g726 ( .A(n_538), .Y(n_726) );
AND2x2_ASAP7_75t_L g739 ( .A(n_538), .B(n_659), .Y(n_739) );
AND2x2_ASAP7_75t_L g780 ( .A(n_538), .B(n_640), .Y(n_780) );
HB1xp67_ASAP7_75t_SL g795 ( .A(n_538), .Y(n_795) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_546), .C(n_550), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_541), .A2(n_559), .B(n_560), .Y(n_558) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_543), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_625) );
AND2x4_ASAP7_75t_L g566 ( .A(n_552), .B(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g722 ( .A(n_552), .B(n_568), .Y(n_722) );
BUFx2_ASAP7_75t_L g743 ( .A(n_552), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_552), .B(n_769), .Y(n_771) );
INVx1_ASAP7_75t_L g865 ( .A(n_552), .Y(n_865) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g689 ( .A(n_553), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g645 ( .A(n_554), .Y(n_645) );
OAI21x1_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_557), .B(n_565), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
O2A1O1Ixp5_ASAP7_75t_L g636 ( .A1(n_566), .A2(n_637), .B(n_642), .C(n_646), .Y(n_636) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g644 ( .A(n_568), .B(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g819 ( .A(n_568), .Y(n_819) );
BUFx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g659 ( .A(n_569), .Y(n_659) );
AOI21x1_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B(n_575), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_579), .Y(n_576) );
INVx2_ASAP7_75t_L g734 ( .A(n_581), .Y(n_734) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_604), .Y(n_581) );
INVx2_ASAP7_75t_L g647 ( .A(n_582), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_582), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g765 ( .A(n_582), .Y(n_765) );
AND2x2_ASAP7_75t_L g813 ( .A(n_582), .B(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g829 ( .A(n_582), .B(n_830), .Y(n_829) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_593), .Y(n_582) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_583), .Y(n_665) );
AND2x4_ASAP7_75t_L g697 ( .A(n_583), .B(n_698), .Y(n_697) );
BUFx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g702 ( .A(n_584), .Y(n_702) );
AND2x2_ASAP7_75t_L g667 ( .A(n_593), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_SL g681 ( .A(n_593), .Y(n_681) );
INVx2_ASAP7_75t_L g698 ( .A(n_593), .Y(n_698) );
AND2x2_ASAP7_75t_L g717 ( .A(n_593), .B(n_702), .Y(n_717) );
INVx1_ASAP7_75t_L g747 ( .A(n_593), .Y(n_747) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g785 ( .A(n_604), .B(n_697), .Y(n_785) );
AND2x4_ASAP7_75t_L g807 ( .A(n_604), .B(n_665), .Y(n_807) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g693 ( .A(n_605), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g870 ( .A(n_605), .Y(n_870) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_623), .Y(n_605) );
AND2x2_ASAP7_75t_L g674 ( .A(n_606), .B(n_623), .Y(n_674) );
INVx2_ASAP7_75t_L g679 ( .A(n_606), .Y(n_679) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g651 ( .A(n_607), .Y(n_651) );
AO21x2_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_615), .B(n_622), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B(n_614), .Y(n_608) );
NOR2x1_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_SL g650 ( .A(n_623), .Y(n_650) );
INVx1_ASAP7_75t_L g668 ( .A(n_623), .Y(n_668) );
AND2x4_ASAP7_75t_L g680 ( .A(n_623), .B(n_681), .Y(n_680) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_623), .Y(n_764) );
AND2x2_ASAP7_75t_L g789 ( .A(n_623), .B(n_702), .Y(n_789) );
AND2x2_ASAP7_75t_L g814 ( .A(n_623), .B(n_679), .Y(n_814) );
OA21x2_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_631), .B(n_635), .Y(n_623) );
AOI322xp5_ASAP7_75t_L g812 ( .A1(n_637), .A2(n_661), .A3(n_783), .B1(n_813), .B2(n_815), .C1(n_816), .C2(n_822), .Y(n_812) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g655 ( .A(n_640), .Y(n_655) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_641), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x4_ASAP7_75t_SL g752 ( .A(n_643), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g793 ( .A(n_643), .Y(n_793) );
BUFx2_ASAP7_75t_L g703 ( .A(n_644), .Y(n_703) );
AND2x2_ASAP7_75t_L g872 ( .A(n_644), .B(n_780), .Y(n_872) );
INVx2_ASAP7_75t_L g661 ( .A(n_645), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_645), .B(n_659), .Y(n_731) );
OR2x6_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVxp67_ASAP7_75t_L g799 ( .A(n_647), .Y(n_799) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_SL g732 ( .A(n_649), .B(n_697), .Y(n_732) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g709 ( .A(n_650), .B(n_702), .Y(n_709) );
INVx2_ASAP7_75t_L g711 ( .A(n_651), .Y(n_711) );
AND2x2_ASAP7_75t_L g777 ( .A(n_651), .B(n_695), .Y(n_777) );
AND2x2_ASAP7_75t_L g849 ( .A(n_651), .B(n_702), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_662), .B(n_669), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
OR2x2_ASAP7_75t_L g670 ( .A(n_655), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g719 ( .A(n_655), .Y(n_719) );
AO32x1_ASAP7_75t_L g713 ( .A1(n_656), .A2(n_714), .A3(n_718), .B1(n_719), .B2(n_720), .Y(n_713) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_657), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g742 ( .A(n_657), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g776 ( .A(n_657), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g837 ( .A(n_657), .Y(n_837) );
BUFx2_ASAP7_75t_L g853 ( .A(n_657), .Y(n_853) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g686 ( .A(n_659), .Y(n_686) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g779 ( .A(n_661), .B(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g783 ( .A(n_661), .B(n_725), .Y(n_783) );
AND2x2_ASAP7_75t_L g804 ( .A(n_661), .B(n_739), .Y(n_804) );
AND2x2_ASAP7_75t_L g832 ( .A(n_661), .B(n_833), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g869 ( .A(n_664), .B(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g745 ( .A(n_665), .Y(n_745) );
OR2x2_ASAP7_75t_L g749 ( .A(n_665), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_665), .B(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g855 ( .A(n_667), .B(n_849), .Y(n_855) );
AND2x2_ASAP7_75t_L g746 ( .A(n_668), .B(n_747), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B1(n_675), .B2(n_682), .Y(n_669) );
BUFx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g736 ( .A(n_674), .B(n_717), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_674), .B(n_700), .Y(n_808) );
INVx2_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g758 ( .A(n_678), .B(n_680), .Y(n_758) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_L g788 ( .A(n_679), .B(n_698), .Y(n_788) );
INVx2_ASAP7_75t_L g750 ( .A(n_680), .Y(n_750) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_680), .Y(n_775) );
AND2x2_ASAP7_75t_L g848 ( .A(n_680), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g712 ( .A(n_681), .Y(n_712) );
AOI211xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_685), .B(n_687), .C(n_689), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_683), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g820 ( .A(n_684), .B(n_821), .Y(n_820) );
AO22x1_ASAP7_75t_L g696 ( .A1(n_685), .A2(n_697), .B1(n_699), .B2(n_703), .Y(n_696) );
INVx1_ASAP7_75t_L g718 ( .A(n_685), .Y(n_718) );
BUFx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_687), .B(n_722), .Y(n_801) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g833 ( .A(n_688), .Y(n_833) );
INVx1_ASAP7_75t_L g707 ( .A(n_689), .Y(n_707) );
AND2x4_ASAP7_75t_L g818 ( .A(n_689), .B(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g695 ( .A(n_690), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_696), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g845 ( .A(n_694), .B(n_846), .Y(n_845) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_694), .Y(n_857) );
OR2x2_ASAP7_75t_L g874 ( .A(n_694), .B(n_772), .Y(n_874) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_SL g720 ( .A(n_697), .B(n_716), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g842 ( .A(n_699), .B(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_L g828 ( .A(n_700), .B(n_788), .Y(n_828) );
OR2x2_ASAP7_75t_L g839 ( .A(n_700), .B(n_750), .Y(n_839) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_702), .B(n_711), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_721), .C(n_740), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .B(n_713), .Y(n_705) );
AND2x4_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
AND2x2_ASAP7_75t_L g811 ( .A(n_709), .B(n_788), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_709), .B(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx2_ASAP7_75t_L g716 ( .A(n_711), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_711), .B(n_712), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_714), .A2(n_779), .B1(n_864), .B2(n_866), .Y(n_863) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g796 ( .A(n_716), .Y(n_796) );
INVx1_ASAP7_75t_L g861 ( .A(n_717), .Y(n_861) );
OAI322xp33_ASAP7_75t_L g840 ( .A1(n_719), .A2(n_841), .A3(n_842), .B1(n_844), .B2(n_847), .C1(n_850), .C2(n_854), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_720), .A2(n_835), .B1(n_836), .B2(n_838), .Y(n_834) );
A2O1A1O1Ixp25_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_727), .C(n_732), .D(n_733), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_722), .B(n_724), .Y(n_835) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_725), .Y(n_760) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
AND2x2_ASAP7_75t_L g767 ( .A(n_730), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_731), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_737), .Y(n_733) );
INVx2_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g772 ( .A(n_739), .Y(n_772) );
NOR2xp67_ASAP7_75t_L g740 ( .A(n_741), .B(n_748), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx2_ASAP7_75t_L g841 ( .A(n_742), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_742), .B(n_815), .Y(n_875) );
INVx1_ASAP7_75t_L g797 ( .A(n_743), .Y(n_797) );
INVxp67_ASAP7_75t_L g873 ( .A(n_744), .Y(n_873) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
AND2x2_ASAP7_75t_L g815 ( .A(n_745), .B(n_814), .Y(n_815) );
INVx2_ASAP7_75t_L g794 ( .A(n_746), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_753), .B(n_791), .C(n_796), .D(n_797), .Y(n_790) );
AND4x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_778), .C(n_798), .D(n_812), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_759), .B(n_761), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_756), .A2(n_779), .B(n_781), .Y(n_778) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI221xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_766), .B1(n_770), .B2(n_773), .C(n_774), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g830 ( .A(n_764), .Y(n_830) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_768), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
OAI211xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_784), .B(n_786), .C(n_790), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_SL g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g792 ( .A(n_789), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_794), .B2(n_795), .Y(n_791) );
AOI221x1_ASAP7_75t_SL g798 ( .A1(n_799), .A2(n_800), .B1(n_802), .B2(n_805), .C(n_809), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_808), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g866 ( .A(n_808), .Y(n_866) );
INVx2_ASAP7_75t_SL g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g862 ( .A(n_814), .Y(n_862) );
NAND2xp5_ASAP7_75t_SL g816 ( .A(n_817), .B(n_820), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NOR4xp25_ASAP7_75t_L g825 ( .A(n_826), .B(n_840), .C(n_856), .D(n_867), .Y(n_825) );
OAI21xp33_ASAP7_75t_SL g826 ( .A1(n_827), .A2(n_831), .B(n_834), .Y(n_826) );
NOR2xp67_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g843 ( .A(n_830), .Y(n_843) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx3_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
AND2x4_ASAP7_75t_L g864 ( .A(n_846), .B(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_853), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_853), .B(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OAI21xp33_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B(n_863), .Y(n_856) );
INVx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
OR2x2_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
OAI221xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_871), .B1(n_873), .B2(n_874), .C(n_875), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVxp67_ASAP7_75t_R g879 ( .A(n_876), .Y(n_879) );
INVx1_ASAP7_75t_L g886 ( .A(n_876), .Y(n_886) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_883), .Y(n_889) );
INVx1_ASAP7_75t_L g896 ( .A(n_884), .Y(n_896) );
INVx1_ASAP7_75t_SL g887 ( .A(n_888), .Y(n_887) );
INVxp33_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_SL g894 ( .A(n_891), .B(n_895), .Y(n_894) );
INVx11_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
BUFx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
BUFx5_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
BUFx4f_ASAP7_75t_L g912 ( .A(n_902), .Y(n_912) );
AND2x2_ASAP7_75t_SL g902 ( .A(n_903), .B(n_908), .Y(n_902) );
INVx4_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVxp67_ASAP7_75t_SL g910 ( .A(n_911), .Y(n_910) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
endmodule