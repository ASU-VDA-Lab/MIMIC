module fake_jpeg_19606_n_39 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_1),
.B(n_2),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_26),
.B(n_2),
.Y(n_27)
);

OAI32xp33_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_8),
.A3(n_13),
.B1(n_10),
.B2(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx12f_ASAP7_75t_SL g32 ( 
.A(n_28),
.Y(n_32)
);

AO221x1_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_28),
.B1(n_24),
.B2(n_26),
.C(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_4),
.B2(n_5),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_7),
.B(n_15),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_5),
.B(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_33),
.Y(n_39)
);


endmodule