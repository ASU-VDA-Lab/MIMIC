module fake_jpeg_745_n_83 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_37),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_30),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_28),
.B1(n_35),
.B2(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_47),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_28),
.B1(n_27),
.B2(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_50),
.B1(n_40),
.B2(n_2),
.Y(n_55)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_12),
.Y(n_60)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_68)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_65),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_58),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_59),
.C(n_20),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_15),
.Y(n_69)
);

XNOR2x1_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_74),
.Y(n_76)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_75),
.A2(n_66),
.A3(n_70),
.B1(n_64),
.B2(n_65),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_76),
.B(n_75),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_72),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_22),
.Y(n_83)
);


endmodule