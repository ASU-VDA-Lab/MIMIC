module fake_ibex_1945_n_2867 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_545, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_568, n_52, n_448, n_99, n_466, n_269, n_156, n_570, n_126, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_558, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_267, n_245, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_572, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_2867);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_2867;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_2847;
wire n_1308;
wire n_1138;
wire n_708;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2347;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2436;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_2090;
wire n_666;
wire n_2260;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_702;
wire n_1326;
wire n_971;
wire n_1350;
wire n_906;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_2723;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_660;
wire n_2590;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_916;
wire n_2298;
wire n_2771;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_961;
wire n_991;
wire n_634;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_2862;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_2617;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_1673;
wire n_2018;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2251;
wire n_722;
wire n_2012;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1871;
wire n_1642;
wire n_2182;
wire n_2447;
wire n_2818;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2861;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_2669;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_2518;
wire n_2784;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_2734;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2652;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_999;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_1142;
wire n_783;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2148;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_2092;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2704;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_2754;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_1534;
wire n_908;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;

INVx1_ASAP7_75t_L g573 ( 
.A(n_76),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_565),
.Y(n_574)
);

BUFx5_ASAP7_75t_L g575 ( 
.A(n_508),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_223),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_511),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_473),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_264),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_557),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_243),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_336),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_357),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_192),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_266),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_78),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_382),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_139),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_480),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_146),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_325),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_525),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_92),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_393),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_412),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_449),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_348),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_153),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_117),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_91),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_324),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_291),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_136),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_436),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_19),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_123),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_109),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_126),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_44),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_300),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_164),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_16),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_498),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_164),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_439),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_2),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_302),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_355),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_359),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_560),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_419),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_255),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_219),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_260),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_500),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_83),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_200),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_492),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_281),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_419),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_150),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_150),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_235),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_110),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_151),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_571),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_548),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_28),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_301),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_193),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_188),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_L g642 ( 
.A(n_541),
.B(n_196),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_12),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_450),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_372),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_442),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_248),
.Y(n_647)
);

CKINVDCx14_ASAP7_75t_R g648 ( 
.A(n_499),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_491),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_302),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_343),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_376),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_280),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_138),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_100),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_145),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_58),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_15),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_183),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_505),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_135),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_556),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_372),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_249),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_L g665 ( 
.A(n_429),
.B(n_572),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_50),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_438),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_347),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_181),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_80),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_330),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_469),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_358),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_544),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_373),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_547),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_358),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_211),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_527),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_416),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_403),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_81),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_530),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_208),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_179),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_451),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_280),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_337),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_271),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_569),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_338),
.B(n_92),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_502),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_38),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_558),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_324),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_268),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_256),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_106),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_495),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_463),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_398),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_549),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_94),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_534),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_353),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_231),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_308),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_562),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_335),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_294),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_414),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_17),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_179),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_115),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_567),
.Y(n_715)
);

NOR2xp67_ASAP7_75t_L g716 ( 
.A(n_112),
.B(n_229),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_404),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_283),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_23),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_182),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_465),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_361),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_550),
.Y(n_723)
);

CKINVDCx14_ASAP7_75t_R g724 ( 
.A(n_189),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_138),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_264),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_414),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_47),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_39),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_239),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_82),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_0),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_361),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_289),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_58),
.Y(n_735)
);

BUFx5_ASAP7_75t_L g736 ( 
.A(n_231),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_507),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_546),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_121),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_80),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_432),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_31),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_104),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_L g744 ( 
.A(n_516),
.B(n_176),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_63),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_134),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_282),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_12),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_295),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_382),
.Y(n_750)
);

BUFx8_ASAP7_75t_SL g751 ( 
.A(n_420),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_35),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_208),
.Y(n_753)
);

NOR2xp67_ASAP7_75t_L g754 ( 
.A(n_169),
.B(n_438),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_54),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_305),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_22),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_40),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_10),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_332),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_493),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_529),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_256),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_363),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_205),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_190),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_568),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_137),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_415),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_308),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_517),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_241),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_228),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_359),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_251),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_459),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_115),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_L g778 ( 
.A(n_199),
.B(n_528),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_237),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_303),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_445),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_563),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_275),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_490),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_141),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_303),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_178),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_200),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_171),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_252),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_427),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_59),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_497),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_535),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_533),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_399),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_430),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_266),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_235),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_118),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_196),
.B(n_401),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_494),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_55),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_521),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_187),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_488),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_250),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_466),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_177),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_145),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_269),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_219),
.Y(n_812)
);

CKINVDCx14_ASAP7_75t_R g813 ( 
.A(n_254),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_161),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_411),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_522),
.Y(n_816)
);

CKINVDCx16_ASAP7_75t_R g817 ( 
.A(n_564),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_49),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_524),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_124),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_222),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_434),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_13),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_136),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_555),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_117),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_449),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_360),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_147),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_224),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_261),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_489),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_496),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_116),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_327),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_2),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_269),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_483),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_526),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_566),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_450),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_177),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_1),
.Y(n_843)
);

BUFx2_ASAP7_75t_SL g844 ( 
.A(n_515),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_559),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_342),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_8),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_345),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_193),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_380),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_369),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_561),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_74),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_283),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_286),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_504),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_337),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_194),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_152),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_197),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_476),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_186),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_481),
.Y(n_863)
);

CKINVDCx14_ASAP7_75t_R g864 ( 
.A(n_570),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_472),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_135),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_202),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_270),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_96),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_531),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_34),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_54),
.Y(n_872)
);

CKINVDCx14_ASAP7_75t_R g873 ( 
.A(n_241),
.Y(n_873)
);

BUFx2_ASAP7_75t_SL g874 ( 
.A(n_159),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_242),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_486),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_41),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_292),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_22),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_341),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_317),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_407),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_25),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_33),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_224),
.Y(n_885)
);

CKINVDCx16_ASAP7_75t_R g886 ( 
.A(n_253),
.Y(n_886)
);

BUFx5_ASAP7_75t_L g887 ( 
.A(n_259),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_418),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_34),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_184),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_296),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_482),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_334),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_1),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_445),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_347),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_130),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_87),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_4),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_226),
.Y(n_900)
);

CKINVDCx16_ASAP7_75t_R g901 ( 
.A(n_81),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_162),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_287),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_40),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_520),
.Y(n_905)
);

BUFx10_ASAP7_75t_L g906 ( 
.A(n_406),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_70),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_385),
.Y(n_908)
);

BUFx10_ASAP7_75t_L g909 ( 
.A(n_160),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_85),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_401),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_234),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_426),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_233),
.B(n_160),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_543),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_514),
.Y(n_916)
);

BUFx12f_ASAP7_75t_L g917 ( 
.A(n_816),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_724),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_918)
);

BUFx12f_ASAP7_75t_L g919 ( 
.A(n_656),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_736),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_580),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_580),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_816),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_736),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_724),
.B(n_3),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_579),
.B(n_5),
.Y(n_926)
);

OAI22x1_ASAP7_75t_SL g927 ( 
.A1(n_595),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_816),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_736),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_618),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_628),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_736),
.Y(n_932)
);

AND2x2_ASAP7_75t_SL g933 ( 
.A(n_676),
.B(n_464),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_736),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_736),
.Y(n_935)
);

BUFx8_ASAP7_75t_SL g936 ( 
.A(n_751),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_579),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_579),
.B(n_639),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_813),
.B(n_6),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_656),
.Y(n_940)
);

BUFx12f_ASAP7_75t_L g941 ( 
.A(n_656),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_736),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_813),
.B(n_9),
.Y(n_943)
);

OA21x2_ASAP7_75t_L g944 ( 
.A1(n_649),
.A2(n_468),
.B(n_467),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_649),
.A2(n_471),
.B(n_470),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_674),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_577),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_618),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_702),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_618),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_639),
.B(n_9),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_873),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_661),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_674),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_887),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_618),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_679),
.B(n_11),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_873),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_703),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_577),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_689),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_887),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_SL g963 ( 
.A1(n_595),
.A2(n_19),
.B1(n_14),
.B2(n_18),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_616),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_679),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_884),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_661),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_730),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_730),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_740),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_808),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_740),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_597),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_689),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_597),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_887),
.Y(n_976)
);

OA21x2_ASAP7_75t_L g977 ( 
.A1(n_683),
.A2(n_475),
.B(n_474),
.Y(n_977)
);

OA21x2_ASAP7_75t_L g978 ( 
.A1(n_683),
.A2(n_478),
.B(n_477),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_750),
.B(n_23),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_703),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_599),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_887),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_689),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_599),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_795),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_811),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_811),
.B(n_24),
.Y(n_987)
);

BUFx8_ASAP7_75t_L g988 ( 
.A(n_914),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_906),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_SL g990 ( 
.A1(n_606),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_833),
.B(n_29),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_897),
.B(n_29),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_887),
.B(n_575),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_903),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_703),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_886),
.B(n_30),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_903),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_887),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_627),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_901),
.B(n_31),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_575),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_703),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_870),
.B(n_32),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_575),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_870),
.B(n_33),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_766),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_SL g1007 ( 
.A1(n_606),
.A2(n_658),
.B1(n_666),
.B2(n_622),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_675),
.Y(n_1008)
);

CKINVDCx6p67_ASAP7_75t_R g1009 ( 
.A(n_919),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_926),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_928),
.B(n_817),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_923),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_926),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_924),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_924),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_946),
.B(n_699),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_923),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_951),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_929),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_964),
.B(n_966),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_921),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_964),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_921),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_923),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_936),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1008),
.B(n_602),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_929),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_946),
.B(n_699),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_992),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_966),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_946),
.B(n_838),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_938),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_932),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_931),
.B(n_838),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_932),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_975),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_925),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_934),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_921),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_975),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_934),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_935),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_931),
.B(n_845),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_981),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_981),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_935),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_974),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_931),
.B(n_845),
.Y(n_1048)
);

INVxp33_ASAP7_75t_L g1049 ( 
.A(n_984),
.Y(n_1049)
);

XOR2x2_ASAP7_75t_L g1050 ( 
.A(n_1007),
.B(n_691),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_942),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_942),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_984),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_955),
.Y(n_1054)
);

OAI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_918),
.A2(n_658),
.B1(n_666),
.B2(n_622),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1008),
.B(n_604),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_953),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_955),
.Y(n_1058)
);

AO21x2_ASAP7_75t_L g1059 ( 
.A1(n_945),
.A2(n_589),
.B(n_574),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_962),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_941),
.Y(n_1061)
);

CKINVDCx16_ASAP7_75t_R g1062 ( 
.A(n_917),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_946),
.B(n_575),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_L g1064 ( 
.A(n_1001),
.B(n_575),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_962),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_973),
.B(n_604),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_976),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_967),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_976),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_917),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_961),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_969),
.Y(n_1072)
);

NOR2x1p5_ASAP7_75t_L g1073 ( 
.A(n_989),
.B(n_607),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_970),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_949),
.B(n_607),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_971),
.B(n_648),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_972),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_982),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_982),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_998),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_994),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_SL g1082 ( 
.A(n_933),
.B(n_672),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_998),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1001),
.Y(n_1084)
);

INVx5_ASAP7_75t_L g1085 ( 
.A(n_921),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1004),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_954),
.B(n_575),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_997),
.B(n_611),
.Y(n_1088)
);

NOR2x1p5_ASAP7_75t_L g1089 ( 
.A(n_936),
.B(n_611),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1004),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_922),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_979),
.Y(n_1092)
);

INVx8_ASAP7_75t_L g1093 ( 
.A(n_954),
.Y(n_1093)
);

OAI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_952),
.A2(n_958),
.B1(n_986),
.B2(n_968),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_922),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_922),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_987),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_922),
.Y(n_1098)
);

BUFx10_ASAP7_75t_L g1099 ( 
.A(n_933),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_SL g1100 ( 
.A(n_939),
.B(n_672),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_947),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_940),
.Y(n_1102)
);

OR2x6_ASAP7_75t_L g1103 ( 
.A(n_990),
.B(n_874),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_937),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_999),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_991),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_960),
.B(n_612),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_930),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_SL g1109 ( 
.A(n_983),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_996),
.B(n_864),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_965),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_985),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_991),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1003),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1003),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_930),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_948),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_948),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_948),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_985),
.B(n_965),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1005),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_950),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_950),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_950),
.Y(n_1124)
);

AND2x6_ASAP7_75t_L g1125 ( 
.A(n_943),
.B(n_1005),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_957),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_944),
.Y(n_1127)
);

INVx5_ASAP7_75t_L g1128 ( 
.A(n_956),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_988),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_1000),
.Y(n_1130)
);

INVx8_ASAP7_75t_L g1131 ( 
.A(n_988),
.Y(n_1131)
);

INVx8_ASAP7_75t_L g1132 ( 
.A(n_993),
.Y(n_1132)
);

BUFx10_ASAP7_75t_L g1133 ( 
.A(n_956),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_944),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1006),
.B(n_614),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_959),
.B(n_660),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_980),
.B(n_662),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_980),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_977),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_980),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_977),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_963),
.B(n_906),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_995),
.B(n_700),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_978),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1006),
.B(n_614),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_995),
.B(n_704),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_995),
.B(n_708),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1002),
.B(n_621),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1002),
.B(n_721),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_978),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1002),
.B(n_723),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1006),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_927),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_945),
.A2(n_793),
.B(n_738),
.Y(n_1154)
);

BUFx10_ASAP7_75t_L g1155 ( 
.A(n_938),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_964),
.B(n_624),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_920),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1092),
.B(n_620),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1057),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1097),
.B(n_620),
.Y(n_1160)
);

AOI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1094),
.A2(n_755),
.B1(n_867),
.B2(n_866),
.C(n_827),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1094),
.A2(n_715),
.B1(n_767),
.B2(n_692),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1022),
.B(n_909),
.Y(n_1163)
);

NAND2xp33_ASAP7_75t_SL g1164 ( 
.A(n_1049),
.B(n_692),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1106),
.B(n_865),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1113),
.B(n_865),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1101),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1101),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1011),
.B(n_876),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1100),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1126),
.B(n_876),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1068),
.Y(n_1172)
);

INVx8_ASAP7_75t_L g1173 ( 
.A(n_1131),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1114),
.B(n_916),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1115),
.B(n_592),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1072),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1102),
.B(n_578),
.Y(n_1177)
);

BUFx5_ASAP7_75t_L g1178 ( 
.A(n_1144),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1066),
.B(n_868),
.C(n_867),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1144),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1032),
.B(n_625),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_L g1182 ( 
.A(n_1055),
.B(n_711),
.C(n_667),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1121),
.B(n_613),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1074),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1077),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1049),
.B(n_696),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1020),
.B(n_909),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1018),
.B(n_701),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1018),
.B(n_752),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1029),
.B(n_769),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1029),
.B(n_769),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1155),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_1131),
.Y(n_1193)
);

AO221x1_ASAP7_75t_L g1194 ( 
.A1(n_1055),
.A2(n_1082),
.B1(n_1061),
.B2(n_1071),
.C(n_1099),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1026),
.B(n_636),
.Y(n_1195)
);

BUFx12f_ASAP7_75t_L g1196 ( 
.A(n_1025),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1156),
.B(n_909),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1130),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1056),
.B(n_637),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1131),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1081),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1093),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1110),
.B(n_690),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1062),
.B(n_868),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1009),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1107),
.B(n_694),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1013),
.B(n_737),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1112),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1070),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1134),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1010),
.B(n_761),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1047),
.B(n_762),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1112),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1105),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_SL g1215 ( 
.A(n_1129),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1104),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_1037),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1036),
.B(n_771),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1135),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1040),
.B(n_782),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1044),
.B(n_794),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1145),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1148),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1088),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1109),
.Y(n_1225)
);

NAND2xp33_ASAP7_75t_L g1226 ( 
.A(n_1132),
.B(n_802),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1045),
.B(n_806),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1053),
.A2(n_767),
.B1(n_784),
.B2(n_715),
.Y(n_1228)
);

AOI22x1_ASAP7_75t_L g1229 ( 
.A1(n_1141),
.A2(n_844),
.B1(n_825),
.B2(n_840),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1075),
.B(n_809),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1084),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1076),
.B(n_819),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1142),
.B(n_869),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1132),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1125),
.B(n_839),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1086),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1073),
.B(n_784),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_SL g1238 ( 
.A(n_1153),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1125),
.B(n_852),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1012),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1064),
.A2(n_581),
.B(n_583),
.C(n_573),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1090),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1136),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1133),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1109),
.B(n_832),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1125),
.B(n_869),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1034),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1017),
.B(n_1024),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1133),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1132),
.A2(n_821),
.B1(n_809),
.B2(n_584),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1099),
.A2(n_861),
.B1(n_804),
.B2(n_871),
.Y(n_1251)
);

AND2x6_ASAP7_75t_SL g1252 ( 
.A(n_1103),
.B(n_586),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1120),
.B(n_915),
.Y(n_1253)
);

AO221x1_ASAP7_75t_L g1254 ( 
.A1(n_1127),
.A2(n_751),
.B1(n_861),
.B2(n_804),
.C(n_773),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1136),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1093),
.B(n_871),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_1043),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_1048),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1111),
.B(n_856),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1064),
.B(n_877),
.C(n_585),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1059),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1048),
.B(n_905),
.Y(n_1262)
);

NAND2xp33_ASAP7_75t_L g1263 ( 
.A(n_1127),
.B(n_863),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1137),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1014),
.A2(n_821),
.B1(n_588),
.B2(n_596),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1016),
.B(n_892),
.Y(n_1266)
);

NOR3xp33_ASAP7_75t_L g1267 ( 
.A(n_1016),
.B(n_659),
.C(n_582),
.Y(n_1267)
);

BUFx5_ASAP7_75t_L g1268 ( 
.A(n_1138),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1015),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1157),
.B(n_587),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1137),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_L g1272 ( 
.A(n_1015),
.B(n_593),
.C(n_590),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1089),
.B(n_594),
.Y(n_1273)
);

INVxp67_ASAP7_75t_L g1274 ( 
.A(n_1103),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1103),
.A2(n_900),
.B1(n_904),
.B2(n_899),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1028),
.B(n_766),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1031),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1019),
.B(n_598),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1031),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_1027),
.B(n_632),
.C(n_600),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1139),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1033),
.B(n_635),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1035),
.B(n_640),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1035),
.B(n_790),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1038),
.B(n_576),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1038),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1041),
.B(n_644),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1139),
.B(n_647),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1042),
.B(n_790),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1046),
.B(n_576),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1046),
.B(n_610),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1150),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1149),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1051),
.B(n_610),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1149),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1052),
.B(n_617),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1154),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1063),
.A2(n_745),
.B1(n_773),
.B2(n_731),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1154),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1052),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1054),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1058),
.B(n_617),
.Y(n_1302)
);

NOR3xp33_ASAP7_75t_L g1303 ( 
.A(n_1087),
.B(n_765),
.C(n_753),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1087),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1060),
.B(n_629),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1065),
.B(n_629),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1065),
.B(n_638),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1067),
.B(n_651),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1050),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1069),
.B(n_638),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1078),
.B(n_652),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1079),
.A2(n_601),
.B1(n_603),
.B2(n_591),
.Y(n_1312)
);

NAND2x1_ASAP7_75t_L g1313 ( 
.A(n_1079),
.B(n_643),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1080),
.A2(n_608),
.B1(n_609),
.B2(n_605),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1083),
.B(n_653),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1143),
.B(n_654),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1143),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1146),
.B(n_643),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1147),
.Y(n_1319)
);

NOR2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1140),
.B(n_663),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1108),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1151),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1039),
.B(n_650),
.Y(n_1323)
);

AO221x1_ASAP7_75t_L g1324 ( 
.A1(n_1108),
.A2(n_786),
.B1(n_792),
.B2(n_745),
.C(n_731),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1039),
.B(n_650),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1039),
.B(n_669),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1039),
.B(n_812),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1085),
.B(n_670),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1116),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1085),
.B(n_671),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1085),
.B(n_859),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1128),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1128),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1085),
.B(n_670),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1128),
.B(n_685),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1091),
.B(n_685),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1021),
.B(n_677),
.Y(n_1337)
);

NOR2x1p5_ASAP7_75t_L g1338 ( 
.A(n_1117),
.B(n_686),
.Y(n_1338)
);

NAND2x1_ASAP7_75t_L g1339 ( 
.A(n_1118),
.B(n_713),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1091),
.B(n_713),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1095),
.B(n_718),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1095),
.B(n_718),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1119),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1119),
.A2(n_619),
.B1(n_623),
.B2(n_615),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1096),
.B(n_722),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1122),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1023),
.B(n_687),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1096),
.B(n_722),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1023),
.B(n_693),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1023),
.B(n_859),
.Y(n_1350)
);

AND2x4_ASAP7_75t_SL g1351 ( 
.A(n_1123),
.B(n_786),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1123),
.A2(n_698),
.B1(n_705),
.B2(n_695),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1124),
.A2(n_894),
.B1(n_895),
.B2(n_893),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1098),
.B(n_789),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1098),
.B(n_789),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1301),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1158),
.B(n_712),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1173),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1198),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1202),
.B(n_714),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1202),
.B(n_720),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1198),
.B(n_792),
.Y(n_1362)
);

BUFx8_ASAP7_75t_L g1363 ( 
.A(n_1215),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1159),
.Y(n_1364)
);

CKINVDCx8_ASAP7_75t_R g1365 ( 
.A(n_1173),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1158),
.B(n_727),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1160),
.B(n_729),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1193),
.B(n_716),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1286),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1160),
.B(n_1224),
.Y(n_1370)
);

OAI21xp33_ASAP7_75t_L g1371 ( 
.A1(n_1163),
.A2(n_739),
.B(n_735),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1186),
.B(n_741),
.Y(n_1372)
);

AOI21xp33_ASAP7_75t_L g1373 ( 
.A1(n_1246),
.A2(n_746),
.B(n_742),
.Y(n_1373)
);

O2A1O1Ixp5_ASAP7_75t_L g1374 ( 
.A1(n_1261),
.A2(n_882),
.B(n_896),
.C(n_824),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1217),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1300),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1161),
.A2(n_890),
.B1(n_831),
.B2(n_630),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1233),
.A2(n_763),
.B1(n_764),
.B2(n_758),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1172),
.Y(n_1379)
);

OR2x6_ASAP7_75t_L g1380 ( 
.A(n_1200),
.B(n_754),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1176),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1241),
.A2(n_631),
.B(n_633),
.C(n_626),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1214),
.Y(n_1383)
);

NOR3xp33_ASAP7_75t_L g1384 ( 
.A(n_1162),
.B(n_818),
.C(n_798),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1165),
.B(n_768),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1184),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1166),
.B(n_774),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1166),
.B(n_775),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1205),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1197),
.A2(n_777),
.B1(n_779),
.B2(n_776),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1174),
.B(n_781),
.Y(n_1391)
);

OAI21xp33_ASAP7_75t_L g1392 ( 
.A1(n_1187),
.A2(n_785),
.B(n_783),
.Y(n_1392)
);

AOI21xp33_ASAP7_75t_L g1393 ( 
.A1(n_1274),
.A2(n_796),
.B(n_791),
.Y(n_1393)
);

NOR3xp33_ASAP7_75t_L g1394 ( 
.A(n_1162),
.B(n_1164),
.C(n_1298),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1185),
.B(n_797),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1288),
.A2(n_665),
.B(n_642),
.Y(n_1396)
);

NAND2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1234),
.B(n_824),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1201),
.B(n_799),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1333),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1192),
.B(n_800),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1175),
.A2(n_890),
.B1(n_831),
.B2(n_641),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1175),
.A2(n_1183),
.B1(n_1216),
.B2(n_1285),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1169),
.A2(n_805),
.B1(n_807),
.B2(n_803),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1182),
.A2(n_645),
.B(n_646),
.C(n_634),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1188),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1196),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1188),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1167),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1228),
.B(n_850),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1219),
.A2(n_778),
.B(n_744),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1222),
.A2(n_657),
.B(n_655),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_L g1412 ( 
.A(n_1178),
.B(n_823),
.Y(n_1412)
);

AOI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1170),
.A2(n_828),
.B(n_826),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1168),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1208),
.Y(n_1415)
);

OR2x6_ASAP7_75t_SL g1416 ( 
.A(n_1298),
.B(n_829),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1320),
.B(n_801),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1230),
.B(n_830),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1209),
.B(n_834),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1204),
.B(n_835),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1285),
.A2(n_668),
.B1(n_673),
.B2(n_664),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1351),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1213),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1290),
.A2(n_680),
.B1(n_681),
.B2(n_678),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1189),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1190),
.A2(n_1152),
.B(n_684),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1251),
.B(n_1275),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1223),
.A2(n_688),
.B(n_697),
.C(n_682),
.Y(n_1428)
);

OAI321xp33_ASAP7_75t_L g1429 ( 
.A1(n_1190),
.A2(n_710),
.A3(n_707),
.B1(n_717),
.B2(n_709),
.C(n_706),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1324),
.B(n_837),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1191),
.A2(n_725),
.B(n_719),
.Y(n_1431)
);

O2A1O1Ixp5_ASAP7_75t_L g1432 ( 
.A1(n_1262),
.A2(n_913),
.B(n_896),
.C(n_728),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1225),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1247),
.A2(n_732),
.B1(n_733),
.B2(n_726),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1290),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1256),
.B(n_842),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1180),
.B(n_847),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1304),
.A2(n_1199),
.B(n_1195),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1243),
.A2(n_743),
.B(n_747),
.C(n_734),
.Y(n_1439)
);

NOR3xp33_ASAP7_75t_L g1440 ( 
.A(n_1309),
.B(n_853),
.C(n_849),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1257),
.A2(n_1258),
.B(n_1255),
.Y(n_1441)
);

AND2x2_ASAP7_75t_SL g1442 ( 
.A(n_1237),
.B(n_913),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1281),
.A2(n_749),
.B(n_748),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1180),
.B(n_858),
.Y(n_1444)
);

AO21x1_ASAP7_75t_L g1445 ( 
.A1(n_1291),
.A2(n_757),
.B(n_756),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1281),
.A2(n_760),
.B(n_759),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1231),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1308),
.B(n_862),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1311),
.B(n_881),
.Y(n_1449)
);

AO21x1_ASAP7_75t_L g1450 ( 
.A1(n_1291),
.A2(n_772),
.B(n_770),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1264),
.A2(n_787),
.B(n_788),
.C(n_780),
.Y(n_1451)
);

NOR2x2_ASAP7_75t_L g1452 ( 
.A(n_1254),
.B(n_907),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1271),
.A2(n_814),
.B(n_810),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1315),
.B(n_883),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1292),
.A2(n_820),
.B(n_815),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1203),
.B(n_889),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1232),
.B(n_910),
.Y(n_1457)
);

INVx11_ASAP7_75t_L g1458 ( 
.A(n_1215),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1211),
.A2(n_836),
.B(n_822),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1293),
.A2(n_843),
.B(n_841),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1218),
.B(n_885),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1294),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1210),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1270),
.B(n_846),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1295),
.A2(n_851),
.B(n_854),
.C(n_848),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1338),
.B(n_855),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1235),
.A2(n_1239),
.B(n_1206),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1322),
.A2(n_860),
.B1(n_872),
.B2(n_857),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1278),
.B(n_875),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1220),
.B(n_879),
.Y(n_1470)
);

AOI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1179),
.A2(n_888),
.B(n_880),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1210),
.A2(n_898),
.B(n_891),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1282),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1210),
.A2(n_908),
.B(n_902),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1283),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1287),
.B(n_911),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1194),
.B(n_1273),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1236),
.A2(n_912),
.B(n_878),
.Y(n_1478)
);

INVx5_ASAP7_75t_L g1479 ( 
.A(n_1333),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1296),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1177),
.B(n_1245),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1303),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1267),
.B(n_36),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1212),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1207),
.A2(n_484),
.B(n_479),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1302),
.Y(n_1486)
);

NOR3xp33_ASAP7_75t_L g1487 ( 
.A(n_1221),
.B(n_1227),
.C(n_1272),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1250),
.B(n_1171),
.Y(n_1488)
);

OAI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1242),
.A2(n_487),
.B(n_485),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1352),
.B(n_37),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1353),
.B(n_38),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1312),
.B(n_39),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1314),
.B(n_41),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1316),
.B(n_1265),
.Y(n_1494)
);

NOR2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1238),
.B(n_42),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1302),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1305),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1305),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1244),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1181),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1259),
.B(n_43),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1260),
.B(n_43),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1306),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1299),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1249),
.B(n_46),
.Y(n_1505)
);

AO21x1_ASAP7_75t_L g1506 ( 
.A1(n_1306),
.A2(n_48),
.B(n_49),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1269),
.A2(n_503),
.B(n_501),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_R g1508 ( 
.A(n_1238),
.B(n_48),
.Y(n_1508)
);

INVx11_ASAP7_75t_L g1509 ( 
.A(n_1252),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1318),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1307),
.Y(n_1511)
);

NAND2xp33_ASAP7_75t_L g1512 ( 
.A(n_1229),
.B(n_506),
.Y(n_1512)
);

BUFx4f_ASAP7_75t_L g1513 ( 
.A(n_1277),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1307),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1279),
.B(n_51),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1344),
.B(n_52),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1310),
.B(n_53),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1323),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1240),
.A2(n_510),
.B(n_509),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1280),
.B(n_56),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1253),
.B(n_56),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1226),
.B(n_57),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1266),
.B(n_57),
.Y(n_1523)
);

AOI21xp33_ASAP7_75t_L g1524 ( 
.A1(n_1248),
.A2(n_59),
.B(n_60),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1332),
.B(n_61),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1318),
.A2(n_513),
.B(n_512),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1313),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1321),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1317),
.A2(n_64),
.B1(n_61),
.B2(n_62),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1323),
.Y(n_1530)
);

BUFx4f_ASAP7_75t_L g1531 ( 
.A(n_1319),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1336),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1325),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1326),
.B(n_65),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1325),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1339),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1337),
.B(n_66),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1336),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1330),
.B(n_67),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1328),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1347),
.B(n_69),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1276),
.A2(n_519),
.B(n_518),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1328),
.Y(n_1543)
);

NAND2xp33_ASAP7_75t_L g1544 ( 
.A(n_1268),
.B(n_523),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1349),
.B(n_69),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1334),
.B(n_70),
.Y(n_1546)
);

AOI21xp33_ASAP7_75t_L g1547 ( 
.A1(n_1335),
.A2(n_71),
.B(n_72),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1340),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1335),
.B(n_73),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1329),
.A2(n_536),
.B(n_532),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1340),
.B(n_75),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1341),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1341),
.B(n_77),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1321),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1342),
.Y(n_1555)
);

OAI321xp33_ASAP7_75t_L g1556 ( 
.A1(n_1345),
.A2(n_83),
.A3(n_85),
.B1(n_79),
.B2(n_82),
.C(n_84),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1327),
.B(n_79),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1345),
.A2(n_1348),
.B1(n_1355),
.B2(n_1354),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1348),
.B(n_84),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1354),
.B(n_86),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1355),
.A2(n_538),
.B(n_537),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1331),
.B(n_86),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1268),
.B(n_87),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1268),
.B(n_88),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1346),
.A2(n_540),
.B(n_539),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1284),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1289),
.A2(n_545),
.B(n_542),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1268),
.B(n_89),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1343),
.B(n_90),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1268),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1350),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1297),
.A2(n_552),
.B(n_551),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1241),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1158),
.B(n_95),
.Y(n_1574)
);

O2A1O1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1217),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1263),
.A2(n_554),
.B(n_553),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1159),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1158),
.B(n_98),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1158),
.B(n_99),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1198),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1205),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1159),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1159),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1427),
.B(n_1370),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1580),
.B(n_101),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1364),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1511),
.B(n_1402),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_L g1588 ( 
.A1(n_1420),
.A2(n_102),
.B(n_103),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1438),
.A2(n_103),
.B(n_104),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1467),
.A2(n_105),
.B(n_106),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_R g1591 ( 
.A(n_1406),
.B(n_105),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1416),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1402),
.B(n_107),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1362),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_SL g1595 ( 
.A1(n_1441),
.A2(n_108),
.B(n_109),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1365),
.Y(n_1596)
);

AND2x6_ASAP7_75t_L g1597 ( 
.A(n_1504),
.B(n_111),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1358),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1379),
.Y(n_1599)
);

OA21x2_ASAP7_75t_L g1600 ( 
.A1(n_1572),
.A2(n_113),
.B(n_114),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1363),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1475),
.B(n_113),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1381),
.B(n_114),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1386),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1441),
.B(n_119),
.Y(n_1605)
);

BUFx12f_ASAP7_75t_L g1606 ( 
.A(n_1363),
.Y(n_1606)
);

BUFx4f_ASAP7_75t_L g1607 ( 
.A(n_1442),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1401),
.B(n_1375),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_SL g1609 ( 
.A(n_1581),
.B(n_120),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1405),
.A2(n_120),
.B(n_121),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1401),
.B(n_122),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1577),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1435),
.A2(n_128),
.B(n_125),
.C(n_127),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1384),
.B(n_127),
.Y(n_1614)
);

AND3x2_ASAP7_75t_L g1615 ( 
.A(n_1394),
.B(n_128),
.C(n_129),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1407),
.A2(n_129),
.B(n_130),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1425),
.A2(n_131),
.B(n_132),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1582),
.B(n_131),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1583),
.B(n_133),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1458),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1480),
.B(n_139),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1486),
.B(n_140),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1383),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_SL g1624 ( 
.A(n_1389),
.B(n_141),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1496),
.B(n_142),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1497),
.A2(n_146),
.B(n_143),
.C(n_144),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1498),
.B(n_148),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1422),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1514),
.B(n_149),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1453),
.B(n_151),
.Y(n_1630)
);

NOR2x1_ASAP7_75t_L g1631 ( 
.A(n_1495),
.B(n_152),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1525),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1494),
.A2(n_154),
.B(n_155),
.Y(n_1633)
);

BUFx4f_ASAP7_75t_L g1634 ( 
.A(n_1523),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1453),
.B(n_156),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1479),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1460),
.B(n_157),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1481),
.B(n_158),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1484),
.B(n_159),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1489),
.A2(n_161),
.B(n_162),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1489),
.A2(n_163),
.B(n_165),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1479),
.B(n_166),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1479),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1487),
.B(n_166),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1507),
.A2(n_167),
.B(n_168),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1558),
.A2(n_167),
.B(n_168),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1555),
.A2(n_169),
.B(n_170),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1554),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1554),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1447),
.Y(n_1650)
);

INVx5_ASAP7_75t_L g1651 ( 
.A(n_1463),
.Y(n_1651)
);

OAI22x1_ASAP7_75t_L g1652 ( 
.A1(n_1466),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1433),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1460),
.B(n_175),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1525),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1478),
.A2(n_180),
.B(n_181),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1478),
.A2(n_184),
.B(n_185),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1409),
.B(n_189),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1488),
.A2(n_190),
.B(n_191),
.Y(n_1659)
);

AOI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1419),
.A2(n_191),
.B(n_192),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1500),
.B(n_195),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1377),
.B(n_198),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1411),
.B(n_1473),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1431),
.A2(n_198),
.B(n_199),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1543),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1463),
.B(n_201),
.Y(n_1666)
);

AO31x2_ASAP7_75t_L g1667 ( 
.A1(n_1506),
.A2(n_203),
.A3(n_201),
.B(n_202),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1357),
.A2(n_203),
.B(n_204),
.Y(n_1668)
);

AO31x2_ASAP7_75t_L g1669 ( 
.A1(n_1445),
.A2(n_206),
.A3(n_204),
.B(n_205),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1477),
.B(n_207),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1366),
.B(n_1367),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1428),
.B(n_209),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1439),
.B(n_210),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1518),
.A2(n_210),
.B(n_211),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1523),
.Y(n_1675)
);

INVx2_ASAP7_75t_SL g1676 ( 
.A(n_1513),
.Y(n_1676)
);

AO21x1_ASAP7_75t_L g1677 ( 
.A1(n_1561),
.A2(n_212),
.B(n_213),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1451),
.B(n_212),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1465),
.B(n_214),
.Y(n_1679)
);

AO31x2_ASAP7_75t_L g1680 ( 
.A1(n_1450),
.A2(n_217),
.A3(n_215),
.B(n_216),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1528),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1568),
.B(n_217),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1385),
.B(n_218),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1563),
.A2(n_218),
.B(n_220),
.Y(n_1684)
);

NOR2x1_ASAP7_75t_L g1685 ( 
.A(n_1483),
.B(n_221),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1526),
.A2(n_1396),
.B(n_1485),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1508),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1534),
.B(n_223),
.C(n_225),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1369),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1492),
.Y(n_1690)
);

AO21x1_ASAP7_75t_L g1691 ( 
.A1(n_1526),
.A2(n_227),
.B(n_228),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1503),
.A2(n_230),
.B(n_227),
.C(n_229),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1391),
.B(n_232),
.Y(n_1694)
);

XNOR2xp5_ASAP7_75t_L g1695 ( 
.A(n_1468),
.B(n_236),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_SL g1696 ( 
.A1(n_1564),
.A2(n_238),
.B(n_239),
.Y(n_1696)
);

O2A1O1Ixp33_ASAP7_75t_L g1697 ( 
.A1(n_1382),
.A2(n_244),
.B(n_240),
.C(n_243),
.Y(n_1697)
);

AO21x1_ASAP7_75t_L g1698 ( 
.A1(n_1396),
.A2(n_244),
.B(n_245),
.Y(n_1698)
);

AOI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1539),
.A2(n_245),
.B(n_246),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1390),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1509),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1418),
.B(n_251),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1493),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1378),
.B(n_252),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1574),
.A2(n_255),
.B(n_257),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1552),
.A2(n_259),
.B(n_257),
.C(n_258),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1573),
.A2(n_262),
.B(n_260),
.C(n_261),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1459),
.B(n_263),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_R g1709 ( 
.A(n_1430),
.B(n_265),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1575),
.A2(n_267),
.B(n_268),
.C(n_271),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1530),
.A2(n_272),
.B(n_273),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1404),
.B(n_1372),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_L g1713 ( 
.A1(n_1510),
.A2(n_273),
.B(n_274),
.C(n_275),
.Y(n_1713)
);

AO21x1_ASAP7_75t_L g1714 ( 
.A1(n_1544),
.A2(n_274),
.B(n_276),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1569),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1578),
.A2(n_277),
.B(n_278),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1579),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1535),
.A2(n_279),
.B(n_282),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1512),
.A2(n_284),
.B(n_285),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1356),
.Y(n_1720)
);

AO31x2_ASAP7_75t_L g1721 ( 
.A1(n_1532),
.A2(n_285),
.A3(n_286),
.B(n_287),
.Y(n_1721)
);

BUFx10_ASAP7_75t_L g1722 ( 
.A(n_1545),
.Y(n_1722)
);

AO21x1_ASAP7_75t_L g1723 ( 
.A1(n_1519),
.A2(n_288),
.B(n_289),
.Y(n_1723)
);

OAI21xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1546),
.A2(n_288),
.B(n_290),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1426),
.A2(n_293),
.B(n_294),
.Y(n_1725)
);

CKINVDCx6p67_ASAP7_75t_R g1726 ( 
.A(n_1380),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1403),
.B(n_1490),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1464),
.B(n_1469),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1397),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1491),
.B(n_297),
.Y(n_1730)
);

A2O1A1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1570),
.A2(n_1520),
.B(n_1476),
.C(n_1429),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1516),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1432),
.A2(n_298),
.B(n_299),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1499),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1429),
.A2(n_300),
.B(n_301),
.C(n_304),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_1393),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1443),
.A2(n_304),
.B(n_305),
.Y(n_1737)
);

AOI21xp33_ASAP7_75t_L g1738 ( 
.A1(n_1457),
.A2(n_306),
.B(n_307),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1499),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1421),
.B(n_309),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1533),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1446),
.A2(n_310),
.B(n_311),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1424),
.B(n_312),
.Y(n_1743)
);

OAI21x1_ASAP7_75t_SL g1744 ( 
.A1(n_1515),
.A2(n_312),
.B(n_313),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1395),
.Y(n_1745)
);

AO31x2_ASAP7_75t_L g1746 ( 
.A1(n_1532),
.A2(n_313),
.A3(n_314),
.B(n_315),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1556),
.A2(n_314),
.B(n_315),
.C(n_316),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1398),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1461),
.B(n_316),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1470),
.B(n_317),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1553),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1434),
.B(n_318),
.Y(n_1752)
);

AO31x2_ASAP7_75t_L g1753 ( 
.A1(n_1538),
.A2(n_318),
.A3(n_319),
.B(n_320),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1360),
.B(n_321),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1412),
.A2(n_321),
.B(n_322),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1540),
.Y(n_1756)
);

CKINVDCx11_ASAP7_75t_R g1757 ( 
.A(n_1380),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1399),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1392),
.B(n_323),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1538),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1399),
.Y(n_1761)
);

OAI21x1_ASAP7_75t_SL g1762 ( 
.A1(n_1548),
.A2(n_325),
.B(n_326),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1456),
.B(n_326),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1436),
.A2(n_327),
.B(n_328),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1455),
.A2(n_328),
.B(n_329),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1448),
.A2(n_329),
.B(n_330),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1371),
.B(n_331),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1536),
.Y(n_1768)
);

BUFx3_ASAP7_75t_L g1769 ( 
.A(n_1513),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1545),
.A2(n_332),
.B(n_333),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1449),
.A2(n_334),
.B(n_335),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1361),
.B(n_339),
.Y(n_1772)
);

INVxp33_ASAP7_75t_SL g1773 ( 
.A(n_1440),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1454),
.A2(n_339),
.B(n_340),
.Y(n_1774)
);

OAI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1472),
.A2(n_340),
.B(n_341),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1471),
.B(n_342),
.Y(n_1776)
);

NOR2x1_ASAP7_75t_SL g1777 ( 
.A(n_1548),
.B(n_344),
.Y(n_1777)
);

A2O1A1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1556),
.A2(n_345),
.B(n_346),
.C(n_348),
.Y(n_1778)
);

AND2x6_ASAP7_75t_L g1779 ( 
.A(n_1527),
.B(n_1376),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1408),
.Y(n_1780)
);

OAI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1474),
.A2(n_349),
.B(n_350),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1521),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1482),
.A2(n_354),
.B(n_355),
.C(n_356),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1517),
.A2(n_354),
.B(n_356),
.Y(n_1784)
);

OA21x2_ASAP7_75t_L g1785 ( 
.A1(n_1410),
.A2(n_1565),
.B(n_1550),
.Y(n_1785)
);

A2O1A1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1547),
.A2(n_362),
.B(n_363),
.C(n_364),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1551),
.A2(n_365),
.B(n_366),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1417),
.B(n_367),
.Y(n_1788)
);

BUFx4f_ASAP7_75t_SL g1789 ( 
.A(n_1437),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1531),
.A2(n_368),
.B(n_369),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1380),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1576),
.A2(n_368),
.B(n_370),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1414),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1415),
.Y(n_1794)
);

AO21x1_ASAP7_75t_L g1795 ( 
.A1(n_1537),
.A2(n_370),
.B(n_371),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1373),
.B(n_371),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1423),
.B(n_373),
.Y(n_1797)
);

AOI21xp33_ASAP7_75t_L g1798 ( 
.A1(n_1400),
.A2(n_1444),
.B(n_1501),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1531),
.A2(n_374),
.B(n_375),
.Y(n_1799)
);

BUFx12f_ASAP7_75t_L g1800 ( 
.A(n_1368),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1571),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1571),
.Y(n_1802)
);

BUFx12f_ASAP7_75t_L g1803 ( 
.A(n_1368),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1417),
.B(n_377),
.Y(n_1804)
);

AO21x1_ASAP7_75t_L g1805 ( 
.A1(n_1541),
.A2(n_377),
.B(n_378),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1505),
.B(n_378),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1413),
.B(n_1524),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_SL g1808 ( 
.A1(n_1522),
.A2(n_379),
.B(n_380),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1559),
.B(n_381),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1549),
.B(n_383),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1560),
.Y(n_1811)
);

BUFx10_ASAP7_75t_L g1812 ( 
.A(n_1557),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1502),
.B(n_384),
.Y(n_1813)
);

AO22x1_ASAP7_75t_L g1814 ( 
.A1(n_1452),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_1814)
);

BUFx8_ASAP7_75t_L g1815 ( 
.A(n_1529),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1562),
.B(n_386),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1566),
.B(n_387),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1542),
.A2(n_388),
.B(n_389),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1567),
.B(n_388),
.Y(n_1819)
);

AO31x2_ASAP7_75t_L g1820 ( 
.A1(n_1506),
.A2(n_390),
.A3(n_391),
.B(n_392),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1370),
.B(n_392),
.Y(n_1821)
);

OAI21x1_ASAP7_75t_SL g1822 ( 
.A1(n_1441),
.A2(n_394),
.B(n_395),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1370),
.A2(n_394),
.B(n_395),
.Y(n_1823)
);

AOI21xp33_ASAP7_75t_L g1824 ( 
.A1(n_1420),
.A2(n_396),
.B(n_397),
.Y(n_1824)
);

INVx2_ASAP7_75t_SL g1825 ( 
.A(n_1359),
.Y(n_1825)
);

A2O1A1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1370),
.A2(n_399),
.B(n_400),
.C(n_402),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1374),
.A2(n_400),
.B(n_402),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1365),
.Y(n_1828)
);

O2A1O1Ixp5_ASAP7_75t_L g1829 ( 
.A1(n_1396),
.A2(n_405),
.B(n_406),
.C(n_407),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1374),
.A2(n_408),
.B(n_409),
.Y(n_1830)
);

AOI221x1_ASAP7_75t_L g1831 ( 
.A1(n_1396),
.A2(n_408),
.B1(n_409),
.B2(n_410),
.C(n_411),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1359),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1394),
.A2(n_413),
.B1(n_415),
.B2(n_416),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_SL g1834 ( 
.A(n_1365),
.B(n_413),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1370),
.B(n_417),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1370),
.A2(n_421),
.B(n_422),
.Y(n_1836)
);

A2O1A1Ixp33_ASAP7_75t_L g1837 ( 
.A1(n_1370),
.A2(n_422),
.B(n_423),
.C(n_424),
.Y(n_1837)
);

INVx1_ASAP7_75t_SL g1838 ( 
.A(n_1359),
.Y(n_1838)
);

A2O1A1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1370),
.A2(n_423),
.B(n_424),
.C(n_425),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1370),
.B(n_426),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1370),
.A2(n_428),
.B(n_429),
.Y(n_1841)
);

NAND2x1p5_ASAP7_75t_L g1842 ( 
.A(n_1358),
.B(n_430),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1402),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1370),
.B(n_434),
.Y(n_1844)
);

A2O1A1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1370),
.A2(n_435),
.B(n_436),
.C(n_437),
.Y(n_1845)
);

AO31x2_ASAP7_75t_L g1846 ( 
.A1(n_1506),
.A2(n_435),
.A3(n_437),
.B(n_439),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1370),
.A2(n_440),
.B(n_441),
.Y(n_1847)
);

A2O1A1Ixp33_ASAP7_75t_L g1848 ( 
.A1(n_1370),
.A2(n_440),
.B(n_441),
.C(n_442),
.Y(n_1848)
);

NOR2x1_ASAP7_75t_L g1849 ( 
.A(n_1406),
.B(n_443),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1359),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1370),
.B(n_444),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1402),
.A2(n_444),
.B(n_446),
.Y(n_1852)
);

NAND2x1_ASAP7_75t_L g1853 ( 
.A(n_1528),
.B(n_447),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1427),
.B(n_448),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1359),
.B(n_448),
.Y(n_1855)
);

A2O1A1Ixp33_ASAP7_75t_L g1856 ( 
.A1(n_1370),
.A2(n_452),
.B(n_453),
.C(n_454),
.Y(n_1856)
);

BUFx12f_ASAP7_75t_L g1857 ( 
.A(n_1363),
.Y(n_1857)
);

A2O1A1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1370),
.A2(n_453),
.B(n_454),
.C(n_455),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1364),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1370),
.B(n_455),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1370),
.B(n_456),
.Y(n_1861)
);

A2O1A1Ixp33_ASAP7_75t_SL g1862 ( 
.A1(n_1396),
.A2(n_457),
.B(n_458),
.C(n_459),
.Y(n_1862)
);

INVx6_ASAP7_75t_L g1863 ( 
.A(n_1363),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1370),
.B(n_460),
.Y(n_1864)
);

A2O1A1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1370),
.A2(n_461),
.B(n_462),
.C(n_1438),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1370),
.B(n_1580),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1427),
.B(n_1099),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1370),
.B(n_1580),
.Y(n_1868)
);

OAI21xp33_ASAP7_75t_L g1869 ( 
.A1(n_1370),
.A2(n_1030),
.B(n_1022),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1370),
.B(n_1359),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1359),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1402),
.A2(n_1511),
.B1(n_1370),
.B2(n_1462),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1370),
.B(n_1580),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1359),
.B(n_1580),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1363),
.Y(n_1875)
);

NOR2xp67_ASAP7_75t_L g1876 ( 
.A(n_1580),
.B(n_1070),
.Y(n_1876)
);

BUFx8_ASAP7_75t_L g1877 ( 
.A(n_1359),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1650),
.Y(n_1878)
);

OR2x6_ASAP7_75t_L g1879 ( 
.A(n_1606),
.B(n_1857),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1586),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1865),
.B(n_1706),
.C(n_1692),
.Y(n_1881)
);

AO21x2_ASAP7_75t_L g1882 ( 
.A1(n_1590),
.A2(n_1830),
.B(n_1827),
.Y(n_1882)
);

INVx2_ASAP7_75t_SL g1883 ( 
.A(n_1606),
.Y(n_1883)
);

BUFx2_ASAP7_75t_L g1884 ( 
.A(n_1877),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1870),
.B(n_1584),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1599),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1838),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1877),
.Y(n_1888)
);

BUFx2_ASAP7_75t_SL g1889 ( 
.A(n_1653),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1681),
.Y(n_1890)
);

OAI21x1_ASAP7_75t_SL g1891 ( 
.A1(n_1872),
.A2(n_1587),
.B(n_1777),
.Y(n_1891)
);

BUFx8_ASAP7_75t_SL g1892 ( 
.A(n_1857),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1604),
.Y(n_1893)
);

NAND3xp33_ASAP7_75t_L g1894 ( 
.A(n_1865),
.B(n_1706),
.C(n_1692),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1870),
.B(n_1675),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1612),
.Y(n_1896)
);

BUFx3_ASAP7_75t_L g1897 ( 
.A(n_1877),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1859),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1603),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1584),
.B(n_1867),
.Y(n_1900)
);

INVx4_ASAP7_75t_L g1901 ( 
.A(n_1875),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1870),
.B(n_1866),
.Y(n_1902)
);

OAI21x1_ASAP7_75t_SL g1903 ( 
.A1(n_1656),
.A2(n_1657),
.B(n_1762),
.Y(n_1903)
);

INVx6_ASAP7_75t_L g1904 ( 
.A(n_1651),
.Y(n_1904)
);

CKINVDCx11_ASAP7_75t_R g1905 ( 
.A(n_1653),
.Y(n_1905)
);

AO31x2_ASAP7_75t_L g1906 ( 
.A1(n_1677),
.A2(n_1691),
.A3(n_1714),
.B(n_1723),
.Y(n_1906)
);

NAND2x1p5_ASAP7_75t_L g1907 ( 
.A(n_1651),
.B(n_1634),
.Y(n_1907)
);

INVx8_ASAP7_75t_L g1908 ( 
.A(n_1597),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1608),
.B(n_1868),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1875),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_L g1911 ( 
.A1(n_1728),
.A2(n_1854),
.B1(n_1869),
.B2(n_1693),
.C(n_1671),
.Y(n_1911)
);

BUFx2_ASAP7_75t_R g1912 ( 
.A(n_1701),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_1687),
.Y(n_1913)
);

BUFx12f_ASAP7_75t_L g1914 ( 
.A(n_1863),
.Y(n_1914)
);

INVx2_ASAP7_75t_SL g1915 ( 
.A(n_1863),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1603),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_SL g1917 ( 
.A1(n_1647),
.A2(n_1711),
.B(n_1674),
.Y(n_1917)
);

CKINVDCx8_ASAP7_75t_R g1918 ( 
.A(n_1701),
.Y(n_1918)
);

OAI21x1_ASAP7_75t_SL g1919 ( 
.A1(n_1718),
.A2(n_1616),
.B(n_1610),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1873),
.B(n_1663),
.Y(n_1920)
);

OR2x6_ASAP7_75t_L g1921 ( 
.A(n_1863),
.B(n_1601),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1681),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1854),
.B(n_1727),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1603),
.Y(n_1924)
);

INVx5_ASAP7_75t_L g1925 ( 
.A(n_1597),
.Y(n_1925)
);

AO31x2_ASAP7_75t_L g1926 ( 
.A1(n_1805),
.A2(n_1698),
.A3(n_1778),
.B(n_1747),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1874),
.B(n_1665),
.Y(n_1927)
);

CKINVDCx20_ASAP7_75t_R g1928 ( 
.A(n_1687),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1867),
.B(n_1745),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1748),
.B(n_1675),
.Y(n_1930)
);

CKINVDCx11_ASAP7_75t_R g1931 ( 
.A(n_1757),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1623),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1594),
.B(n_1712),
.Y(n_1933)
);

OR2x6_ASAP7_75t_L g1934 ( 
.A(n_1620),
.B(n_1842),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1756),
.B(n_1636),
.Y(n_1935)
);

NAND3xp33_ASAP7_75t_L g1936 ( 
.A(n_1829),
.B(n_1710),
.C(n_1831),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1618),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1756),
.B(n_1636),
.Y(n_1938)
);

OAI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1607),
.A2(n_1638),
.B1(n_1592),
.B2(n_1752),
.C(n_1724),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1638),
.B(n_1658),
.Y(n_1940)
);

AOI22x1_ASAP7_75t_L g1941 ( 
.A1(n_1589),
.A2(n_1646),
.B1(n_1807),
.B2(n_1755),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1871),
.B(n_1611),
.Y(n_1942)
);

OAI21x1_ASAP7_75t_SL g1943 ( 
.A1(n_1617),
.A2(n_1822),
.B(n_1595),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1643),
.B(n_1751),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1686),
.A2(n_1785),
.B(n_1731),
.Y(n_1945)
);

INVx4_ASAP7_75t_L g1946 ( 
.A(n_1651),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1619),
.Y(n_1947)
);

INVx5_ASAP7_75t_L g1948 ( 
.A(n_1597),
.Y(n_1948)
);

OAI21x1_ASAP7_75t_SL g1949 ( 
.A1(n_1593),
.A2(n_1787),
.B(n_1784),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1643),
.B(n_1844),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1661),
.Y(n_1951)
);

NOR2xp67_ASAP7_75t_L g1952 ( 
.A(n_1596),
.B(n_1828),
.Y(n_1952)
);

NAND3xp33_ASAP7_75t_L g1953 ( 
.A(n_1829),
.B(n_1710),
.C(n_1707),
.Y(n_1953)
);

AO21x2_ASAP7_75t_L g1954 ( 
.A1(n_1862),
.A2(n_1627),
.B(n_1622),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1850),
.Y(n_1955)
);

AO21x2_ASAP7_75t_L g1956 ( 
.A1(n_1862),
.A2(n_1733),
.B(n_1792),
.Y(n_1956)
);

NAND2x1p5_ASAP7_75t_L g1957 ( 
.A(n_1651),
.B(n_1634),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1661),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1686),
.A2(n_1785),
.B(n_1731),
.Y(n_1959)
);

INVx4_ASAP7_75t_L g1960 ( 
.A(n_1597),
.Y(n_1960)
);

AO21x2_ASAP7_75t_L g1961 ( 
.A1(n_1818),
.A2(n_1810),
.B(n_1682),
.Y(n_1961)
);

NAND2x1p5_ASAP7_75t_L g1962 ( 
.A(n_1729),
.B(n_1769),
.Y(n_1962)
);

INVxp33_ASAP7_75t_L g1963 ( 
.A(n_1741),
.Y(n_1963)
);

NAND2x1p5_ASAP7_75t_L g1964 ( 
.A(n_1729),
.B(n_1769),
.Y(n_1964)
);

BUFx12f_ASAP7_75t_L g1965 ( 
.A(n_1757),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1773),
.B(n_1632),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1825),
.B(n_1695),
.Y(n_1967)
);

NAND3xp33_ASAP7_75t_L g1968 ( 
.A(n_1707),
.B(n_1688),
.C(n_1713),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1661),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1844),
.B(n_1864),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1821),
.A2(n_1840),
.B(n_1835),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1785),
.A2(n_1811),
.B(n_1717),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1662),
.B(n_1760),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1800),
.Y(n_1974)
);

AO21x2_ASAP7_75t_L g1975 ( 
.A1(n_1810),
.A2(n_1719),
.B(n_1744),
.Y(n_1975)
);

BUFx12f_ASAP7_75t_L g1976 ( 
.A(n_1800),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1842),
.Y(n_1977)
);

OA21x2_ASAP7_75t_L g1978 ( 
.A1(n_1747),
.A2(n_1778),
.B(n_1725),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1844),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_L g1980 ( 
.A1(n_1666),
.A2(n_1642),
.B(n_1699),
.Y(n_1980)
);

OAI21x1_ASAP7_75t_L g1981 ( 
.A1(n_1853),
.A2(n_1802),
.B(n_1600),
.Y(n_1981)
);

INVx1_ASAP7_75t_SL g1982 ( 
.A(n_1628),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_SL g1983 ( 
.A(n_1644),
.Y(n_1983)
);

INVx3_ASAP7_75t_SL g1984 ( 
.A(n_1726),
.Y(n_1984)
);

OA21x2_ASAP7_75t_L g1985 ( 
.A1(n_1659),
.A2(n_1664),
.B(n_1633),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1864),
.B(n_1730),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1864),
.Y(n_1987)
);

INVx6_ASAP7_75t_L g1988 ( 
.A(n_1722),
.Y(n_1988)
);

AO21x2_ASAP7_75t_L g1989 ( 
.A1(n_1808),
.A2(n_1809),
.B(n_1605),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1741),
.B(n_1780),
.Y(n_1990)
);

AOI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1736),
.A2(n_1773),
.B1(n_1639),
.B2(n_1602),
.Y(n_1991)
);

BUFx2_ASAP7_75t_L g1992 ( 
.A(n_1803),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1655),
.B(n_1715),
.Y(n_1993)
);

OAI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1851),
.A2(n_1861),
.B(n_1860),
.Y(n_1994)
);

OA21x2_ASAP7_75t_L g1995 ( 
.A1(n_1588),
.A2(n_1626),
.B(n_1613),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_R g1996 ( 
.A(n_1834),
.B(n_1791),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1794),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1702),
.A2(n_1694),
.B(n_1683),
.Y(n_1998)
);

INVx8_ASAP7_75t_L g1999 ( 
.A(n_1803),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1793),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1639),
.B(n_1602),
.Y(n_2001)
);

OA21x2_ASAP7_75t_L g2002 ( 
.A1(n_1613),
.A2(n_1626),
.B(n_1735),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1797),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1648),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1598),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1648),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1797),
.Y(n_2007)
);

NAND2x1p5_ASAP7_75t_L g2008 ( 
.A(n_1649),
.B(n_1797),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1734),
.B(n_1720),
.Y(n_2009)
);

OA21x2_ASAP7_75t_L g2010 ( 
.A1(n_1735),
.A2(n_1742),
.B(n_1737),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1855),
.Y(n_2011)
);

OAI21x1_ASAP7_75t_L g2012 ( 
.A1(n_1621),
.A2(n_1629),
.B(n_1625),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1649),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1791),
.Y(n_2014)
);

AOI22x1_ASAP7_75t_L g2015 ( 
.A1(n_1766),
.A2(n_1774),
.B1(n_1771),
.B2(n_1668),
.Y(n_2015)
);

INVx8_ASAP7_75t_L g2016 ( 
.A(n_1779),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1763),
.A2(n_1703),
.B(n_1690),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1689),
.Y(n_2018)
);

NOR2x1p5_ASAP7_75t_L g2019 ( 
.A(n_1644),
.B(n_1740),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1732),
.Y(n_2020)
);

OAI21x1_ASAP7_75t_L g2021 ( 
.A1(n_1768),
.A2(n_1716),
.B(n_1705),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1743),
.Y(n_2022)
);

AO21x1_ASAP7_75t_L g2023 ( 
.A1(n_1644),
.A2(n_1843),
.B(n_1670),
.Y(n_2023)
);

OA21x2_ASAP7_75t_L g2024 ( 
.A1(n_1765),
.A2(n_1845),
.B(n_1826),
.Y(n_2024)
);

BUFx2_ASAP7_75t_L g2025 ( 
.A(n_1598),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1758),
.Y(n_2026)
);

INVxp67_ASAP7_75t_SL g2027 ( 
.A(n_1815),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1720),
.B(n_1739),
.Y(n_2028)
);

OAI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1749),
.A2(n_1750),
.B(n_1630),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1754),
.Y(n_2030)
);

AND2x2_ASAP7_75t_SL g2031 ( 
.A(n_1624),
.B(n_1754),
.Y(n_2031)
);

NOR3xp33_ASAP7_75t_L g2032 ( 
.A(n_1814),
.B(n_1709),
.C(n_1824),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1585),
.Y(n_2033)
);

INVx8_ASAP7_75t_L g2034 ( 
.A(n_1779),
.Y(n_2034)
);

CKINVDCx16_ASAP7_75t_R g2035 ( 
.A(n_1609),
.Y(n_2035)
);

INVx4_ASAP7_75t_L g2036 ( 
.A(n_1761),
.Y(n_2036)
);

BUFx2_ASAP7_75t_SL g2037 ( 
.A(n_1876),
.Y(n_2037)
);

BUFx12f_ASAP7_75t_L g2038 ( 
.A(n_1676),
.Y(n_2038)
);

AOI21x1_ASAP7_75t_L g2039 ( 
.A1(n_1635),
.A2(n_1654),
.B(n_1637),
.Y(n_2039)
);

BUFx3_ASAP7_75t_L g2040 ( 
.A(n_1761),
.Y(n_2040)
);

INVxp67_ASAP7_75t_L g2041 ( 
.A(n_1591),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1815),
.Y(n_2042)
);

CKINVDCx14_ASAP7_75t_R g2043 ( 
.A(n_1722),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1761),
.Y(n_2044)
);

AO21x2_ASAP7_75t_L g2045 ( 
.A1(n_1775),
.A2(n_1781),
.B(n_1858),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1704),
.B(n_1614),
.Y(n_2046)
);

OA21x2_ASAP7_75t_L g2047 ( 
.A1(n_1826),
.A2(n_1839),
.B(n_1848),
.Y(n_2047)
);

OAI221xp5_ASAP7_75t_SL g2048 ( 
.A1(n_1833),
.A2(n_1783),
.B1(n_1700),
.B2(n_1856),
.C(n_1848),
.Y(n_2048)
);

OAI21x1_ASAP7_75t_L g2049 ( 
.A1(n_1685),
.A2(n_1847),
.B(n_1841),
.Y(n_2049)
);

OA21x2_ASAP7_75t_L g2050 ( 
.A1(n_1837),
.A2(n_1845),
.B(n_1839),
.Y(n_2050)
);

OA21x2_ASAP7_75t_L g2051 ( 
.A1(n_1837),
.A2(n_1858),
.B(n_1856),
.Y(n_2051)
);

INVxp67_ASAP7_75t_SL g2052 ( 
.A(n_1815),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1823),
.A2(n_1836),
.B(n_1764),
.Y(n_2053)
);

AND2x6_ASAP7_75t_L g2054 ( 
.A(n_1801),
.B(n_1772),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1736),
.A2(n_1833),
.B1(n_1817),
.B2(n_1852),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1779),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1779),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_1789),
.Y(n_2058)
);

AND2x6_ASAP7_75t_L g2059 ( 
.A(n_1801),
.B(n_1772),
.Y(n_2059)
);

OAI21x1_ASAP7_75t_L g2060 ( 
.A1(n_1795),
.A2(n_1813),
.B(n_1799),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1788),
.B(n_1804),
.Y(n_2061)
);

OAI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1790),
.A2(n_1819),
.B(n_1708),
.Y(n_2062)
);

NAND2x1p5_ASAP7_75t_L g2063 ( 
.A(n_1754),
.B(n_1772),
.Y(n_2063)
);

O2A1O1Ixp33_ASAP7_75t_L g2064 ( 
.A1(n_1783),
.A2(n_1786),
.B(n_1697),
.C(n_1679),
.Y(n_2064)
);

INVx6_ASAP7_75t_L g2065 ( 
.A(n_1812),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_SL g2066 ( 
.A1(n_1631),
.A2(n_1673),
.B(n_1678),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_1672),
.A2(n_1660),
.B1(n_1806),
.B2(n_1738),
.Y(n_2067)
);

OA21x2_ASAP7_75t_L g2068 ( 
.A1(n_1786),
.A2(n_1776),
.B(n_1796),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1669),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1669),
.Y(n_2070)
);

AO21x2_ASAP7_75t_L g2071 ( 
.A1(n_1684),
.A2(n_1816),
.B(n_1782),
.Y(n_2071)
);

BUFx2_ASAP7_75t_L g2072 ( 
.A(n_1789),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_1798),
.B(n_1812),
.Y(n_2073)
);

OAI21x1_ASAP7_75t_L g2074 ( 
.A1(n_1696),
.A2(n_1759),
.B(n_1767),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1667),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1770),
.A2(n_1779),
.B(n_1849),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1652),
.B(n_1806),
.Y(n_2077)
);

A2O1A1Ixp33_ASAP7_75t_L g2078 ( 
.A1(n_1806),
.A2(n_1615),
.B(n_1746),
.C(n_1753),
.Y(n_2078)
);

OA21x2_ASAP7_75t_L g2079 ( 
.A1(n_1667),
.A2(n_1820),
.B(n_1846),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1669),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1801),
.Y(n_2081)
);

BUFx2_ASAP7_75t_SL g2082 ( 
.A(n_1615),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1721),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1669),
.Y(n_2084)
);

BUFx12f_ASAP7_75t_L g2085 ( 
.A(n_1721),
.Y(n_2085)
);

NAND2xp33_ASAP7_75t_R g2086 ( 
.A(n_1721),
.B(n_1746),
.Y(n_2086)
);

OAI21x1_ASAP7_75t_SL g2087 ( 
.A1(n_1721),
.A2(n_1746),
.B(n_1753),
.Y(n_2087)
);

O2A1O1Ixp33_ASAP7_75t_L g2088 ( 
.A1(n_1680),
.A2(n_1783),
.B(n_1872),
.C(n_1865),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1753),
.A2(n_1162),
.B1(n_1082),
.B2(n_1869),
.Y(n_2089)
);

OA21x2_ASAP7_75t_L g2090 ( 
.A1(n_1846),
.A2(n_1680),
.B(n_1753),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_1680),
.Y(n_2091)
);

NAND3xp33_ASAP7_75t_L g2092 ( 
.A(n_1865),
.B(n_1396),
.C(n_1692),
.Y(n_2092)
);

INVx4_ASAP7_75t_L g2093 ( 
.A(n_1606),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_1606),
.Y(n_2094)
);

INVx4_ASAP7_75t_L g2095 ( 
.A(n_1606),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_1877),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_1584),
.B(n_1867),
.Y(n_2097)
);

NAND2x1p5_ASAP7_75t_L g2098 ( 
.A(n_1651),
.B(n_1202),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1650),
.Y(n_2099)
);

INVxp67_ASAP7_75t_SL g2100 ( 
.A(n_1872),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1606),
.Y(n_2101)
);

AND2x4_ASAP7_75t_L g2102 ( 
.A(n_1870),
.B(n_1675),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1870),
.B(n_1584),
.Y(n_2103)
);

CKINVDCx16_ASAP7_75t_R g2104 ( 
.A(n_1606),
.Y(n_2104)
);

AOI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_1869),
.A2(n_1162),
.B1(n_1082),
.B2(n_1584),
.Y(n_2105)
);

INVxp33_ASAP7_75t_L g2106 ( 
.A(n_1832),
.Y(n_2106)
);

CKINVDCx6p67_ASAP7_75t_R g2107 ( 
.A(n_1606),
.Y(n_2107)
);

OA21x2_ASAP7_75t_L g2108 ( 
.A1(n_1640),
.A2(n_1645),
.B(n_1641),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1584),
.B(n_1870),
.Y(n_2109)
);

INVx4_ASAP7_75t_L g2110 ( 
.A(n_1606),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1584),
.B(n_1867),
.Y(n_2111)
);

INVx5_ASAP7_75t_L g2112 ( 
.A(n_1597),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1586),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1586),
.Y(n_2114)
);

OAI21x1_ASAP7_75t_SL g2115 ( 
.A1(n_1872),
.A2(n_1587),
.B(n_1777),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1586),
.Y(n_2116)
);

AO21x1_ASAP7_75t_SL g2117 ( 
.A1(n_1587),
.A2(n_1760),
.B(n_1593),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1584),
.B(n_1870),
.Y(n_2118)
);

AO21x2_ASAP7_75t_L g2119 ( 
.A1(n_1590),
.A2(n_1830),
.B(n_1827),
.Y(n_2119)
);

AO21x2_ASAP7_75t_L g2120 ( 
.A1(n_1590),
.A2(n_1830),
.B(n_1827),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_1885),
.B(n_2103),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1973),
.B(n_2100),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1878),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_1900),
.A2(n_2111),
.B1(n_2097),
.B2(n_2032),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1880),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_L g2126 ( 
.A1(n_2031),
.A2(n_2100),
.B1(n_2063),
.B2(n_2089),
.Y(n_2126)
);

CKINVDCx6p67_ASAP7_75t_R g2127 ( 
.A(n_1879),
.Y(n_2127)
);

INVx2_ASAP7_75t_SL g2128 ( 
.A(n_1879),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_1942),
.B(n_1909),
.Y(n_2129)
);

CKINVDCx6p67_ASAP7_75t_R g2130 ( 
.A(n_1879),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1927),
.B(n_2046),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1886),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1893),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1896),
.Y(n_2134)
);

BUFx2_ASAP7_75t_L g2135 ( 
.A(n_1934),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_1900),
.A2(n_2097),
.B1(n_2111),
.B2(n_2032),
.Y(n_2136)
);

OAI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_2031),
.A2(n_2063),
.B1(n_2083),
.B2(n_1939),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1983),
.A2(n_2019),
.B1(n_1911),
.B2(n_2082),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_SL g2139 ( 
.A1(n_1983),
.A2(n_2052),
.B1(n_2027),
.B2(n_1939),
.Y(n_2139)
);

INVx2_ASAP7_75t_SL g2140 ( 
.A(n_1999),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_1929),
.B(n_1923),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1898),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2113),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_1935),
.Y(n_2144)
);

OAI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2083),
.A2(n_1960),
.B1(n_2105),
.B2(n_1925),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_1911),
.A2(n_2001),
.B1(n_2023),
.B2(n_1933),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2001),
.A2(n_1991),
.B1(n_2055),
.B2(n_1933),
.Y(n_2147)
);

AO21x1_ASAP7_75t_L g2148 ( 
.A1(n_2088),
.A2(n_1960),
.B(n_2086),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2114),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_1935),
.Y(n_2150)
);

INVx2_ASAP7_75t_SL g2151 ( 
.A(n_1999),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2116),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1932),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1997),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_2077),
.A2(n_2118),
.B1(n_2109),
.B2(n_2052),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1993),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1993),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1946),
.Y(n_2158)
);

CKINVDCx20_ASAP7_75t_R g2159 ( 
.A(n_1892),
.Y(n_2159)
);

INVx4_ASAP7_75t_L g2160 ( 
.A(n_1914),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1925),
.B(n_1948),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_1938),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2022),
.B(n_1920),
.Y(n_2163)
);

AO21x2_ASAP7_75t_L g2164 ( 
.A1(n_1945),
.A2(n_1959),
.B(n_2087),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_L g2165 ( 
.A1(n_2027),
.A2(n_2092),
.B1(n_1940),
.B2(n_1894),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1990),
.B(n_1963),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_1938),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2020),
.Y(n_2168)
);

OAI21x1_ASAP7_75t_SL g2169 ( 
.A1(n_1891),
.A2(n_2115),
.B(n_1943),
.Y(n_2169)
);

CKINVDCx20_ASAP7_75t_R g2170 ( 
.A(n_1892),
.Y(n_2170)
);

INVx4_ASAP7_75t_L g2171 ( 
.A(n_1914),
.Y(n_2171)
);

BUFx2_ASAP7_75t_SL g2172 ( 
.A(n_2093),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2020),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_1990),
.B(n_1963),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_1934),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_1934),
.Y(n_2176)
);

OAI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_1925),
.A2(n_1948),
.B1(n_2112),
.B2(n_1908),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1930),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1902),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_2107),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_2008),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2017),
.B(n_1979),
.Y(n_2182)
);

INVx3_ASAP7_75t_L g2183 ( 
.A(n_1946),
.Y(n_2183)
);

HB1xp67_ASAP7_75t_L g2184 ( 
.A(n_2008),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_L g2185 ( 
.A1(n_1881),
.A2(n_2085),
.B1(n_1986),
.B2(n_1949),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2000),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2000),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2099),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2099),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2106),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_1996),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_1996),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2106),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2030),
.Y(n_2194)
);

BUFx3_ASAP7_75t_L g2195 ( 
.A(n_1907),
.Y(n_2195)
);

INVx1_ASAP7_75t_SL g2196 ( 
.A(n_2081),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1977),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1944),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_1970),
.Y(n_2199)
);

INVx2_ASAP7_75t_SL g2200 ( 
.A(n_1999),
.Y(n_2200)
);

INVx3_ASAP7_75t_SL g2201 ( 
.A(n_2101),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2061),
.B(n_1967),
.Y(n_2202)
);

BUFx12f_ASAP7_75t_L g2203 ( 
.A(n_1905),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1951),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1958),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_2011),
.B(n_1966),
.Y(n_2206)
);

OR2x6_ASAP7_75t_L g2207 ( 
.A(n_1908),
.B(n_2016),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1969),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1899),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2018),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1916),
.Y(n_2211)
);

BUFx2_ASAP7_75t_L g2212 ( 
.A(n_1897),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1905),
.Y(n_2213)
);

OR2x2_ASAP7_75t_L g2214 ( 
.A(n_1955),
.B(n_1887),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_1925),
.Y(n_2215)
);

OR2x6_ASAP7_75t_L g2216 ( 
.A(n_1908),
.B(n_2016),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1924),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1966),
.Y(n_2218)
);

AO21x2_ASAP7_75t_L g2219 ( 
.A1(n_1917),
.A2(n_1919),
.B(n_2078),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1890),
.Y(n_2220)
);

BUFx2_ASAP7_75t_L g2221 ( 
.A(n_1897),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1890),
.Y(n_2222)
);

BUFx2_ASAP7_75t_L g2223 ( 
.A(n_2096),
.Y(n_2223)
);

BUFx2_ASAP7_75t_L g2224 ( 
.A(n_2096),
.Y(n_2224)
);

OAI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_1953),
.A2(n_1936),
.B(n_1968),
.Y(n_2225)
);

AOI22xp33_ASAP7_75t_L g2226 ( 
.A1(n_2085),
.A2(n_1937),
.B1(n_1947),
.B2(n_2071),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1922),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1922),
.Y(n_2228)
);

BUFx2_ASAP7_75t_R g2229 ( 
.A(n_2101),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_2104),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_2098),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2025),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_1931),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2005),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_2098),
.Y(n_2235)
);

AO21x1_ASAP7_75t_SL g2236 ( 
.A1(n_1948),
.A2(n_2112),
.B(n_1987),
.Y(n_2236)
);

NOR2x1_ASAP7_75t_R g2237 ( 
.A(n_1931),
.B(n_2093),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_1948),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2003),
.Y(n_2239)
);

OR2x6_ASAP7_75t_L g2240 ( 
.A(n_2016),
.B(n_2034),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2007),
.Y(n_2241)
);

BUFx3_ASAP7_75t_L g2242 ( 
.A(n_1907),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2033),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_1957),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_1957),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2112),
.A2(n_2048),
.B1(n_2078),
.B2(n_2067),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2004),
.Y(n_2247)
);

AOI22xp33_ASAP7_75t_L g2248 ( 
.A1(n_2071),
.A2(n_2051),
.B1(n_2050),
.B2(n_2047),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2006),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_1895),
.B(n_2102),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_SL g2251 ( 
.A(n_2042),
.Y(n_2251)
);

AOI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_2102),
.A2(n_2035),
.B1(n_2073),
.B2(n_2041),
.Y(n_2252)
);

BUFx2_ASAP7_75t_L g2253 ( 
.A(n_2043),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2006),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2013),
.Y(n_2255)
);

BUFx2_ASAP7_75t_SL g2256 ( 
.A(n_2095),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1952),
.Y(n_2257)
);

HB1xp67_ASAP7_75t_L g2258 ( 
.A(n_1950),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_1904),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2013),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_1904),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2069),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2070),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2080),
.Y(n_2264)
);

AOI222xp33_ASAP7_75t_L g2265 ( 
.A1(n_2041),
.A2(n_1965),
.B1(n_2042),
.B2(n_1888),
.C1(n_1884),
.C2(n_2110),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2084),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_1950),
.Y(n_2267)
);

INVx3_ASAP7_75t_L g2268 ( 
.A(n_1904),
.Y(n_2268)
);

NAND2x1p5_ASAP7_75t_L g2269 ( 
.A(n_2072),
.B(n_1901),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2090),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2043),
.Y(n_2271)
);

OR2x6_ASAP7_75t_L g2272 ( 
.A(n_2034),
.B(n_1889),
.Y(n_2272)
);

INVx2_ASAP7_75t_SL g2273 ( 
.A(n_2095),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2017),
.B(n_1972),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2090),
.Y(n_2275)
);

AOI22xp33_ASAP7_75t_L g2276 ( 
.A1(n_2047),
.A2(n_2050),
.B1(n_2051),
.B2(n_2067),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2090),
.Y(n_2277)
);

INVx3_ASAP7_75t_L g2278 ( 
.A(n_2034),
.Y(n_2278)
);

AOI22xp33_ASAP7_75t_SL g2279 ( 
.A1(n_1903),
.A2(n_2059),
.B1(n_2054),
.B2(n_2024),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2037),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1962),
.Y(n_2281)
);

BUFx12f_ASAP7_75t_L g2282 ( 
.A(n_2110),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_1976),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1962),
.Y(n_2284)
);

BUFx3_ASAP7_75t_L g2285 ( 
.A(n_1964),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1964),
.Y(n_2286)
);

BUFx2_ASAP7_75t_L g2287 ( 
.A(n_1921),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2048),
.A2(n_1978),
.B1(n_2010),
.B2(n_2002),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1972),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2079),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_1982),
.B(n_2073),
.Y(n_2291)
);

BUFx4f_ASAP7_75t_SL g2292 ( 
.A(n_1976),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2058),
.B(n_2065),
.Y(n_2293)
);

INVx2_ASAP7_75t_SL g2294 ( 
.A(n_1883),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2079),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2044),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2065),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2065),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_1988),
.B(n_2014),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2075),
.Y(n_2300)
);

OR2x2_ASAP7_75t_L g2301 ( 
.A(n_1921),
.B(n_1992),
.Y(n_2301)
);

BUFx4f_ASAP7_75t_L g2302 ( 
.A(n_1965),
.Y(n_2302)
);

HB1xp67_ASAP7_75t_L g2303 ( 
.A(n_2044),
.Y(n_2303)
);

OR2x6_ASAP7_75t_L g2304 ( 
.A(n_2056),
.B(n_1988),
.Y(n_2304)
);

CKINVDCx8_ASAP7_75t_R g2305 ( 
.A(n_1974),
.Y(n_2305)
);

BUFx2_ASAP7_75t_L g2306 ( 
.A(n_2038),
.Y(n_2306)
);

BUFx12f_ASAP7_75t_L g2307 ( 
.A(n_1901),
.Y(n_2307)
);

OAI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_1978),
.A2(n_2010),
.B1(n_2002),
.B2(n_2088),
.Y(n_2308)
);

OR2x6_ASAP7_75t_L g2309 ( 
.A(n_2056),
.B(n_1988),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2014),
.B(n_1984),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2122),
.B(n_2146),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_2231),
.Y(n_2312)
);

INVxp33_ASAP7_75t_SL g2313 ( 
.A(n_2237),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2122),
.B(n_2091),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2123),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2125),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2132),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2146),
.B(n_2163),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_2124),
.A2(n_2068),
.B1(n_2024),
.B2(n_1941),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2129),
.B(n_2131),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2163),
.B(n_2045),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2133),
.Y(n_2322)
);

BUFx3_ASAP7_75t_L g2323 ( 
.A(n_2195),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2134),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2142),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2143),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2121),
.B(n_2028),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2202),
.B(n_2028),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2149),
.Y(n_2329)
);

OAI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_2137),
.A2(n_2002),
.B1(n_1978),
.B2(n_2010),
.Y(n_2330)
);

INVx4_ASAP7_75t_L g2331 ( 
.A(n_2127),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2218),
.B(n_2081),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2152),
.Y(n_2333)
);

OAI211xp5_ASAP7_75t_SL g2334 ( 
.A1(n_2124),
.A2(n_2136),
.B(n_2265),
.C(n_2252),
.Y(n_2334)
);

AOI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2136),
.A2(n_2117),
.B1(n_2029),
.B2(n_1971),
.Y(n_2335)
);

AOI222xp33_ASAP7_75t_L g2336 ( 
.A1(n_2141),
.A2(n_2059),
.B1(n_1984),
.B2(n_2094),
.C1(n_1915),
.C2(n_1994),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2153),
.Y(n_2337)
);

INVx1_ASAP7_75t_SL g2338 ( 
.A(n_2196),
.Y(n_2338)
);

AOI22xp33_ASAP7_75t_L g2339 ( 
.A1(n_2137),
.A2(n_2066),
.B1(n_2059),
.B2(n_1961),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2154),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2141),
.B(n_2038),
.Y(n_2341)
);

OAI21xp5_ASAP7_75t_SL g2342 ( 
.A1(n_2139),
.A2(n_2064),
.B(n_1998),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2291),
.B(n_2009),
.Y(n_2343)
);

HB1xp67_ASAP7_75t_L g2344 ( 
.A(n_2144),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2243),
.Y(n_2345)
);

BUFx2_ASAP7_75t_L g2346 ( 
.A(n_2285),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2168),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2139),
.A2(n_1961),
.B1(n_2015),
.B2(n_1995),
.Y(n_2348)
);

INVx5_ASAP7_75t_L g2349 ( 
.A(n_2207),
.Y(n_2349)
);

BUFx6f_ASAP7_75t_L g2350 ( 
.A(n_2236),
.Y(n_2350)
);

INVx2_ASAP7_75t_SL g2351 ( 
.A(n_2292),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2173),
.Y(n_2352)
);

BUFx2_ASAP7_75t_L g2353 ( 
.A(n_2285),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2206),
.B(n_2196),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2178),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_2195),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2156),
.Y(n_2357)
);

OR2x2_ASAP7_75t_L g2358 ( 
.A(n_2214),
.B(n_1910),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2166),
.B(n_2036),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2157),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2190),
.Y(n_2361)
);

INVx5_ASAP7_75t_L g2362 ( 
.A(n_2207),
.Y(n_2362)
);

INVxp67_ASAP7_75t_SL g2363 ( 
.A(n_2144),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_2231),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_2242),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2193),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2174),
.B(n_2036),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2299),
.B(n_2076),
.Y(n_2368)
);

INVx3_ASAP7_75t_L g2369 ( 
.A(n_2235),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2212),
.B(n_1989),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2221),
.B(n_1989),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2223),
.B(n_2062),
.Y(n_2372)
);

OR2x2_ASAP7_75t_L g2373 ( 
.A(n_2179),
.B(n_1910),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2224),
.B(n_2062),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2199),
.B(n_2049),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2165),
.B(n_1926),
.Y(n_2376)
);

BUFx2_ASAP7_75t_L g2377 ( 
.A(n_2272),
.Y(n_2377)
);

OAI21xp5_ASAP7_75t_SL g2378 ( 
.A1(n_2138),
.A2(n_2057),
.B(n_1912),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2276),
.B(n_1926),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2199),
.B(n_2049),
.Y(n_2380)
);

OR2x2_ASAP7_75t_L g2381 ( 
.A(n_2301),
.B(n_2150),
.Y(n_2381)
);

OAI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2138),
.A2(n_1995),
.B1(n_2039),
.B2(n_2108),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2150),
.B(n_1926),
.Y(n_2383)
);

INVx3_ASAP7_75t_L g2384 ( 
.A(n_2242),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2272),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2287),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2197),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2232),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2250),
.B(n_2074),
.Y(n_2389)
);

BUFx2_ASAP7_75t_L g2390 ( 
.A(n_2272),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2209),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2293),
.B(n_2147),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2155),
.B(n_1906),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2211),
.Y(n_2394)
);

INVx2_ASAP7_75t_SL g2395 ( 
.A(n_2292),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_2155),
.B(n_1974),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2253),
.B(n_1906),
.Y(n_2397)
);

OR2x2_ASAP7_75t_L g2398 ( 
.A(n_2162),
.B(n_1926),
.Y(n_2398)
);

INVx2_ASAP7_75t_SL g2399 ( 
.A(n_2180),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2271),
.B(n_1906),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2160),
.B(n_1975),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2217),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2204),
.Y(n_2403)
);

INVx4_ASAP7_75t_R g2404 ( 
.A(n_2251),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2297),
.B(n_1906),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2298),
.B(n_2040),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_2162),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2167),
.B(n_2040),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2205),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2208),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2186),
.Y(n_2411)
);

HB1xp67_ASAP7_75t_L g2412 ( 
.A(n_2296),
.Y(n_2412)
);

HB1xp67_ASAP7_75t_L g2413 ( 
.A(n_2296),
.Y(n_2413)
);

INVxp67_ASAP7_75t_L g2414 ( 
.A(n_2182),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2303),
.Y(n_2415)
);

HB1xp67_ASAP7_75t_L g2416 ( 
.A(n_2303),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2187),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_L g2418 ( 
.A1(n_2246),
.A2(n_2130),
.B1(n_2126),
.B2(n_2191),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2245),
.B(n_2026),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2269),
.B(n_2135),
.Y(n_2420)
);

BUFx3_ASAP7_75t_L g2421 ( 
.A(n_2140),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2188),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2189),
.Y(n_2423)
);

AOI222xp33_ASAP7_75t_L g2424 ( 
.A1(n_2302),
.A2(n_1928),
.B1(n_1913),
.B2(n_1980),
.C1(n_2060),
.C2(n_2012),
.Y(n_2424)
);

HB1xp67_ASAP7_75t_L g2425 ( 
.A(n_2300),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2269),
.B(n_2060),
.Y(n_2426)
);

OAI21xp5_ASAP7_75t_SL g2427 ( 
.A1(n_2265),
.A2(n_1912),
.B(n_1918),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2175),
.B(n_1975),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2244),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2262),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2290),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2185),
.B(n_2194),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2185),
.B(n_1954),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2176),
.B(n_2021),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2263),
.Y(n_2435)
);

AOI22xp33_ASAP7_75t_L g2436 ( 
.A1(n_2246),
.A2(n_1882),
.B1(n_2119),
.B2(n_2120),
.Y(n_2436)
);

BUFx2_ASAP7_75t_L g2437 ( 
.A(n_2158),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_2180),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2234),
.B(n_2053),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2160),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_2126),
.A2(n_1882),
.B1(n_2119),
.B2(n_2120),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2264),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2266),
.Y(n_2443)
);

HB1xp67_ASAP7_75t_L g2444 ( 
.A(n_2182),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2239),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2183),
.B(n_2053),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2183),
.B(n_1985),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2258),
.B(n_2267),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2241),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2257),
.Y(n_2450)
);

INVx4_ASAP7_75t_L g2451 ( 
.A(n_2171),
.Y(n_2451)
);

INVx3_ASAP7_75t_L g2452 ( 
.A(n_2244),
.Y(n_2452)
);

OR2x6_ASAP7_75t_L g2453 ( 
.A(n_2207),
.B(n_1981),
.Y(n_2453)
);

HB1xp67_ASAP7_75t_L g2454 ( 
.A(n_2274),
.Y(n_2454)
);

INVx2_ASAP7_75t_SL g2455 ( 
.A(n_2171),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2281),
.B(n_2284),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2220),
.Y(n_2457)
);

CKINVDCx5p33_ASAP7_75t_R g2458 ( 
.A(n_2159),
.Y(n_2458)
);

NOR2x1_ASAP7_75t_L g2459 ( 
.A(n_2172),
.B(n_1928),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_2334),
.B(n_2128),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2318),
.B(n_2288),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2345),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2320),
.B(n_2267),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2316),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2318),
.B(n_2288),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2317),
.Y(n_2466)
);

INVxp67_ASAP7_75t_L g2467 ( 
.A(n_2412),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2334),
.B(n_2192),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2343),
.B(n_2354),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2322),
.Y(n_2470)
);

OAI21xp33_ASAP7_75t_L g2471 ( 
.A1(n_2342),
.A2(n_2226),
.B(n_2248),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_2336),
.B(n_2279),
.Y(n_2472)
);

AOI222xp33_ASAP7_75t_L g2473 ( 
.A1(n_2427),
.A2(n_2302),
.B1(n_2203),
.B2(n_2226),
.C1(n_2225),
.C2(n_2248),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2311),
.B(n_2308),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2324),
.Y(n_2475)
);

INVxp67_ASAP7_75t_SL g2476 ( 
.A(n_2425),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2325),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2326),
.Y(n_2478)
);

INVxp67_ASAP7_75t_SL g2479 ( 
.A(n_2444),
.Y(n_2479)
);

BUFx3_ASAP7_75t_L g2480 ( 
.A(n_2350),
.Y(n_2480)
);

INVxp67_ASAP7_75t_L g2481 ( 
.A(n_2412),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2329),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2333),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2337),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2340),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2355),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2328),
.B(n_2327),
.Y(n_2487)
);

INVx4_ASAP7_75t_L g2488 ( 
.A(n_2350),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2311),
.B(n_2270),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2392),
.B(n_2198),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2387),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2388),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2357),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2360),
.Y(n_2494)
);

INVxp67_ASAP7_75t_L g2495 ( 
.A(n_2413),
.Y(n_2495)
);

AOI22xp33_ASAP7_75t_L g2496 ( 
.A1(n_2313),
.A2(n_2148),
.B1(n_2145),
.B2(n_2219),
.Y(n_2496)
);

AND2x2_ASAP7_75t_L g2497 ( 
.A(n_2338),
.B(n_2247),
.Y(n_2497)
);

INVxp67_ASAP7_75t_L g2498 ( 
.A(n_2413),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2321),
.B(n_2275),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2338),
.B(n_2249),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2391),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2394),
.Y(n_2502)
);

OR2x2_ASAP7_75t_L g2503 ( 
.A(n_2381),
.B(n_2164),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2402),
.Y(n_2504)
);

INVxp67_ASAP7_75t_L g2505 ( 
.A(n_2415),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2359),
.B(n_2254),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2403),
.Y(n_2507)
);

BUFx2_ASAP7_75t_L g2508 ( 
.A(n_2350),
.Y(n_2508)
);

AOI22xp33_ASAP7_75t_L g2509 ( 
.A1(n_2313),
.A2(n_2145),
.B1(n_2219),
.B2(n_2280),
.Y(n_2509)
);

HB1xp67_ASAP7_75t_L g2510 ( 
.A(n_2415),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2367),
.B(n_2255),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2321),
.B(n_2277),
.Y(n_2512)
);

NOR2xp67_ASAP7_75t_L g2513 ( 
.A(n_2451),
.B(n_2282),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2397),
.B(n_2260),
.Y(n_2514)
);

AND2x4_ASAP7_75t_SL g2515 ( 
.A(n_2350),
.B(n_2159),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2400),
.B(n_2181),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2409),
.Y(n_2517)
);

AOI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2335),
.A2(n_1985),
.B1(n_2279),
.B2(n_1956),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_2448),
.B(n_2164),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2414),
.B(n_2225),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2410),
.Y(n_2521)
);

OR2x6_ASAP7_75t_L g2522 ( 
.A(n_2453),
.B(n_2216),
.Y(n_2522)
);

OAI22xp5_ASAP7_75t_L g2523 ( 
.A1(n_2418),
.A2(n_2216),
.B1(n_2240),
.B2(n_2184),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2414),
.B(n_2295),
.Y(n_2524)
);

NOR2xp33_ASAP7_75t_L g2525 ( 
.A(n_2396),
.B(n_2286),
.Y(n_2525)
);

AND2x2_ASAP7_75t_SL g2526 ( 
.A(n_2339),
.B(n_2161),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2456),
.B(n_2181),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2445),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2449),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2332),
.B(n_2184),
.Y(n_2530)
);

INVxp67_ASAP7_75t_SL g2531 ( 
.A(n_2444),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2315),
.Y(n_2532)
);

OAI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2418),
.A2(n_2216),
.B1(n_2240),
.B2(n_2215),
.Y(n_2533)
);

OR2x2_ASAP7_75t_L g2534 ( 
.A(n_2361),
.B(n_2366),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2430),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2315),
.Y(n_2536)
);

INVx1_ASAP7_75t_SL g2537 ( 
.A(n_2421),
.Y(n_2537)
);

BUFx2_ASAP7_75t_L g2538 ( 
.A(n_2437),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2405),
.B(n_2435),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2336),
.B(n_2424),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2335),
.A2(n_1985),
.B1(n_2169),
.B2(n_2294),
.Y(n_2541)
);

AND2x4_ASAP7_75t_L g2542 ( 
.A(n_2372),
.B(n_2161),
.Y(n_2542)
);

HB1xp67_ASAP7_75t_L g2543 ( 
.A(n_2416),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2386),
.B(n_2347),
.Y(n_2544)
);

INVx2_ASAP7_75t_SL g2545 ( 
.A(n_2404),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2450),
.B(n_2210),
.Y(n_2546)
);

INVx2_ASAP7_75t_SL g2547 ( 
.A(n_2451),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2442),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2421),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2443),
.B(n_2289),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2457),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2349),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2416),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2352),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2411),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2408),
.B(n_2222),
.Y(n_2556)
);

BUFx2_ASAP7_75t_L g2557 ( 
.A(n_2323),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2417),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2422),
.Y(n_2559)
);

OR2x2_ASAP7_75t_L g2560 ( 
.A(n_2344),
.B(n_2274),
.Y(n_2560)
);

BUFx3_ASAP7_75t_L g2561 ( 
.A(n_2323),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2344),
.B(n_2310),
.Y(n_2562)
);

AND2x2_ASAP7_75t_SL g2563 ( 
.A(n_2339),
.B(n_2215),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2423),
.Y(n_2564)
);

NAND2x1p5_ASAP7_75t_L g2565 ( 
.A(n_2349),
.B(n_2278),
.Y(n_2565)
);

INVxp67_ASAP7_75t_L g2566 ( 
.A(n_2538),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2532),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2514),
.B(n_2393),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2539),
.B(n_2383),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2516),
.B(n_2447),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2462),
.Y(n_2571)
);

OAI21xp33_ASAP7_75t_SL g2572 ( 
.A1(n_2540),
.A2(n_2424),
.B(n_2331),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2489),
.B(n_2439),
.Y(n_2573)
);

INVx2_ASAP7_75t_SL g2574 ( 
.A(n_2480),
.Y(n_2574)
);

OR2x2_ASAP7_75t_L g2575 ( 
.A(n_2539),
.B(n_2398),
.Y(n_2575)
);

INVx2_ASAP7_75t_SL g2576 ( 
.A(n_2480),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2536),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2493),
.B(n_2374),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2494),
.B(n_2432),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2464),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2537),
.B(n_2440),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2489),
.B(n_2454),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2463),
.B(n_2432),
.Y(n_2583)
);

BUFx2_ASAP7_75t_L g2584 ( 
.A(n_2476),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2524),
.Y(n_2585)
);

OAI221xp5_ASAP7_75t_SL g2586 ( 
.A1(n_2473),
.A2(n_2378),
.B1(n_2396),
.B2(n_2441),
.C(n_2348),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2486),
.B(n_2370),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2524),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2492),
.B(n_2371),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2469),
.B(n_2454),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2461),
.B(n_2375),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2554),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2461),
.B(n_2380),
.Y(n_2593)
);

NOR2xp33_ASAP7_75t_L g2594 ( 
.A(n_2549),
.B(n_2455),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2465),
.B(n_2389),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2465),
.B(n_2428),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2503),
.B(n_2314),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2490),
.B(n_2407),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_2522),
.B(n_2453),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2474),
.B(n_2441),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2466),
.B(n_2407),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2555),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2522),
.B(n_2453),
.Y(n_2603)
);

NAND2x1p5_ASAP7_75t_L g2604 ( 
.A(n_2488),
.B(n_2349),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2474),
.B(n_2542),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2470),
.B(n_2368),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2542),
.B(n_2379),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2520),
.B(n_2499),
.Y(n_2608)
);

AOI32xp33_ASAP7_75t_L g2609 ( 
.A1(n_2515),
.A2(n_2459),
.A3(n_2331),
.B1(n_2341),
.B2(n_2390),
.Y(n_2609)
);

AND2x4_ASAP7_75t_L g2610 ( 
.A(n_2522),
.B(n_2446),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2520),
.B(n_2379),
.Y(n_2611)
);

OR2x2_ASAP7_75t_L g2612 ( 
.A(n_2560),
.B(n_2314),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2475),
.B(n_2363),
.Y(n_2613)
);

AND2x4_ASAP7_75t_L g2614 ( 
.A(n_2488),
.B(n_2401),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2558),
.Y(n_2615)
);

AND2x4_ASAP7_75t_L g2616 ( 
.A(n_2519),
.B(n_2434),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2499),
.B(n_2431),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2512),
.B(n_2431),
.Y(n_2618)
);

INVx2_ASAP7_75t_SL g2619 ( 
.A(n_2508),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2497),
.B(n_2376),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2477),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2478),
.Y(n_2622)
);

OR2x2_ASAP7_75t_L g2623 ( 
.A(n_2476),
.B(n_2376),
.Y(n_2623)
);

OR2x2_ASAP7_75t_L g2624 ( 
.A(n_2590),
.B(n_2510),
.Y(n_2624)
);

OR2x2_ASAP7_75t_L g2625 ( 
.A(n_2590),
.B(n_2510),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2592),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2567),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_L g2628 ( 
.A(n_2572),
.B(n_2460),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2592),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2567),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2605),
.B(n_2487),
.Y(n_2631)
);

OAI21xp33_ASAP7_75t_L g2632 ( 
.A1(n_2586),
.A2(n_2540),
.B(n_2472),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2602),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2605),
.B(n_2500),
.Y(n_2634)
);

OR2x2_ASAP7_75t_L g2635 ( 
.A(n_2569),
.B(n_2543),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2608),
.B(n_2433),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2611),
.B(n_2482),
.Y(n_2637)
);

OR2x2_ASAP7_75t_L g2638 ( 
.A(n_2569),
.B(n_2543),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2581),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2602),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2570),
.B(n_2553),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_2575),
.B(n_2553),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2615),
.Y(n_2643)
);

NOR2xp33_ASAP7_75t_L g2644 ( 
.A(n_2566),
.B(n_2460),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2615),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2570),
.B(n_2506),
.Y(n_2646)
);

OAI21xp5_ASAP7_75t_L g2647 ( 
.A1(n_2594),
.A2(n_2513),
.B(n_2341),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2620),
.B(n_2511),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2571),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2599),
.B(n_2603),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2575),
.B(n_2479),
.Y(n_2651)
);

NAND2x1p5_ASAP7_75t_L g2652 ( 
.A(n_2599),
.B(n_2561),
.Y(n_2652)
);

INVxp67_ASAP7_75t_L g2653 ( 
.A(n_2584),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2620),
.B(n_2526),
.Y(n_2654)
);

BUFx2_ASAP7_75t_L g2655 ( 
.A(n_2604),
.Y(n_2655)
);

OR2x2_ASAP7_75t_L g2656 ( 
.A(n_2597),
.B(n_2479),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2580),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2599),
.B(n_2531),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2611),
.B(n_2483),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2577),
.Y(n_2660)
);

INVx3_ASAP7_75t_L g2661 ( 
.A(n_2614),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2621),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2607),
.B(n_2526),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2600),
.B(n_2484),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2622),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2585),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2585),
.Y(n_2667)
);

AOI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2600),
.A2(n_2468),
.B1(n_2533),
.B2(n_2472),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2607),
.B(n_2556),
.Y(n_2669)
);

AND2x4_ASAP7_75t_L g2670 ( 
.A(n_2603),
.B(n_2531),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2588),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2577),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2608),
.B(n_2485),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2588),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2617),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2635),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2636),
.B(n_2596),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2638),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2642),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2627),
.Y(n_2680)
);

OAI22xp33_ASAP7_75t_SL g2681 ( 
.A1(n_2628),
.A2(n_2655),
.B1(n_2652),
.B2(n_2668),
.Y(n_2681)
);

OAI21xp33_ASAP7_75t_L g2682 ( 
.A1(n_2632),
.A2(n_2496),
.B(n_2468),
.Y(n_2682)
);

AOI211xp5_ASAP7_75t_L g2683 ( 
.A1(n_2628),
.A2(n_2533),
.B(n_2523),
.C(n_2603),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2666),
.Y(n_2684)
);

HB1xp67_ASAP7_75t_L g2685 ( 
.A(n_2653),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2667),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2636),
.B(n_2596),
.Y(n_2687)
);

AND4x1_ASAP7_75t_L g2688 ( 
.A(n_2647),
.B(n_2496),
.C(n_2509),
.D(n_2229),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2671),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2674),
.Y(n_2690)
);

INVx1_ASAP7_75t_SL g2691 ( 
.A(n_2639),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2624),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2641),
.B(n_2616),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2644),
.B(n_2233),
.Y(n_2694)
);

OAI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_2652),
.A2(n_2523),
.B1(n_2557),
.B2(n_2561),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2664),
.B(n_2591),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2627),
.Y(n_2697)
);

INVxp67_ASAP7_75t_SL g2698 ( 
.A(n_2653),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2630),
.Y(n_2699)
);

OR2x2_ASAP7_75t_L g2700 ( 
.A(n_2625),
.B(n_2623),
.Y(n_2700)
);

OAI22xp5_ASAP7_75t_L g2701 ( 
.A1(n_2658),
.A2(n_2509),
.B1(n_2609),
.B2(n_2670),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2626),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2629),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2630),
.Y(n_2704)
);

INVxp33_ASAP7_75t_L g2705 ( 
.A(n_2644),
.Y(n_2705)
);

AND2x2_ASAP7_75t_SL g2706 ( 
.A(n_2650),
.B(n_2563),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2658),
.Y(n_2707)
);

INVxp67_ASAP7_75t_L g2708 ( 
.A(n_2656),
.Y(n_2708)
);

NAND4xp75_ASAP7_75t_L g2709 ( 
.A(n_2663),
.B(n_2545),
.C(n_2563),
.D(n_2547),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2633),
.Y(n_2710)
);

NAND3xp33_ASAP7_75t_L g2711 ( 
.A(n_2651),
.B(n_2541),
.C(n_2471),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2664),
.B(n_2675),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2640),
.Y(n_2713)
);

OR2x2_ASAP7_75t_L g2714 ( 
.A(n_2637),
.B(n_2623),
.Y(n_2714)
);

OAI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2658),
.A2(n_2604),
.B1(n_2541),
.B2(n_2385),
.Y(n_2715)
);

HB1xp67_ASAP7_75t_L g2716 ( 
.A(n_2660),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2637),
.B(n_2591),
.Y(n_2717)
);

AND2x4_ASAP7_75t_SL g2718 ( 
.A(n_2646),
.B(n_2170),
.Y(n_2718)
);

AOI21xp33_ASAP7_75t_L g2719 ( 
.A1(n_2649),
.A2(n_2358),
.B(n_2562),
.Y(n_2719)
);

OAI22xp33_ASAP7_75t_SL g2720 ( 
.A1(n_2650),
.A2(n_2604),
.B1(n_2670),
.B2(n_2661),
.Y(n_2720)
);

NOR2xp33_ASAP7_75t_SL g2721 ( 
.A(n_2670),
.B(n_2229),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2660),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2707),
.B(n_2650),
.Y(n_2723)
);

NOR3xp33_ASAP7_75t_L g2724 ( 
.A(n_2681),
.B(n_2682),
.C(n_2701),
.Y(n_2724)
);

AOI22xp33_ASAP7_75t_L g2725 ( 
.A1(n_2706),
.A2(n_2654),
.B1(n_2610),
.B2(n_2616),
.Y(n_2725)
);

AOI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2683),
.A2(n_2659),
.B1(n_2595),
.B2(n_2593),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2700),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2714),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2712),
.Y(n_2729)
);

OAI21xp5_ASAP7_75t_L g2730 ( 
.A1(n_2711),
.A2(n_2584),
.B(n_2518),
.Y(n_2730)
);

AOI22xp5_ASAP7_75t_L g2731 ( 
.A1(n_2721),
.A2(n_2659),
.B1(n_2595),
.B2(n_2593),
.Y(n_2731)
);

OAI21xp33_ASAP7_75t_L g2732 ( 
.A1(n_2705),
.A2(n_2673),
.B(n_2582),
.Y(n_2732)
);

NAND2xp33_ASAP7_75t_SL g2733 ( 
.A(n_2707),
.B(n_2170),
.Y(n_2733)
);

OAI32xp33_ASAP7_75t_L g2734 ( 
.A1(n_2691),
.A2(n_2661),
.A3(n_2673),
.B1(n_2631),
.B2(n_2648),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2712),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2708),
.B(n_2677),
.Y(n_2736)
);

OAI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2698),
.A2(n_2518),
.B(n_2619),
.Y(n_2737)
);

AOI21xp5_ASAP7_75t_L g2738 ( 
.A1(n_2720),
.A2(n_2576),
.B(n_2574),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_SL g2739 ( 
.A(n_2695),
.B(n_2614),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2684),
.Y(n_2740)
);

OAI221xp5_ASAP7_75t_L g2741 ( 
.A1(n_2688),
.A2(n_2657),
.B1(n_2665),
.B2(n_2662),
.C(n_2606),
.Y(n_2741)
);

NOR2xp33_ASAP7_75t_L g2742 ( 
.A(n_2718),
.B(n_2233),
.Y(n_2742)
);

OAI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2715),
.A2(n_2698),
.B1(n_2708),
.B2(n_2687),
.Y(n_2743)
);

AOI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2709),
.A2(n_2582),
.B1(n_2616),
.B2(n_2525),
.Y(n_2744)
);

OAI21xp5_ASAP7_75t_L g2745 ( 
.A1(n_2685),
.A2(n_2619),
.B(n_2614),
.Y(n_2745)
);

OAI21xp33_ASAP7_75t_L g2746 ( 
.A1(n_2692),
.A2(n_2634),
.B(n_2583),
.Y(n_2746)
);

A2O1A1Ixp33_ASAP7_75t_L g2747 ( 
.A1(n_2694),
.A2(n_2351),
.B(n_2395),
.C(n_2256),
.Y(n_2747)
);

AOI21xp33_ASAP7_75t_L g2748 ( 
.A1(n_2686),
.A2(n_2273),
.B(n_2399),
.Y(n_2748)
);

AOI21xp5_ASAP7_75t_L g2749 ( 
.A1(n_2719),
.A2(n_2576),
.B(n_2574),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2689),
.Y(n_2750)
);

AOI32xp33_ASAP7_75t_L g2751 ( 
.A1(n_2693),
.A2(n_2669),
.A3(n_2377),
.B1(n_2525),
.B2(n_2552),
.Y(n_2751)
);

OAI21xp33_ASAP7_75t_L g2752 ( 
.A1(n_2724),
.A2(n_2719),
.B(n_2678),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_2742),
.B(n_2458),
.Y(n_2753)
);

INVxp67_ASAP7_75t_L g2754 ( 
.A(n_2733),
.Y(n_2754)
);

OAI222xp33_ASAP7_75t_L g2755 ( 
.A1(n_2741),
.A2(n_2679),
.B1(n_2676),
.B2(n_2696),
.C1(n_2717),
.C2(n_2677),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_SL g2756 ( 
.A(n_2743),
.B(n_2716),
.Y(n_2756)
);

AOI211xp5_ASAP7_75t_L g2757 ( 
.A1(n_2734),
.A2(n_2201),
.B(n_2213),
.C(n_2230),
.Y(n_2757)
);

A2O1A1Ixp33_ASAP7_75t_L g2758 ( 
.A1(n_2751),
.A2(n_2717),
.B(n_2696),
.C(n_2230),
.Y(n_2758)
);

NOR2x1_ASAP7_75t_SL g2759 ( 
.A(n_2739),
.B(n_2552),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2726),
.B(n_2687),
.Y(n_2760)
);

AOI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2738),
.A2(n_2716),
.B(n_2213),
.Y(n_2761)
);

OAI21xp5_ASAP7_75t_SL g2762 ( 
.A1(n_2747),
.A2(n_2306),
.B(n_2200),
.Y(n_2762)
);

AOI221xp5_ASAP7_75t_L g2763 ( 
.A1(n_2730),
.A2(n_2690),
.B1(n_2713),
.B2(n_2710),
.C(n_2703),
.Y(n_2763)
);

OAI21xp33_ASAP7_75t_SL g2764 ( 
.A1(n_2725),
.A2(n_2744),
.B(n_2745),
.Y(n_2764)
);

OAI221xp5_ASAP7_75t_L g2765 ( 
.A1(n_2737),
.A2(n_2702),
.B1(n_2579),
.B2(n_2645),
.C(n_2643),
.Y(n_2765)
);

NAND4xp25_ASAP7_75t_L g2766 ( 
.A(n_2748),
.B(n_2348),
.C(n_2319),
.D(n_2420),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2727),
.Y(n_2767)
);

AOI211xp5_ASAP7_75t_L g2768 ( 
.A1(n_2748),
.A2(n_2201),
.B(n_2283),
.C(n_2330),
.Y(n_2768)
);

NAND2xp33_ASAP7_75t_L g2769 ( 
.A(n_2749),
.B(n_2283),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2728),
.Y(n_2770)
);

AOI22x1_ASAP7_75t_L g2771 ( 
.A1(n_2723),
.A2(n_2438),
.B1(n_2307),
.B2(n_2565),
.Y(n_2771)
);

OAI21xp5_ASAP7_75t_SL g2772 ( 
.A1(n_2731),
.A2(n_2732),
.B(n_2736),
.Y(n_2772)
);

NOR2xp67_ASAP7_75t_L g2773 ( 
.A(n_2729),
.B(n_2680),
.Y(n_2773)
);

BUFx2_ASAP7_75t_L g2774 ( 
.A(n_2735),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2746),
.B(n_2568),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2740),
.B(n_2568),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2750),
.B(n_2573),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2726),
.B(n_2573),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2729),
.B(n_2597),
.Y(n_2779)
);

OAI211xp5_ASAP7_75t_L g2780 ( 
.A1(n_2724),
.A2(n_2305),
.B(n_2151),
.C(n_2349),
.Y(n_2780)
);

AOI211xp5_ASAP7_75t_L g2781 ( 
.A1(n_2724),
.A2(n_2330),
.B(n_2177),
.C(n_2612),
.Y(n_2781)
);

AOI211xp5_ASAP7_75t_L g2782 ( 
.A1(n_2780),
.A2(n_2177),
.B(n_2382),
.C(n_2373),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2754),
.Y(n_2783)
);

AOI221xp5_ASAP7_75t_SL g2784 ( 
.A1(n_2752),
.A2(n_1913),
.B1(n_2601),
.B2(n_2535),
.C(n_2528),
.Y(n_2784)
);

NOR4xp25_ASAP7_75t_L g2785 ( 
.A(n_2756),
.B(n_2501),
.C(n_2502),
.D(n_2491),
.Y(n_2785)
);

A2O1A1Ixp33_ASAP7_75t_L g2786 ( 
.A1(n_2754),
.A2(n_2365),
.B(n_2356),
.C(n_2610),
.Y(n_2786)
);

AOI211xp5_ASAP7_75t_L g2787 ( 
.A1(n_2762),
.A2(n_2382),
.B(n_2433),
.C(n_2426),
.Y(n_2787)
);

NOR3xp33_ASAP7_75t_L g2788 ( 
.A(n_2764),
.B(n_2261),
.C(n_2259),
.Y(n_2788)
);

AOI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2769),
.A2(n_2610),
.B1(n_2699),
.B2(n_2697),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2774),
.Y(n_2790)
);

NOR3xp33_ASAP7_75t_L g2791 ( 
.A(n_2755),
.B(n_2261),
.C(n_2259),
.Y(n_2791)
);

NAND3xp33_ASAP7_75t_L g2792 ( 
.A(n_2781),
.B(n_2757),
.C(n_2763),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_2761),
.B(n_2362),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2759),
.B(n_2617),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2767),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2770),
.Y(n_2796)
);

NOR3xp33_ASAP7_75t_L g2797 ( 
.A(n_2755),
.B(n_2772),
.C(n_2758),
.Y(n_2797)
);

OAI21xp5_ASAP7_75t_SL g2798 ( 
.A1(n_2760),
.A2(n_2565),
.B(n_2436),
.Y(n_2798)
);

OAI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_2771),
.A2(n_2251),
.B1(n_2362),
.B2(n_2356),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2778),
.B(n_2704),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2779),
.Y(n_2801)
);

AOI221xp5_ASAP7_75t_L g2802 ( 
.A1(n_2765),
.A2(n_2504),
.B1(n_2507),
.B2(n_2517),
.C(n_2521),
.Y(n_2802)
);

NOR3xp33_ASAP7_75t_L g2803 ( 
.A(n_2768),
.B(n_2268),
.C(n_2384),
.Y(n_2803)
);

NAND3xp33_ASAP7_75t_L g2804 ( 
.A(n_2797),
.B(n_2773),
.C(n_2753),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2783),
.B(n_2775),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_2785),
.B(n_2362),
.Y(n_2806)
);

NOR3xp33_ASAP7_75t_SL g2807 ( 
.A(n_2792),
.B(n_2766),
.C(n_2777),
.Y(n_2807)
);

NOR2x1_ASAP7_75t_L g2808 ( 
.A(n_2793),
.B(n_2365),
.Y(n_2808)
);

NAND4xp75_ASAP7_75t_L g2809 ( 
.A(n_2784),
.B(n_2776),
.C(n_2406),
.D(n_2419),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2790),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2801),
.Y(n_2811)
);

AOI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2788),
.A2(n_2798),
.B1(n_2791),
.B2(n_2789),
.Y(n_2812)
);

AOI21xp5_ASAP7_75t_L g2813 ( 
.A1(n_2786),
.A2(n_2362),
.B(n_2550),
.Y(n_2813)
);

NOR3xp33_ASAP7_75t_L g2814 ( 
.A(n_2795),
.B(n_2268),
.C(n_2384),
.Y(n_2814)
);

OAI211xp5_ASAP7_75t_L g2815 ( 
.A1(n_2787),
.A2(n_2346),
.B(n_2353),
.C(n_2319),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2802),
.B(n_2722),
.Y(n_2816)
);

NOR2x1_ASAP7_75t_SL g2817 ( 
.A(n_2799),
.B(n_2240),
.Y(n_2817)
);

INVx1_ASAP7_75t_SL g2818 ( 
.A(n_2796),
.Y(n_2818)
);

NAND3xp33_ASAP7_75t_L g2819 ( 
.A(n_2782),
.B(n_2228),
.C(n_2227),
.Y(n_2819)
);

INVx2_ASAP7_75t_SL g2820 ( 
.A(n_2794),
.Y(n_2820)
);

OAI322xp33_ASAP7_75t_L g2821 ( 
.A1(n_2800),
.A2(n_2548),
.A3(n_2529),
.B1(n_2544),
.B2(n_2551),
.C1(n_2495),
.C2(n_2505),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2810),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2807),
.B(n_2803),
.Y(n_2823)
);

NOR4xp75_ASAP7_75t_L g2824 ( 
.A(n_2805),
.B(n_2799),
.C(n_2598),
.D(n_2278),
.Y(n_2824)
);

NOR2x1p5_ASAP7_75t_L g2825 ( 
.A(n_2804),
.B(n_2429),
.Y(n_2825)
);

NAND3xp33_ASAP7_75t_L g2826 ( 
.A(n_2811),
.B(n_2564),
.C(n_2559),
.Y(n_2826)
);

NAND3xp33_ASAP7_75t_SL g2827 ( 
.A(n_2812),
.B(n_2238),
.C(n_2436),
.Y(n_2827)
);

NAND2x1p5_ASAP7_75t_L g2828 ( 
.A(n_2808),
.B(n_2429),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2818),
.Y(n_2829)
);

NOR4xp25_ASAP7_75t_L g2830 ( 
.A(n_2818),
.B(n_2815),
.C(n_2820),
.D(n_2821),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2809),
.A2(n_2612),
.B1(n_2587),
.B2(n_2589),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2817),
.B(n_2534),
.Y(n_2832)
);

INVx2_ASAP7_75t_SL g2833 ( 
.A(n_2816),
.Y(n_2833)
);

NAND4xp25_ASAP7_75t_L g2834 ( 
.A(n_2806),
.B(n_2452),
.C(n_2312),
.D(n_2364),
.Y(n_2834)
);

NAND3xp33_ASAP7_75t_L g2835 ( 
.A(n_2819),
.B(n_2481),
.C(n_2467),
.Y(n_2835)
);

NOR2xp67_ASAP7_75t_SL g2836 ( 
.A(n_2829),
.B(n_2813),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2823),
.A2(n_2833),
.B1(n_2825),
.B2(n_2830),
.Y(n_2837)
);

NOR2x1_ASAP7_75t_L g2838 ( 
.A(n_2822),
.B(n_2834),
.Y(n_2838)
);

AND2x2_ASAP7_75t_SL g2839 ( 
.A(n_2832),
.B(n_2814),
.Y(n_2839)
);

NAND4xp75_ASAP7_75t_L g2840 ( 
.A(n_2824),
.B(n_2530),
.C(n_2546),
.D(n_2527),
.Y(n_2840)
);

AO22x2_ASAP7_75t_L g2841 ( 
.A1(n_2827),
.A2(n_2452),
.B1(n_2312),
.B2(n_2364),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2826),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2835),
.Y(n_2843)
);

NOR2x1_ASAP7_75t_L g2844 ( 
.A(n_2831),
.B(n_2304),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2828),
.B(n_2618),
.Y(n_2845)
);

OAI22xp33_ASAP7_75t_L g2846 ( 
.A1(n_2823),
.A2(n_2304),
.B1(n_2309),
.B2(n_2613),
.Y(n_2846)
);

INVx2_ASAP7_75t_SL g2847 ( 
.A(n_2844),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2842),
.B(n_2672),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2843),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2839),
.Y(n_2850)
);

NAND3xp33_ASAP7_75t_L g2851 ( 
.A(n_2837),
.B(n_2309),
.C(n_2304),
.Y(n_2851)
);

NOR2x1_ASAP7_75t_L g2852 ( 
.A(n_2838),
.B(n_2309),
.Y(n_2852)
);

XNOR2x1_ASAP7_75t_L g2853 ( 
.A(n_2840),
.B(n_2369),
.Y(n_2853)
);

OR2x2_ASAP7_75t_L g2854 ( 
.A(n_2845),
.B(n_2578),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2846),
.B(n_2672),
.Y(n_2855)
);

AO21x2_ASAP7_75t_L g2856 ( 
.A1(n_2849),
.A2(n_2836),
.B(n_2841),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2848),
.Y(n_2857)
);

OAI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2851),
.A2(n_2481),
.B1(n_2498),
.B2(n_2495),
.Y(n_2858)
);

XNOR2xp5_ASAP7_75t_L g2859 ( 
.A(n_2853),
.B(n_2238),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2847),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2860),
.Y(n_2861)
);

OAI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2861),
.A2(n_2850),
.B1(n_2857),
.B2(n_2859),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2862),
.Y(n_2863)
);

AO21x2_ASAP7_75t_L g2864 ( 
.A1(n_2863),
.A2(n_2857),
.B(n_2856),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2864),
.B(n_2852),
.Y(n_2865)
);

OR2x6_ASAP7_75t_L g2866 ( 
.A(n_2865),
.B(n_2854),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_SL g2867 ( 
.A1(n_2866),
.A2(n_2855),
.B1(n_2858),
.B2(n_2369),
.Y(n_2867)
);


endmodule