module real_aes_13488_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_0), .B(n_10), .C(n_21), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g43 ( .A(n_1), .Y(n_43) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_2), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g37 ( .A(n_2), .B(n_38), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_3), .Y(n_28) );
NAND2xp33_ASAP7_75t_R g29 ( .A(n_3), .B(n_14), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_3), .B(n_14), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g34 ( .A(n_3), .B(n_35), .Y(n_34) );
OAI22xp33_ASAP7_75t_SL g30 ( .A1(n_4), .A2(n_13), .B1(n_31), .B2(n_33), .Y(n_30) );
NAND5xp2_ASAP7_75t_SL g17 ( .A(n_5), .B(n_9), .C(n_18), .D(n_23), .E(n_24), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_5), .Y(n_39) );
OAI22xp33_ASAP7_75t_SL g25 ( .A1(n_6), .A2(n_8), .B1(n_26), .B2(n_29), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g41 ( .A(n_7), .Y(n_41) );
NOR2xp33_ASAP7_75t_R g40 ( .A(n_9), .B(n_19), .Y(n_40) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_11), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_12), .Y(n_24) );
NAND3xp33_ASAP7_75t_SL g38 ( .A(n_12), .B(n_39), .C(n_40), .Y(n_38) );
NOR2xp33_ASAP7_75t_R g27 ( .A(n_14), .B(n_28), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_14), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_15), .Y(n_21) );
OAI322xp33_ASAP7_75t_L g16 ( .A1(n_17), .A2(n_25), .A3(n_30), .B1(n_36), .B2(n_41), .C1(n_42), .C2(n_43), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
NAND2xp33_ASAP7_75t_R g19 ( .A(n_20), .B(n_22), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_27), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_32), .Y(n_31) );
NAND2xp33_ASAP7_75t_R g36 ( .A(n_32), .B(n_37), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_34), .Y(n_33) );
NAND2xp33_ASAP7_75t_R g42 ( .A(n_34), .B(n_37), .Y(n_42) );
endmodule