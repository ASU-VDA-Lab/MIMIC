module fake_jpeg_32051_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_11),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx8_ASAP7_75t_SL g57 ( 
.A(n_5),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_60),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_20),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_55),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_55),
.B(n_60),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_43),
.B(n_46),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_78),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_55),
.B1(n_58),
.B2(n_44),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_81),
.B1(n_56),
.B2(n_2),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_58),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_73),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_51),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_93),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_39),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_53),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_74),
.B1(n_53),
.B2(n_41),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_96),
.B1(n_97),
.B2(n_6),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_42),
.B1(n_54),
.B2(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_21),
.B1(n_37),
.B2(n_36),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_100),
.B1(n_108),
.B2(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_115),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_114),
.B1(n_15),
.B2(n_16),
.Y(n_124)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_31),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_23),
.B1(n_33),
.B2(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_8),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_9),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_35),
.B1(n_22),
.B2(n_13),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_10),
.B(n_12),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_120),
.C(n_125),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_103),
.C(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_111),
.B(n_12),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_122),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_14),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_124),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_17),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_127),
.B1(n_102),
.B2(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_130),
.C(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_125),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_135),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_137),
.C(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_137),
.C(n_108),
.Y(n_143)
);

AOI221xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_127),
.B1(n_104),
.B2(n_131),
.C(n_128),
.Y(n_144)
);


endmodule