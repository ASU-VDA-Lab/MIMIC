module real_aes_1069_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_0), .B(n_217), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_1), .A2(n_200), .B(n_250), .Y(n_249) );
AO22x2_ASAP7_75t_L g87 ( .A1(n_2), .A2(n_54), .B1(n_88), .B2(n_89), .Y(n_87) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_3), .B(n_207), .Y(n_263) );
INVx1_ASAP7_75t_L g183 ( .A(n_4), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_5), .B(n_207), .Y(n_227) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_6), .A2(n_25), .B1(n_88), .B2(n_92), .Y(n_91) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_7), .A2(n_24), .B1(n_153), .B2(n_155), .Y(n_152) );
AOI22xp5_ASAP7_75t_SL g138 ( .A1(n_8), .A2(n_62), .B1(n_139), .B2(n_141), .Y(n_138) );
NAND2xp33_ASAP7_75t_L g244 ( .A(n_9), .B(n_211), .Y(n_244) );
INVx2_ASAP7_75t_L g197 ( .A(n_10), .Y(n_197) );
AOI221x1_ASAP7_75t_L g286 ( .A1(n_11), .A2(n_20), .B1(n_200), .B2(n_217), .C(n_287), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_12), .A2(n_52), .B1(n_107), .B2(n_115), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_13), .B(n_217), .Y(n_240) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_14), .A2(n_238), .B(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_15), .B(n_230), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_16), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_17), .B(n_134), .Y(n_133) );
AO21x1_ASAP7_75t_L g258 ( .A1(n_18), .A2(n_217), .B(n_259), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_19), .A2(n_71), .B1(n_168), .B2(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g169 ( .A(n_19), .Y(n_169) );
NAND2x1_ASAP7_75t_L g272 ( .A(n_21), .B(n_207), .Y(n_272) );
NAND2x1_ASAP7_75t_L g226 ( .A(n_22), .B(n_211), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_23), .A2(n_80), .B1(n_81), .B2(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_23), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g175 ( .A1(n_25), .A2(n_54), .B1(n_58), .B2(n_176), .C(n_178), .Y(n_175) );
OR2x2_ASAP7_75t_L g196 ( .A(n_26), .B(n_65), .Y(n_196) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_26), .A2(n_65), .B(n_197), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_27), .B(n_211), .Y(n_252) );
INVx3_ASAP7_75t_L g88 ( .A(n_28), .Y(n_88) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_29), .B(n_207), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_30), .A2(n_64), .B1(n_119), .B2(n_122), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_31), .B(n_211), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_32), .A2(n_47), .B1(n_126), .B2(n_130), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g83 ( .A1(n_33), .A2(n_40), .B1(n_84), .B2(n_101), .Y(n_83) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_34), .A2(n_200), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g99 ( .A(n_35), .Y(n_99) );
INVx1_ASAP7_75t_L g185 ( .A(n_36), .Y(n_185) );
AND2x2_ASAP7_75t_L g201 ( .A(n_36), .B(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g215 ( .A(n_36), .B(n_183), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_37), .B(n_217), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_37), .A2(n_80), .B1(n_81), .B2(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_37), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_38), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_39), .B(n_211), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_41), .A2(n_80), .B1(n_81), .B2(n_160), .Y(n_79) );
INVx1_ASAP7_75t_L g160 ( .A(n_41), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_42), .A2(n_200), .B(n_225), .Y(n_224) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_43), .A2(n_58), .B1(n_88), .B2(n_95), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_44), .B(n_211), .Y(n_273) );
INVx1_ASAP7_75t_L g204 ( .A(n_45), .Y(n_204) );
INVx1_ASAP7_75t_L g213 ( .A(n_45), .Y(n_213) );
INVx1_ASAP7_75t_L g100 ( .A(n_46), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_48), .B(n_207), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_49), .A2(n_200), .B(n_271), .Y(n_270) );
AO21x1_ASAP7_75t_L g260 ( .A1(n_50), .A2(n_200), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_51), .B(n_217), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_53), .B(n_217), .Y(n_228) );
INVxp33_ASAP7_75t_L g180 ( .A(n_54), .Y(n_180) );
AND2x2_ASAP7_75t_L g309 ( .A(n_55), .B(n_231), .Y(n_309) );
INVx1_ASAP7_75t_L g202 ( .A(n_56), .Y(n_202) );
INVx1_ASAP7_75t_L g209 ( .A(n_56), .Y(n_209) );
AND2x2_ASAP7_75t_L g232 ( .A(n_57), .B(n_233), .Y(n_232) );
INVxp67_ASAP7_75t_L g179 ( .A(n_58), .Y(n_179) );
INVx1_ASAP7_75t_L g163 ( .A(n_59), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_59), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g246 ( .A(n_60), .B(n_233), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_61), .A2(n_69), .B1(n_146), .B2(n_148), .Y(n_145) );
AND2x2_ASAP7_75t_L g259 ( .A(n_63), .B(n_195), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_66), .B(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g276 ( .A(n_67), .B(n_233), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_68), .B(n_207), .Y(n_307) );
INVx1_ASAP7_75t_L g529 ( .A(n_68), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_70), .A2(n_200), .B(n_205), .Y(n_199) );
INVx1_ASAP7_75t_L g168 ( .A(n_71), .Y(n_168) );
INVx1_ASAP7_75t_L g171 ( .A(n_72), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_73), .B(n_211), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_74), .B(n_207), .Y(n_251) );
BUFx2_ASAP7_75t_SL g177 ( .A(n_75), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_76), .A2(n_200), .B(n_242), .Y(n_241) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_172), .B1(n_186), .B2(n_503), .C(n_509), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_161), .Y(n_78) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_81), .Y(n_80) );
OR2x2_ASAP7_75t_L g81 ( .A(n_82), .B(n_132), .Y(n_81) );
NAND4xp25_ASAP7_75t_L g82 ( .A(n_83), .B(n_106), .C(n_118), .D(n_125), .Y(n_82) );
BUFx6f_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_93), .Y(n_85) );
AND2x4_ASAP7_75t_L g124 ( .A(n_86), .B(n_113), .Y(n_124) );
AND2x2_ASAP7_75t_L g154 ( .A(n_86), .B(n_129), .Y(n_154) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_90), .Y(n_86) );
AND2x2_ASAP7_75t_L g105 ( .A(n_87), .B(n_91), .Y(n_105) );
INVx2_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
INVx1_ASAP7_75t_L g89 ( .A(n_88), .Y(n_89) );
INVx2_ASAP7_75t_L g92 ( .A(n_88), .Y(n_92) );
INVx1_ASAP7_75t_L g95 ( .A(n_88), .Y(n_95) );
OAI22x1_ASAP7_75t_L g97 ( .A1(n_88), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_88), .Y(n_98) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_90), .Y(n_159) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g111 ( .A(n_91), .Y(n_111) );
AND2x4_ASAP7_75t_L g117 ( .A(n_91), .B(n_112), .Y(n_117) );
AND2x2_ASAP7_75t_L g121 ( .A(n_93), .B(n_110), .Y(n_121) );
AND2x4_ASAP7_75t_L g140 ( .A(n_93), .B(n_117), .Y(n_140) );
AND2x2_ASAP7_75t_L g93 ( .A(n_94), .B(n_96), .Y(n_93) );
BUFx2_ASAP7_75t_L g104 ( .A(n_94), .Y(n_104) );
INVx2_ASAP7_75t_L g114 ( .A(n_94), .Y(n_114) );
AND2x2_ASAP7_75t_L g137 ( .A(n_94), .B(n_97), .Y(n_137) );
AND2x4_ASAP7_75t_L g113 ( .A(n_96), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g129 ( .A(n_97), .B(n_114), .Y(n_129) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_97), .Y(n_151) );
INVx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx5_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x4_ASAP7_75t_L g131 ( .A(n_105), .B(n_113), .Y(n_131) );
AND2x2_ASAP7_75t_L g150 ( .A(n_105), .B(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx8_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_113), .Y(n_109) );
AND2x4_ASAP7_75t_L g128 ( .A(n_110), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g136 ( .A(n_110), .B(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVxp67_ASAP7_75t_L g144 ( .A(n_112), .Y(n_144) );
AND2x4_ASAP7_75t_L g116 ( .A(n_113), .B(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g147 ( .A(n_117), .B(n_129), .Y(n_147) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx8_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx6_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND4xp25_ASAP7_75t_SL g132 ( .A(n_133), .B(n_138), .C(n_145), .D(n_152), .Y(n_132) );
INVx4_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx6_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g143 ( .A(n_137), .B(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g157 ( .A(n_137), .B(n_158), .Y(n_157) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx6_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B1(n_164), .B2(n_165), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g165 ( .A1(n_166), .A2(n_167), .B1(n_170), .B2(n_171), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
AND3x1_ASAP7_75t_SL g174 ( .A(n_175), .B(n_181), .C(n_184), .Y(n_174) );
INVxp67_ASAP7_75t_L g517 ( .A(n_175), .Y(n_517) );
CKINVDCx8_ASAP7_75t_R g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_181), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_181), .A2(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OR2x2_ASAP7_75t_SL g522 ( .A(n_182), .B(n_184), .Y(n_522) );
AND2x2_ASAP7_75t_L g527 ( .A(n_182), .B(n_528), .Y(n_527) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g203 ( .A(n_183), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_184), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2x1p5_ASAP7_75t_L g506 ( .A(n_185), .B(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_401), .Y(n_187) );
NAND3xp33_ASAP7_75t_SL g188 ( .A(n_189), .B(n_313), .C(n_368), .Y(n_188) );
AOI221xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_253), .B1(n_277), .B2(n_281), .C(n_291), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_236), .Y(n_190) );
AND2x2_ASAP7_75t_SL g279 ( .A(n_191), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g312 ( .A(n_191), .Y(n_312) );
AND2x2_ASAP7_75t_L g357 ( .A(n_191), .B(n_294), .Y(n_357) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_221), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g345 ( .A(n_193), .Y(n_345) );
INVx1_ASAP7_75t_L g355 ( .A(n_193), .Y(n_355) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_198), .B(n_219), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_194), .B(n_220), .Y(n_219) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_194), .A2(n_198), .B(n_219), .Y(n_319) );
INVx1_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_195), .A2(n_240), .B(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_195), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
AND2x2_ASAP7_75t_SL g231 ( .A(n_196), .B(n_197), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_216), .Y(n_198) );
AND2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_203), .Y(n_200) );
AND2x6_ASAP7_75t_L g211 ( .A(n_202), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g508 ( .A(n_202), .Y(n_508) );
AND2x4_ASAP7_75t_L g505 ( .A(n_203), .B(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g207 ( .A(n_204), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g528 ( .A(n_204), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_210), .B(n_214), .Y(n_205) );
AND2x4_ASAP7_75t_L g218 ( .A(n_208), .B(n_212), .Y(n_218) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_214), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_214), .A2(n_243), .B(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_214), .A2(n_251), .B(n_252), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_214), .A2(n_262), .B(n_263), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_214), .A2(n_272), .B(n_273), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_214), .A2(n_288), .B(n_289), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_214), .A2(n_306), .B(n_307), .Y(n_305) );
INVx5_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g217 ( .A(n_215), .B(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g334 ( .A(n_221), .B(n_237), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_221), .B(n_280), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_221), .B(n_245), .Y(n_378) );
INVx2_ASAP7_75t_L g387 ( .A(n_221), .Y(n_387) );
AND2x2_ASAP7_75t_L g408 ( .A(n_221), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g492 ( .A(n_221), .B(n_311), .Y(n_492) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g320 ( .A(n_222), .B(n_245), .Y(n_320) );
AND2x2_ASAP7_75t_L g453 ( .A(n_222), .B(n_280), .Y(n_453) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_222), .Y(n_479) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_232), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_228), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_230), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_230), .A2(n_248), .B(n_249), .Y(n_247) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_230), .A2(n_286), .B(n_290), .Y(n_285) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_230), .A2(n_286), .B(n_290), .Y(n_297) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g275 ( .A(n_233), .Y(n_275) );
INVx4_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
BUFx4f_ASAP7_75t_L g238 ( .A(n_235), .Y(n_238) );
AND2x4_ASAP7_75t_L g407 ( .A(n_236), .B(n_408), .Y(n_407) );
AOI321xp33_ASAP7_75t_L g421 ( .A1(n_236), .A2(n_350), .A3(n_351), .B1(n_383), .B2(n_422), .C(n_425), .Y(n_421) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_245), .Y(n_236) );
BUFx3_ASAP7_75t_L g278 ( .A(n_237), .Y(n_278) );
INVx2_ASAP7_75t_L g311 ( .A(n_237), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_237), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g344 ( .A(n_237), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g377 ( .A(n_237), .Y(n_377) );
INVx5_ASAP7_75t_L g280 ( .A(n_245), .Y(n_280) );
NOR2x1_ASAP7_75t_SL g329 ( .A(n_245), .B(n_319), .Y(n_329) );
BUFx2_ASAP7_75t_L g424 ( .A(n_245), .Y(n_424) );
OR2x6_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVxp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_266), .Y(n_254) );
NOR2xp33_ASAP7_75t_SL g322 ( .A(n_255), .B(n_323), .Y(n_322) );
NOR4xp25_ASAP7_75t_L g425 ( .A(n_255), .B(n_419), .C(n_423), .D(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g463 ( .A(n_255), .Y(n_463) );
AND2x2_ASAP7_75t_L g497 ( .A(n_255), .B(n_437), .Y(n_497) );
BUFx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g298 ( .A(n_256), .Y(n_298) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g352 ( .A(n_257), .Y(n_352) );
OAI21x1_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_260), .B(n_264), .Y(n_257) );
INVx1_ASAP7_75t_L g265 ( .A(n_259), .Y(n_265) );
AOI33xp33_ASAP7_75t_L g493 ( .A1(n_266), .A2(n_295), .A3(n_326), .B1(n_342), .B2(n_448), .B3(n_494), .Y(n_493) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g283 ( .A(n_267), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g293 ( .A(n_267), .B(n_294), .Y(n_293) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g300 ( .A(n_268), .Y(n_300) );
INVxp67_ASAP7_75t_L g381 ( .A(n_268), .Y(n_381) );
AND2x2_ASAP7_75t_L g437 ( .A(n_268), .B(n_302), .Y(n_437) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_275), .B(n_276), .Y(n_268) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_269), .A2(n_275), .B(n_276), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_275), .A2(n_303), .B(n_309), .Y(n_302) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_275), .A2(n_303), .B(n_309), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_277), .A2(n_459), .B(n_460), .Y(n_458) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g446 ( .A(n_278), .B(n_320), .Y(n_446) );
AND3x2_ASAP7_75t_L g448 ( .A(n_278), .B(n_332), .C(n_387), .Y(n_448) );
INVx3_ASAP7_75t_SL g400 ( .A(n_279), .Y(n_400) );
INVx4_ASAP7_75t_L g294 ( .A(n_280), .Y(n_294) );
AND2x2_ASAP7_75t_L g332 ( .A(n_280), .B(n_319), .Y(n_332) );
INVxp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g326 ( .A(n_284), .Y(n_326) );
AND2x4_ASAP7_75t_L g351 ( .A(n_284), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g414 ( .A(n_284), .B(n_302), .Y(n_414) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g384 ( .A(n_285), .Y(n_384) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_285), .Y(n_406) );
O2A1O1Ixp33_ASAP7_75t_R g291 ( .A1(n_292), .A2(n_295), .B(n_299), .C(n_310), .Y(n_291) );
CKINVDCx16_ASAP7_75t_R g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g343 ( .A(n_294), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_294), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_294), .B(n_311), .Y(n_472) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g454 ( .A(n_296), .B(n_444), .Y(n_454) );
AND2x2_ASAP7_75t_SL g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g301 ( .A(n_297), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g323 ( .A(n_297), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g339 ( .A(n_297), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g372 ( .A(n_297), .B(n_352), .Y(n_372) );
AND2x4_ASAP7_75t_L g337 ( .A(n_298), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g361 ( .A(n_298), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g399 ( .A(n_298), .B(n_324), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g327 ( .A(n_300), .B(n_324), .Y(n_327) );
AND2x2_ASAP7_75t_L g342 ( .A(n_300), .B(n_302), .Y(n_342) );
BUFx2_ASAP7_75t_L g398 ( .A(n_300), .Y(n_398) );
AND2x2_ASAP7_75t_L g412 ( .A(n_300), .B(n_323), .Y(n_412) );
INVx2_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_304), .B(n_308), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_310), .A2(n_361), .B1(n_363), .B2(n_367), .Y(n_360) );
INVx2_ASAP7_75t_SL g391 ( .A(n_310), .Y(n_391) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AND2x2_ASAP7_75t_L g366 ( .A(n_311), .B(n_319), .Y(n_366) );
INVx1_ASAP7_75t_L g473 ( .A(n_312), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_346), .C(n_360), .Y(n_313) );
OAI221xp5_ASAP7_75t_SL g314 ( .A1(n_315), .A2(n_321), .B1(n_325), .B2(n_328), .C(n_330), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_320), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g374 ( .A(n_318), .Y(n_374) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_318), .Y(n_502) );
INVx1_ASAP7_75t_L g465 ( .A(n_320), .Y(n_465) );
AND2x2_ASAP7_75t_SL g475 ( .A(n_320), .B(n_344), .Y(n_475) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_324), .B(n_352), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OR2x2_ASAP7_75t_L g358 ( .A(n_326), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g436 ( .A(n_326), .Y(n_436) );
AND2x2_ASAP7_75t_L g371 ( .A(n_327), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g417 ( .A(n_329), .B(n_377), .Y(n_417) );
AND2x2_ASAP7_75t_L g494 ( .A(n_329), .B(n_492), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B1(n_342), .B2(n_343), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g353 ( .A(n_334), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx2_ASAP7_75t_L g359 ( .A(n_337), .Y(n_359) );
AND2x4_ASAP7_75t_L g383 ( .A(n_337), .B(n_384), .Y(n_383) );
OAI21xp33_ASAP7_75t_SL g413 ( .A1(n_337), .A2(n_414), .B(n_415), .Y(n_413) );
AND2x2_ASAP7_75t_L g440 ( .A(n_337), .B(n_398), .Y(n_440) );
INVx2_ASAP7_75t_L g362 ( .A(n_338), .Y(n_362) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_338), .Y(n_395) );
INVx1_ASAP7_75t_SL g419 ( .A(n_339), .Y(n_419) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g350 ( .A(n_341), .Y(n_350) );
AND2x4_ASAP7_75t_SL g444 ( .A(n_341), .B(n_362), .Y(n_444) );
AND2x2_ASAP7_75t_L g441 ( .A(n_344), .B(n_387), .Y(n_441) );
AND2x2_ASAP7_75t_L g467 ( .A(n_344), .B(n_453), .Y(n_467) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_345), .Y(n_389) );
INVx1_ASAP7_75t_L g409 ( .A(n_345), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_353), .B1(n_356), .B2(n_358), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_351), .B(n_362), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_351), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g490 ( .A(n_351), .Y(n_490) );
INVx2_ASAP7_75t_SL g415 ( .A(n_353), .Y(n_415) );
AND2x2_ASAP7_75t_L g427 ( .A(n_355), .B(n_387), .Y(n_427) );
INVx2_ASAP7_75t_L g433 ( .A(n_355), .Y(n_433) );
INVxp33_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_361), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g483 ( .A(n_361), .Y(n_483) );
INVx1_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_364), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g422 ( .A(n_366), .B(n_423), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_366), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_390), .C(n_393), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B1(n_375), .B2(n_379), .C(n_382), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_SL g488 ( .A(n_373), .Y(n_488) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g457 ( .A(n_374), .B(n_423), .Y(n_457) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g388 ( .A(n_377), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g459 ( .A(n_379), .Y(n_459) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g456 ( .A(n_380), .Y(n_456) );
INVx1_ASAP7_75t_L g462 ( .A(n_381), .Y(n_462) );
OR2x2_ASAP7_75t_L g485 ( .A(n_381), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_SL g394 ( .A(n_384), .Y(n_394) );
AND2x2_ASAP7_75t_L g464 ( .A(n_384), .B(n_444), .Y(n_464) );
AND2x2_ASAP7_75t_SL g496 ( .A(n_384), .B(n_397), .Y(n_496) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g501 ( .A(n_387), .Y(n_501) );
INVx1_ASAP7_75t_L g451 ( .A(n_389), .Y(n_451) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_396), .C(n_400), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_394), .B(n_444), .Y(n_468) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_397), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
AND2x2_ASAP7_75t_L g405 ( .A(n_399), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g486 ( .A(n_399), .Y(n_486) );
NAND4xp75_ASAP7_75t_L g401 ( .A(n_402), .B(n_458), .C(n_474), .D(n_495), .Y(n_401) );
NOR3x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_420), .C(n_442), .Y(n_402) );
NAND4xp75_ASAP7_75t_L g403 ( .A(n_404), .B(n_410), .C(n_413), .D(n_416), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_405), .B(n_407), .Y(n_404) );
AND2x2_ASAP7_75t_L g455 ( .A(n_406), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_SL g480 ( .A(n_407), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_SL g469 ( .A(n_412), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_428), .Y(n_420) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_424), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_434), .B(n_438), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI322xp33_ASAP7_75t_L g460 ( .A1(n_432), .A2(n_461), .A3(n_465), .B1(n_466), .B2(n_468), .C1(n_469), .C2(n_470), .Y(n_460) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_433), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_436), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_437), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_445), .B(n_447), .C(n_449), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_454), .B1(n_455), .B2(n_457), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_464), .Y(n_461) );
INVxp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_467), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g477 ( .A(n_472), .B(n_478), .Y(n_477) );
O2A1O1Ixp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_481), .C(n_484), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_477), .B(n_480), .Y(n_476) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_SL g484 ( .A1(n_485), .A2(n_487), .B1(n_489), .B2(n_491), .C(n_493), .Y(n_484) );
INVxp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_506), .Y(n_525) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI222xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .B1(n_518), .B2(n_520), .C1(n_523), .C2(n_529), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
endmodule