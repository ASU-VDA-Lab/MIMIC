module real_aes_6189_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g250 ( .A1(n_0), .A2(n_251), .B(n_252), .C(n_255), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_1), .B(n_192), .Y(n_256) );
INVx1_ASAP7_75t_L g430 ( .A(n_2), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_3), .B(n_162), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_4), .A2(n_132), .B(n_135), .C(n_471), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_5), .A2(n_152), .B(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_6), .A2(n_152), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_7), .B(n_192), .Y(n_517) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_8), .A2(n_119), .B(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_9), .A2(n_451), .B1(n_454), .B2(n_455), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_9), .Y(n_455) );
AND2x6_ASAP7_75t_L g132 ( .A(n_10), .B(n_133), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_11), .A2(n_132), .B(n_135), .C(n_138), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_12), .A2(n_47), .B1(n_452), .B2(n_453), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_12), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_13), .B(n_42), .Y(n_431) );
INVx1_ASAP7_75t_L g487 ( .A(n_14), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_15), .B(n_142), .Y(n_473) );
INVx1_ASAP7_75t_L g124 ( .A(n_16), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_17), .B(n_162), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_18), .A2(n_140), .B(n_495), .C(n_497), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_19), .B(n_192), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_20), .B(n_216), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_21), .A2(n_135), .B(n_179), .C(n_212), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_22), .A2(n_144), .B(n_254), .C(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_23), .B(n_142), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_24), .B(n_142), .Y(n_538) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_25), .Y(n_545) );
INVx1_ASAP7_75t_L g537 ( .A(n_26), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_27), .A2(n_135), .B(n_175), .C(n_179), .Y(n_174) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_28), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_29), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_30), .B(n_435), .Y(n_436) );
INVx1_ASAP7_75t_L g528 ( .A(n_31), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_32), .A2(n_152), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g130 ( .A(n_33), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_34), .A2(n_154), .B(n_165), .C(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_35), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_36), .A2(n_254), .B(n_514), .C(n_516), .Y(n_513) );
INVxp67_ASAP7_75t_L g529 ( .A(n_37), .Y(n_529) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_38), .A2(n_103), .B1(n_437), .B2(n_445), .C1(n_448), .C2(n_738), .Y(n_102) );
OAI321xp33_ASAP7_75t_L g103 ( .A1(n_38), .A2(n_104), .A3(n_426), .B1(n_432), .B2(n_433), .C(n_436), .Y(n_103) );
INVx1_ASAP7_75t_L g432 ( .A(n_38), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_39), .B(n_177), .Y(n_176) );
CKINVDCx14_ASAP7_75t_R g512 ( .A(n_40), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_41), .A2(n_135), .B(n_179), .C(n_536), .Y(n_535) );
AOI222xp33_ASAP7_75t_SL g449 ( .A1(n_43), .A2(n_450), .B1(n_456), .B2(n_730), .C1(n_731), .C2(n_735), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_44), .A2(n_255), .B(n_485), .C(n_486), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_45), .B(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_46), .Y(n_147) );
INVx1_ASAP7_75t_L g453 ( .A(n_47), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_48), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_49), .B(n_152), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_50), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_51), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_52), .A2(n_154), .B(n_156), .C(n_165), .Y(n_153) );
INVx1_ASAP7_75t_L g253 ( .A(n_53), .Y(n_253) );
INVx1_ASAP7_75t_L g157 ( .A(n_54), .Y(n_157) );
INVx1_ASAP7_75t_L g502 ( .A(n_55), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_56), .B(n_152), .Y(n_151) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_57), .A2(n_60), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_57), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_58), .Y(n_219) );
CKINVDCx14_ASAP7_75t_R g483 ( .A(n_59), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_60), .Y(n_107) );
INVx1_ASAP7_75t_L g133 ( .A(n_61), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_62), .B(n_152), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_63), .B(n_192), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_64), .A2(n_186), .B(n_188), .C(n_190), .Y(n_185) );
INVx1_ASAP7_75t_L g123 ( .A(n_65), .Y(n_123) );
INVx1_ASAP7_75t_SL g515 ( .A(n_66), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_67), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_68), .B(n_162), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_69), .B(n_192), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_70), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g548 ( .A(n_71), .Y(n_548) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_72), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_73), .B(n_159), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_74), .A2(n_135), .B(n_165), .C(n_226), .Y(n_225) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_75), .Y(n_184) );
INVx1_ASAP7_75t_L g444 ( .A(n_76), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_77), .A2(n_152), .B(n_482), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_78), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_79), .A2(n_152), .B(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_80), .A2(n_210), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g493 ( .A(n_81), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_82), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_83), .B(n_158), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_84), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_85), .A2(n_152), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g496 ( .A(n_86), .Y(n_496) );
INVx2_ASAP7_75t_L g121 ( .A(n_87), .Y(n_121) );
INVx1_ASAP7_75t_L g472 ( .A(n_88), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_89), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_90), .B(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g427 ( .A(n_91), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g459 ( .A(n_91), .B(n_429), .Y(n_459) );
INVx2_ASAP7_75t_L g729 ( .A(n_91), .Y(n_729) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_92), .A2(n_135), .B(n_165), .C(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_93), .B(n_152), .Y(n_198) );
INVx1_ASAP7_75t_L g201 ( .A(n_94), .Y(n_201) );
INVxp67_ASAP7_75t_L g189 ( .A(n_95), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_96), .B(n_119), .Y(n_488) );
INVx1_ASAP7_75t_L g126 ( .A(n_97), .Y(n_126) );
INVx1_ASAP7_75t_L g227 ( .A(n_98), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_99), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g505 ( .A(n_100), .Y(n_505) );
AND2x2_ASAP7_75t_L g168 ( .A(n_101), .B(n_167), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_104), .B(n_434), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_106), .B1(n_109), .B2(n_110), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22x1_ASAP7_75t_SL g731 ( .A1(n_109), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g456 ( .A1(n_110), .A2(n_457), .B1(n_460), .B2(n_726), .Y(n_456) );
OR3x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_324), .C(n_389), .Y(n_110) );
NAND4xp25_ASAP7_75t_SL g111 ( .A(n_112), .B(n_265), .C(n_291), .D(n_314), .Y(n_111) );
AOI221xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_193), .B1(n_234), .B2(n_241), .C(n_257), .Y(n_112) );
CKINVDCx14_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_114), .A2(n_258), .B1(n_282), .B2(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_169), .Y(n_114) );
INVx1_ASAP7_75t_SL g318 ( .A(n_115), .Y(n_318) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_149), .Y(n_115) );
OR2x2_ASAP7_75t_L g239 ( .A(n_116), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g260 ( .A(n_116), .B(n_170), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_116), .B(n_180), .Y(n_273) );
AND2x2_ASAP7_75t_L g290 ( .A(n_116), .B(n_149), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_116), .B(n_237), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_116), .B(n_289), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_116), .B(n_169), .Y(n_411) );
AOI211xp5_ASAP7_75t_SL g422 ( .A1(n_116), .A2(n_328), .B(n_423), .C(n_424), .Y(n_422) );
INVx5_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_117), .B(n_170), .Y(n_294) );
AND2x2_ASAP7_75t_L g297 ( .A(n_117), .B(n_171), .Y(n_297) );
OR2x2_ASAP7_75t_L g342 ( .A(n_117), .B(n_170), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_117), .B(n_180), .Y(n_351) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_125), .B(n_146), .Y(n_117) );
INVx3_ASAP7_75t_L g192 ( .A(n_118), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_118), .B(n_204), .Y(n_203) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_118), .A2(n_224), .B(n_232), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_118), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_118), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_118), .B(n_540), .Y(n_539) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_118), .A2(n_544), .B(n_550), .Y(n_543) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_119), .A2(n_173), .B(n_174), .Y(n_172) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_119), .Y(n_181) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_121), .B(n_122), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B(n_134), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_127), .A2(n_469), .B(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_127), .A2(n_167), .B(n_534), .C(n_535), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_127), .A2(n_545), .B(n_546), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
AND2x4_ASAP7_75t_L g152 ( .A(n_128), .B(n_132), .Y(n_152) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx1_ASAP7_75t_L g145 ( .A(n_130), .Y(n_145) );
INVx1_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx3_ASAP7_75t_L g140 ( .A(n_131), .Y(n_140) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_131), .Y(n_142) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
INVx1_ASAP7_75t_L g177 ( .A(n_131), .Y(n_177) );
INVx4_ASAP7_75t_SL g166 ( .A(n_132), .Y(n_166) );
BUFx3_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
INVx5_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx3_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_136), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_141), .B(n_143), .Y(n_138) );
INVx5_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_140), .B(n_487), .Y(n_486) );
INVx4_ASAP7_75t_L g254 ( .A(n_142), .Y(n_254) );
INVx2_ASAP7_75t_L g485 ( .A(n_142), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_143), .A2(n_176), .B(n_178), .Y(n_175) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx2_ASAP7_75t_L g522 ( .A(n_148), .Y(n_522) );
INVx5_ASAP7_75t_SL g240 ( .A(n_149), .Y(n_240) );
AND2x2_ASAP7_75t_L g259 ( .A(n_149), .B(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_149), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g345 ( .A(n_149), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g377 ( .A(n_149), .B(n_180), .Y(n_377) );
OR2x2_ASAP7_75t_L g383 ( .A(n_149), .B(n_273), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_149), .B(n_333), .Y(n_392) );
OR2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_168), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_153), .B(n_167), .Y(n_150) );
BUFx2_ASAP7_75t_L g210 ( .A(n_152), .Y(n_210) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_155), .A2(n_166), .B(n_184), .C(n_185), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_SL g248 ( .A1(n_155), .A2(n_166), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_155), .A2(n_166), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_155), .A2(n_166), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_155), .A2(n_166), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_155), .A2(n_166), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_SL g524 ( .A1(n_155), .A2(n_166), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_161), .C(n_163), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_158), .A2(n_163), .B(n_201), .C(n_202), .Y(n_200) );
O2A1O1Ixp5_ASAP7_75t_L g471 ( .A1(n_158), .A2(n_472), .B(n_473), .C(n_474), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_158), .A2(n_474), .B(n_548), .C(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx4_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_162), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g251 ( .A(n_162), .Y(n_251) );
OAI22xp33_ASAP7_75t_L g527 ( .A1(n_162), .A2(n_187), .B1(n_528), .B2(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_162), .A2(n_215), .B(n_537), .C(n_538), .Y(n_536) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g255 ( .A(n_164), .Y(n_255) );
INVx1_ASAP7_75t_L g497 ( .A(n_164), .Y(n_497) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_167), .A2(n_198), .B(n_199), .Y(n_197) );
INVx2_ASAP7_75t_L g217 ( .A(n_167), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_167), .A2(n_481), .B(n_488), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_180), .Y(n_169) );
AND2x2_ASAP7_75t_L g274 ( .A(n_170), .B(n_240), .Y(n_274) );
INVx1_ASAP7_75t_SL g287 ( .A(n_170), .Y(n_287) );
OR2x2_ASAP7_75t_L g322 ( .A(n_170), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g328 ( .A(n_170), .B(n_180), .Y(n_328) );
AND2x2_ASAP7_75t_L g386 ( .A(n_170), .B(n_237), .Y(n_386) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_171), .B(n_240), .Y(n_313) );
INVx3_ASAP7_75t_L g237 ( .A(n_180), .Y(n_237) );
OR2x2_ASAP7_75t_L g279 ( .A(n_180), .B(n_240), .Y(n_279) );
AND2x2_ASAP7_75t_L g289 ( .A(n_180), .B(n_287), .Y(n_289) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_180), .Y(n_337) );
AND2x2_ASAP7_75t_L g346 ( .A(n_180), .B(n_260), .Y(n_346) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_191), .Y(n_180) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_181), .A2(n_491), .B(n_498), .Y(n_490) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_181), .A2(n_500), .B(n_506), .Y(n_499) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_181), .A2(n_510), .B(n_517), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_186), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_187), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_187), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g215 ( .A(n_190), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_190), .B(n_527), .Y(n_526) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_192), .A2(n_247), .B(n_256), .Y(n_246) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_193), .A2(n_363), .B1(n_365), .B2(n_367), .C(n_370), .Y(n_362) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_205), .Y(n_194) );
AND2x2_ASAP7_75t_L g336 ( .A(n_195), .B(n_317), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_195), .B(n_395), .Y(n_399) );
OR2x2_ASAP7_75t_L g420 ( .A(n_195), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_195), .B(n_425), .Y(n_424) );
BUFx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx5_ASAP7_75t_L g267 ( .A(n_196), .Y(n_267) );
AND2x2_ASAP7_75t_L g344 ( .A(n_196), .B(n_207), .Y(n_344) );
AND2x2_ASAP7_75t_L g405 ( .A(n_196), .B(n_284), .Y(n_405) );
AND2x2_ASAP7_75t_L g418 ( .A(n_196), .B(n_237), .Y(n_418) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_203), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_221), .Y(n_205) );
AND2x4_ASAP7_75t_L g244 ( .A(n_206), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g263 ( .A(n_206), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g270 ( .A(n_206), .Y(n_270) );
AND2x2_ASAP7_75t_L g339 ( .A(n_206), .B(n_317), .Y(n_339) );
AND2x2_ASAP7_75t_L g349 ( .A(n_206), .B(n_267), .Y(n_349) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_206), .Y(n_357) );
AND2x2_ASAP7_75t_L g369 ( .A(n_206), .B(n_246), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_206), .B(n_301), .Y(n_373) );
AND2x2_ASAP7_75t_L g410 ( .A(n_206), .B(n_405), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_206), .B(n_284), .Y(n_421) );
OR2x2_ASAP7_75t_L g423 ( .A(n_206), .B(n_359), .Y(n_423) );
INVx5_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g309 ( .A(n_207), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g319 ( .A(n_207), .B(n_264), .Y(n_319) );
AND2x2_ASAP7_75t_L g331 ( .A(n_207), .B(n_246), .Y(n_331) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_207), .Y(n_361) );
AND2x4_ASAP7_75t_L g395 ( .A(n_207), .B(n_245), .Y(n_395) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_211), .B(n_216), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_217), .B(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_220), .A2(n_468), .B(n_475), .Y(n_467) );
BUFx2_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g284 ( .A(n_222), .Y(n_284) );
AND2x2_ASAP7_75t_L g317 ( .A(n_222), .B(n_246), .Y(n_317) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g264 ( .A(n_223), .B(n_246), .Y(n_264) );
BUFx2_ASAP7_75t_L g310 ( .A(n_223), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_231), .Y(n_224) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx3_ASAP7_75t_L g516 ( .A(n_230), .Y(n_516) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_236), .B(n_318), .Y(n_397) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_237), .B(n_260), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_237), .B(n_240), .Y(n_299) );
AND2x2_ASAP7_75t_L g354 ( .A(n_237), .B(n_290), .Y(n_354) );
AOI221xp5_ASAP7_75t_SL g291 ( .A1(n_238), .A2(n_292), .B1(n_300), .B2(n_302), .C(n_306), .Y(n_291) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g286 ( .A(n_239), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g327 ( .A(n_239), .B(n_328), .Y(n_327) );
OAI321xp33_ASAP7_75t_L g334 ( .A1(n_239), .A2(n_293), .A3(n_335), .B1(n_337), .B2(n_338), .C(n_340), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_240), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_243), .B(n_395), .Y(n_413) );
AND2x2_ASAP7_75t_L g300 ( .A(n_244), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_244), .B(n_304), .Y(n_303) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_245), .Y(n_276) );
AND2x2_ASAP7_75t_L g283 ( .A(n_245), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_245), .B(n_358), .Y(n_388) );
INVx1_ASAP7_75t_L g425 ( .A(n_245), .Y(n_425) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_254), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g474 ( .A(n_255), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B(n_262), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_259), .A2(n_369), .B(n_418), .C(n_419), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_260), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_260), .B(n_298), .Y(n_364) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g307 ( .A(n_264), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_264), .B(n_267), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_264), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_264), .B(n_349), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_268), .B1(n_280), .B2(n_285), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g281 ( .A(n_267), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g304 ( .A(n_267), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g316 ( .A(n_267), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_267), .B(n_310), .Y(n_352) );
OR2x2_ASAP7_75t_L g359 ( .A(n_267), .B(n_284), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_267), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g409 ( .A(n_267), .B(n_395), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .B1(n_275), .B2(n_277), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g315 ( .A(n_270), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
OAI22xp33_ASAP7_75t_L g355 ( .A1(n_273), .A2(n_288), .B1(n_356), .B2(n_360), .Y(n_355) );
INVx1_ASAP7_75t_L g403 ( .A(n_274), .Y(n_403) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_278), .A2(n_315), .B1(n_318), .B2(n_319), .C(n_320), .Y(n_314) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g293 ( .A(n_279), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_283), .B(n_349), .Y(n_381) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_284), .Y(n_301) );
INVx1_ASAP7_75t_L g305 ( .A(n_284), .Y(n_305) );
NAND2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g323 ( .A(n_290), .Y(n_323) );
AND2x2_ASAP7_75t_L g332 ( .A(n_290), .B(n_333), .Y(n_332) );
NAND2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g376 ( .A(n_297), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_300), .A2(n_326), .B1(n_329), .B2(n_332), .C(n_334), .Y(n_325) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_304), .B(n_361), .Y(n_360) );
AOI21xp33_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_308), .B(n_311), .Y(n_306) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_311), .Y(n_408) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
OR2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g371 ( .A(n_316), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_316), .B(n_376), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_319), .B(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND4xp25_ASAP7_75t_L g324 ( .A(n_325), .B(n_343), .C(n_362), .D(n_375), .Y(n_324) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g333 ( .A(n_328), .Y(n_333) );
INVxp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g366 ( .A(n_337), .B(n_342), .Y(n_366) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_345), .B(n_347), .C(n_355), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g414 ( .A1(n_345), .A2(n_387), .B(n_415), .C(n_422), .Y(n_414) );
INVx1_ASAP7_75t_SL g374 ( .A(n_346), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B1(n_352), .B2(n_353), .Y(n_347) );
INVx1_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_358), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_358), .B(n_369), .Y(n_402) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g379 ( .A(n_369), .Y(n_379) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B(n_374), .Y(n_370) );
INVxp33_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI322xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_378), .A3(n_379), .B1(n_380), .B2(n_382), .C1(n_384), .C2(n_387), .Y(n_375) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND3xp33_ASAP7_75t_SL g389 ( .A(n_390), .B(n_407), .C(n_414), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B1(n_396), .B2(n_398), .C(n_400), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g406 ( .A(n_395), .Y(n_406) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_403), .B2(n_404), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_410), .B2(n_411), .C(n_412), .Y(n_407) );
NAND2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g435 ( .A(n_427), .Y(n_435) );
BUFx2_ASAP7_75t_L g447 ( .A(n_427), .Y(n_447) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_428), .B(n_729), .Y(n_737) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g728 ( .A(n_429), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
NAND2xp33_ASAP7_75t_L g739 ( .A(n_434), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_441), .A2(n_442), .B(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_SL g740 ( .A(n_441), .B(n_443), .Y(n_740) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_450), .Y(n_730) );
INVx1_ASAP7_75t_L g454 ( .A(n_451), .Y(n_454) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g732 ( .A(n_458), .Y(n_732) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g733 ( .A(n_460), .Y(n_733) );
OR2x2_ASAP7_75t_SL g460 ( .A(n_461), .B(n_681), .Y(n_460) );
NAND5xp2_ASAP7_75t_L g461 ( .A(n_462), .B(n_593), .C(n_631), .D(n_652), .E(n_669), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_565), .C(n_586), .Y(n_462) );
OAI221xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_507), .B1(n_531), .B2(n_552), .C(n_556), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_477), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_466), .B(n_554), .Y(n_573) );
OR2x2_ASAP7_75t_L g600 ( .A(n_466), .B(n_490), .Y(n_600) );
AND2x2_ASAP7_75t_L g614 ( .A(n_466), .B(n_490), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_466), .B(n_480), .Y(n_628) );
AND2x2_ASAP7_75t_L g666 ( .A(n_466), .B(n_630), .Y(n_666) );
AND2x2_ASAP7_75t_L g695 ( .A(n_466), .B(n_605), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_466), .B(n_577), .Y(n_712) );
INVx4_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g592 ( .A(n_467), .B(n_489), .Y(n_592) );
BUFx3_ASAP7_75t_L g617 ( .A(n_467), .Y(n_617) );
AND2x2_ASAP7_75t_L g646 ( .A(n_467), .B(n_490), .Y(n_646) );
AND3x2_ASAP7_75t_L g659 ( .A(n_467), .B(n_660), .C(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g582 ( .A(n_477), .Y(n_582) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_489), .Y(n_477) );
AOI32xp33_ASAP7_75t_L g637 ( .A1(n_478), .A2(n_589), .A3(n_638), .B1(n_641), .B2(n_642), .Y(n_637) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g564 ( .A(n_479), .B(n_489), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_479), .B(n_592), .Y(n_635) );
AND2x2_ASAP7_75t_L g642 ( .A(n_479), .B(n_614), .Y(n_642) );
OR2x2_ASAP7_75t_L g648 ( .A(n_479), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_479), .B(n_603), .Y(n_673) );
OR2x2_ASAP7_75t_L g691 ( .A(n_479), .B(n_519), .Y(n_691) );
BUFx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g555 ( .A(n_480), .B(n_499), .Y(n_555) );
INVx2_ASAP7_75t_L g577 ( .A(n_480), .Y(n_577) );
OR2x2_ASAP7_75t_L g599 ( .A(n_480), .B(n_499), .Y(n_599) );
AND2x2_ASAP7_75t_L g604 ( .A(n_480), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_480), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g660 ( .A(n_480), .B(n_554), .Y(n_660) );
INVx1_ASAP7_75t_SL g711 ( .A(n_489), .Y(n_711) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
INVx1_ASAP7_75t_SL g554 ( .A(n_490), .Y(n_554) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_490), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_490), .B(n_640), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_490), .B(n_577), .C(n_695), .Y(n_706) );
INVx2_ASAP7_75t_L g605 ( .A(n_499), .Y(n_605) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_499), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
INVx1_ASAP7_75t_L g641 ( .A(n_508), .Y(n_641) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g559 ( .A(n_509), .B(n_542), .Y(n_559) );
INVx2_ASAP7_75t_L g576 ( .A(n_509), .Y(n_576) );
AND2x2_ASAP7_75t_L g581 ( .A(n_509), .B(n_543), .Y(n_581) );
AND2x2_ASAP7_75t_L g596 ( .A(n_509), .B(n_532), .Y(n_596) );
AND2x2_ASAP7_75t_L g608 ( .A(n_509), .B(n_580), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_518), .B(n_624), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g680 ( .A(n_518), .B(n_581), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_518), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_518), .B(n_575), .Y(n_703) );
BUFx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g541 ( .A(n_519), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_519), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g585 ( .A(n_519), .B(n_532), .Y(n_585) );
AND2x2_ASAP7_75t_L g611 ( .A(n_519), .B(n_542), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_519), .B(n_651), .Y(n_650) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_523), .B(n_530), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_521), .A2(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g570 ( .A(n_523), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_530), .Y(n_571) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_532), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g575 ( .A(n_532), .B(n_576), .Y(n_575) );
INVx3_ASAP7_75t_SL g580 ( .A(n_532), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_532), .B(n_567), .Y(n_633) );
OR2x2_ASAP7_75t_L g643 ( .A(n_532), .B(n_569), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_532), .B(n_611), .Y(n_671) );
OR2x2_ASAP7_75t_L g701 ( .A(n_532), .B(n_542), .Y(n_701) );
AND2x2_ASAP7_75t_L g705 ( .A(n_532), .B(n_543), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_532), .B(n_581), .Y(n_718) );
AND2x2_ASAP7_75t_L g725 ( .A(n_532), .B(n_607), .Y(n_725) );
OR2x6_ASAP7_75t_L g532 ( .A(n_533), .B(n_539), .Y(n_532) );
INVx1_ASAP7_75t_SL g668 ( .A(n_541), .Y(n_668) );
AND2x2_ASAP7_75t_L g607 ( .A(n_542), .B(n_569), .Y(n_607) );
AND2x2_ASAP7_75t_L g621 ( .A(n_542), .B(n_576), .Y(n_621) );
AND2x2_ASAP7_75t_L g624 ( .A(n_542), .B(n_580), .Y(n_624) );
INVx1_ASAP7_75t_L g651 ( .A(n_542), .Y(n_651) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g563 ( .A(n_543), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g722 ( .A1(n_553), .A2(n_599), .B(n_723), .C(n_724), .Y(n_722) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g629 ( .A(n_554), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_555), .B(n_572), .Y(n_587) );
AND2x2_ASAP7_75t_L g613 ( .A(n_555), .B(n_614), .Y(n_613) );
OAI21xp5_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_560), .B(n_564), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_558), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g584 ( .A(n_559), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_559), .B(n_580), .Y(n_625) );
AND2x2_ASAP7_75t_L g716 ( .A(n_559), .B(n_567), .Y(n_716) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g589 ( .A(n_563), .B(n_576), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_563), .B(n_574), .Y(n_590) );
OAI322xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_573), .A3(n_574), .B1(n_577), .B2(n_578), .C1(n_582), .C2(n_583), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_572), .Y(n_566) );
AND2x2_ASAP7_75t_L g677 ( .A(n_567), .B(n_589), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_567), .B(n_641), .Y(n_723) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g620 ( .A(n_569), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g686 ( .A(n_573), .B(n_599), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_574), .B(n_668), .Y(n_667) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_575), .B(n_607), .Y(n_664) );
AND2x2_ASAP7_75t_L g610 ( .A(n_576), .B(n_580), .Y(n_610) );
AND2x2_ASAP7_75t_L g618 ( .A(n_577), .B(n_619), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_577), .A2(n_656), .B(n_716), .C(n_717), .Y(n_715) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_578), .A2(n_591), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_580), .B(n_607), .Y(n_647) );
AND2x2_ASAP7_75t_L g653 ( .A(n_580), .B(n_621), .Y(n_653) );
AND2x2_ASAP7_75t_L g687 ( .A(n_580), .B(n_589), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_581), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_SL g697 ( .A(n_581), .Y(n_697) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_585), .A2(n_613), .B1(n_615), .B2(n_620), .Y(n_612) );
OAI22xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_588), .B1(n_590), .B2(n_591), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_587), .A2(n_623), .B1(n_625), .B2(n_626), .Y(n_622) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_592), .A2(n_694), .B1(n_696), .B2(n_698), .C(n_702), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B(n_601), .C(n_622), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
OR2x2_ASAP7_75t_L g663 ( .A(n_599), .B(n_616), .Y(n_663) );
INVx1_ASAP7_75t_L g714 ( .A(n_599), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_600), .A2(n_602), .B1(n_606), .B2(n_609), .C(n_612), .Y(n_601) );
INVx2_ASAP7_75t_SL g656 ( .A(n_600), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g721 ( .A(n_603), .Y(n_721) );
AND2x2_ASAP7_75t_L g645 ( .A(n_604), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g630 ( .A(n_605), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g692 ( .A(n_608), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_616), .B(n_718), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g616 ( .A(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_L g661 ( .A(n_619), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_620), .A2(n_632), .B(n_634), .C(n_636), .Y(n_631) );
INVx1_ASAP7_75t_L g709 ( .A(n_623), .Y(n_709) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_627), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx2_ASAP7_75t_L g640 ( .A(n_630), .Y(n_640) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI222xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_643), .B1(n_644), .B2(n_647), .C1(n_648), .C2(n_650), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g676 ( .A(n_640), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_643), .B(n_697), .Y(n_696) );
NAND2xp33_ASAP7_75t_SL g674 ( .A(n_644), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g649 ( .A(n_646), .Y(n_649) );
AND2x2_ASAP7_75t_L g713 ( .A(n_646), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g679 ( .A(n_649), .B(n_676), .Y(n_679) );
INVx1_ASAP7_75t_L g708 ( .A(n_650), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_657), .C(n_662), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_656), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
AOI322xp5_ASAP7_75t_L g707 ( .A1(n_659), .A2(n_687), .A3(n_692), .B1(n_708), .B2(n_709), .C1(n_710), .C2(n_713), .Y(n_707) );
AND2x2_ASAP7_75t_L g694 ( .A(n_660), .B(n_695), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_665), .B2(n_667), .Y(n_662) );
INVxp33_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B1(n_674), .B2(n_677), .C(n_678), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
NAND5xp2_ASAP7_75t_L g681 ( .A(n_682), .B(n_693), .C(n_707), .D(n_715), .E(n_719), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B(n_688), .Y(n_682) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVxp33_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_695), .A2(n_720), .B(n_721), .C(n_722), .Y(n_719) );
AOI31xp33_ASAP7_75t_L g702 ( .A1(n_697), .A2(n_703), .A3(n_704), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g734 ( .A(n_727), .Y(n_734) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
endmodule