module fake_jpeg_7353_n_107 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_107);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_30),
.B1(n_21),
.B2(n_13),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_17),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_12),
.B(n_20),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_32),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_15),
.B1(n_18),
.B2(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_24),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_29),
.B(n_30),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_54),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_53),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_29),
.B1(n_32),
.B2(n_28),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_58),
.C(n_54),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_16),
.C(n_12),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_12),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_25),
.B1(n_27),
.B2(n_21),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_68),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_65),
.B(n_51),
.C(n_49),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_27),
.B(n_19),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_69),
.C(n_52),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_16),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_56),
.B1(n_50),
.B2(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_78),
.B1(n_74),
.B2(n_69),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_59),
.C(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_77),
.Y(n_82)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

XOR2x2_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_44),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_78),
.B(n_58),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_65),
.B1(n_61),
.B2(n_60),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_48),
.C(n_55),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_22),
.C(n_25),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_85),
.C(n_86),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_47),
.C(n_75),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_25),
.C(n_18),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.C(n_72),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_79),
.B(n_76),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_20),
.B(n_5),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_79),
.B1(n_92),
.B2(n_20),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.C(n_9),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_79),
.C(n_16),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_6),
.C(n_8),
.Y(n_101)
);

OAI321xp33_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_8),
.C(n_4),
.Y(n_98)
);

AOI31xp67_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_11),
.A3(n_7),
.B(n_8),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_102),
.B(n_101),
.CI(n_99),
.CON(n_105),
.SN(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_104),
.C(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);


endmodule