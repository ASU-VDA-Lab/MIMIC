module fake_aes_4598_n_542 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_542);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_542;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_165;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_51), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_46), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_35), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_63), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_52), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_12), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_15), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_32), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_21), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_58), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_77), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_18), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_8), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_66), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_42), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_57), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_62), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_34), .Y(n_96) );
INVxp33_ASAP7_75t_SL g97 ( .A(n_13), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_43), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_14), .Y(n_99) );
BUFx2_ASAP7_75t_L g100 ( .A(n_0), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_13), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_10), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_74), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_45), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_64), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_23), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_38), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_76), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_24), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_27), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_5), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_9), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_78), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_0), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_100), .B(n_84), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_106), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_106), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_87), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_106), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_106), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_106), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_106), .Y(n_124) );
NOR2xp33_ASAP7_75t_SL g125 ( .A(n_86), .B(n_31), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_79), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_105), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_105), .B(n_1), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_83), .B(n_1), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_83), .B(n_2), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_89), .B(n_2), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_114), .B(n_109), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_134), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_123), .Y(n_141) );
NOR3xp33_ASAP7_75t_L g142 ( .A(n_115), .B(n_112), .C(n_89), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
BUFx3_ASAP7_75t_L g144 ( .A(n_132), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g146 ( .A1(n_119), .A2(n_112), .B1(n_90), .B2(n_101), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
INVx1_ASAP7_75t_SL g148 ( .A(n_134), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
INVx2_ASAP7_75t_SL g151 ( .A(n_114), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_134), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_123), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_135), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_121), .B(n_103), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_135), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_121), .B(n_126), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_123), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_142), .B(n_135), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_143), .B(n_131), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
AO22x1_ASAP7_75t_L g166 ( .A1(n_160), .A2(n_85), .B1(n_96), .B2(n_104), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_151), .B(n_126), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_147), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_142), .B(n_131), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_160), .B(n_94), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_151), .B(n_133), .Y(n_176) );
AO22x1_ASAP7_75t_L g177 ( .A1(n_148), .A2(n_108), .B1(n_130), .B2(n_129), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_140), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_140), .Y(n_179) );
CKINVDCx6p67_ASAP7_75t_R g180 ( .A(n_143), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_140), .B(n_129), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_148), .B(n_81), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
INVx5_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_157), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_139), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
INVxp67_ASAP7_75t_SL g192 ( .A(n_151), .Y(n_192) );
INVx5_ASAP7_75t_L g193 ( .A(n_159), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_139), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_139), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_159), .A2(n_139), .B1(n_152), .B2(n_137), .Y(n_196) );
INVx1_ASAP7_75t_SL g197 ( .A(n_180), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_186), .B(n_159), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_186), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_173), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_163), .A2(n_159), .B1(n_139), .B2(n_152), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_180), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_186), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_180), .A2(n_152), .B1(n_137), .B2(n_161), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_173), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_189), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_186), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_164), .B(n_161), .Y(n_208) );
BUFx8_ASAP7_75t_SL g209 ( .A(n_174), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_186), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_189), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_186), .B(n_152), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_194), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_186), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_194), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_193), .B(n_152), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_193), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_193), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_193), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_164), .B(n_146), .Y(n_220) );
INVxp67_ASAP7_75t_SL g221 ( .A(n_191), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_193), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_163), .A2(n_158), .B1(n_130), .B2(n_133), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_195), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_169), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_174), .A2(n_146), .B1(n_158), .B2(n_97), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_181), .A2(n_156), .B(n_154), .C(n_128), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_193), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_187), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_225), .B(n_174), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_225), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_206), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_206), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_199), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_229), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_199), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_211), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_211), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_199), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_227), .A2(n_192), .B(n_168), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_213), .A2(n_176), .B(n_168), .C(n_172), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_204), .A2(n_163), .B(n_175), .C(n_174), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_213), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_201), .A2(n_195), .B(n_171), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_215), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_223), .A2(n_163), .B1(n_184), .B2(n_177), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_220), .A2(n_184), .B1(n_191), .B2(n_182), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_208), .A2(n_166), .B1(n_90), .B2(n_101), .C(n_102), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_220), .B(n_200), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_224), .Y(n_251) );
BUFx12f_ASAP7_75t_L g252 ( .A(n_202), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_203), .B(n_217), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_224), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_226), .A2(n_184), .B1(n_177), .B2(n_176), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_198), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_232), .Y(n_257) );
AOI22xp33_ASAP7_75t_SL g258 ( .A1(n_235), .A2(n_197), .B1(n_205), .B2(n_184), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_246), .A2(n_184), .B1(n_201), .B2(n_221), .Y(n_259) );
AOI211xp5_ASAP7_75t_L g260 ( .A1(n_249), .A2(n_166), .B(n_102), .C(n_113), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_250), .A2(n_209), .B1(n_184), .B2(n_216), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_232), .Y(n_262) );
NAND3xp33_ASAP7_75t_L g263 ( .A(n_249), .B(n_125), .C(n_132), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_230), .B(n_219), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_231), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_250), .B(n_232), .Y(n_266) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_240), .A2(n_120), .B(n_117), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_245), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_246), .A2(n_184), .B1(n_212), .B2(n_216), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_255), .A2(n_184), .B1(n_212), .B2(n_216), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_255), .A2(n_216), .B1(n_212), .B2(n_219), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_230), .A2(n_212), .B1(n_203), .B2(n_217), .Y(n_272) );
AO31x2_ASAP7_75t_L g273 ( .A1(n_245), .A2(n_127), .A3(n_117), .B(n_118), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_245), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_248), .A2(n_198), .B1(n_196), .B2(n_214), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_253), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_231), .A2(n_222), .B1(n_214), .B2(n_217), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_257), .B(n_231), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_260), .B(n_132), .C(n_82), .Y(n_280) );
AOI31xp33_ASAP7_75t_L g281 ( .A1(n_258), .A2(n_252), .A3(n_253), .B(n_99), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_261), .A2(n_252), .B1(n_254), .B2(n_238), .Y(n_282) );
AND2x4_ASAP7_75t_L g283 ( .A(n_257), .B(n_233), .Y(n_283) );
INVxp67_ASAP7_75t_L g284 ( .A(n_266), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_262), .Y(n_285) );
NAND3xp33_ASAP7_75t_SL g286 ( .A(n_259), .B(n_242), .C(n_110), .Y(n_286) );
OAI221xp5_ASAP7_75t_SL g287 ( .A1(n_259), .A2(n_256), .B1(n_107), .B2(n_110), .C(n_88), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g288 ( .A1(n_269), .A2(n_244), .B1(n_256), .B2(n_251), .C(n_247), .Y(n_288) );
AOI33xp33_ASAP7_75t_L g289 ( .A1(n_270), .A2(n_98), .A3(n_82), .B1(n_88), .B2(n_111), .B3(n_107), .Y(n_289) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_262), .A2(n_244), .B(n_251), .Y(n_290) );
AND2x4_ASAP7_75t_SL g291 ( .A(n_277), .B(n_253), .Y(n_291) );
AOI22xp33_ASAP7_75t_SL g292 ( .A1(n_263), .A2(n_252), .B1(n_253), .B2(n_254), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g293 ( .A1(n_266), .A2(n_247), .B1(n_243), .B2(n_233), .Y(n_293) );
NAND4xp25_ASAP7_75t_L g294 ( .A(n_271), .B(n_92), .C(n_93), .D(n_95), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_264), .A2(n_243), .B1(n_238), .B2(n_237), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_272), .A2(n_237), .B1(n_234), .B2(n_239), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_268), .Y(n_297) );
OAI211xp5_ASAP7_75t_L g298 ( .A1(n_276), .A2(n_98), .B(n_92), .C(n_93), .Y(n_298) );
OAI221xp5_ASAP7_75t_L g299 ( .A1(n_268), .A2(n_241), .B1(n_222), .B2(n_203), .C(n_228), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_274), .B(n_236), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_279), .Y(n_301) );
AND2x2_ASAP7_75t_SL g302 ( .A(n_289), .B(n_274), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_297), .B(n_265), .Y(n_303) );
AOI221xp5_ASAP7_75t_SL g304 ( .A1(n_281), .A2(n_95), .B1(n_111), .B2(n_264), .C(n_154), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_284), .B(n_265), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_297), .B(n_275), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_285), .Y(n_308) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_294), .B(n_132), .C(n_91), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_290), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_290), .Y(n_311) );
AOI33xp33_ASAP7_75t_L g312 ( .A1(n_295), .A2(n_156), .A3(n_118), .B1(n_120), .B2(n_122), .B3(n_124), .Y(n_312) );
OAI21xp33_ASAP7_75t_L g313 ( .A1(n_289), .A2(n_117), .B(n_124), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_283), .B(n_275), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_293), .A2(n_132), .B1(n_278), .B2(n_118), .C(n_120), .Y(n_315) );
AOI33xp33_ASAP7_75t_L g316 ( .A1(n_282), .A2(n_122), .A3(n_124), .B1(n_5), .B2(n_6), .B3(n_7), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_286), .A2(n_275), .B1(n_234), .B2(n_239), .Y(n_317) );
NOR2x1p5_ASAP7_75t_L g318 ( .A(n_283), .B(n_236), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_283), .B(n_273), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_300), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_300), .B(n_273), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_291), .B(n_273), .Y(n_324) );
AOI33xp33_ASAP7_75t_L g325 ( .A1(n_292), .A2(n_122), .A3(n_4), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_325) );
AOI21xp5_ASAP7_75t_SL g326 ( .A1(n_288), .A2(n_267), .B(n_198), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_287), .A2(n_123), .B1(n_172), .B2(n_183), .C(n_167), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_291), .B(n_273), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_298), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_322), .B(n_273), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_322), .B(n_267), .Y(n_332) );
OAI21xp33_ASAP7_75t_L g333 ( .A1(n_325), .A2(n_280), .B(n_123), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_321), .B(n_267), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_308), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_308), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_301), .B(n_267), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g339 ( .A(n_304), .B(n_239), .C(n_236), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g340 ( .A(n_316), .B(n_239), .C(n_236), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_321), .B(n_3), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_307), .B(n_22), .Y(n_342) );
NAND4xp25_ASAP7_75t_L g343 ( .A(n_330), .B(n_144), .C(n_145), .D(n_9), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_307), .B(n_3), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_320), .B(n_4), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_305), .B(n_10), .Y(n_348) );
OAI33xp33_ASAP7_75t_L g349 ( .A1(n_330), .A2(n_11), .A3(n_12), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_310), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_323), .B(n_11), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_323), .B(n_16), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_328), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_306), .B(n_17), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_319), .B(n_17), .Y(n_357) );
OAI33xp33_ASAP7_75t_L g358 ( .A1(n_319), .A2(n_18), .A3(n_19), .B1(n_20), .B2(n_150), .B3(n_155), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_314), .B(n_19), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_314), .B(n_20), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_324), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_302), .B(n_183), .Y(n_362) );
AO211x2_ASAP7_75t_L g363 ( .A1(n_309), .A2(n_25), .B(n_26), .C(n_28), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_324), .B(n_145), .Y(n_364) );
NAND4xp25_ASAP7_75t_L g365 ( .A(n_326), .B(n_144), .C(n_145), .D(n_198), .Y(n_365) );
OAI21xp33_ASAP7_75t_L g366 ( .A1(n_326), .A2(n_145), .B(n_150), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_318), .Y(n_367) );
NOR3xp33_ASAP7_75t_L g368 ( .A(n_329), .B(n_228), .C(n_218), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_302), .B(n_188), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_318), .B(n_29), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_329), .B(n_210), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_302), .Y(n_372) );
INVx2_ASAP7_75t_SL g373 ( .A(n_329), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_313), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_317), .B(n_30), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_335), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_355), .B(n_33), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_351), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
XNOR2xp5_ASAP7_75t_L g380 ( .A(n_359), .B(n_327), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
AND3x1_ASAP7_75t_L g382 ( .A(n_373), .B(n_312), .C(n_315), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_347), .B(n_37), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_372), .B(n_150), .C(n_155), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_359), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_361), .B(n_39), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_336), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_361), .B(n_40), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_347), .B(n_41), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_336), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_352), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_351), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_360), .B(n_44), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_352), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_331), .B(n_47), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_331), .B(n_48), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_332), .B(n_49), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_338), .B(n_50), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_346), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_343), .A2(n_373), .B1(n_368), .B2(n_349), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g402 ( .A1(n_366), .A2(n_162), .B(n_155), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_350), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_332), .B(n_53), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_350), .B(n_54), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_334), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_334), .B(n_55), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_353), .B(n_56), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_337), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_357), .B(n_199), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_357), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_353), .B(n_354), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_364), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_364), .B(n_59), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g415 ( .A1(n_365), .A2(n_228), .B(n_218), .C(n_210), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_345), .B(n_60), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_354), .B(n_61), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g418 ( .A1(n_339), .A2(n_228), .B(n_218), .C(n_210), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_356), .B(n_65), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_341), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_356), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_345), .B(n_67), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_341), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_348), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_348), .B(n_367), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_362), .B(n_68), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_369), .B(n_70), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_406), .B(n_342), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_391), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_406), .B(n_342), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_394), .Y(n_431) );
NOR2xp33_ASAP7_75t_SL g432 ( .A(n_385), .B(n_370), .Y(n_432) );
OAI32xp33_ASAP7_75t_L g433 ( .A1(n_385), .A2(n_371), .A3(n_370), .B1(n_374), .B2(n_375), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_421), .A2(n_358), .B1(n_333), .B2(n_340), .C(n_342), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_403), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_399), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_413), .B(n_371), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_376), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_413), .B(n_374), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_379), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_418), .A2(n_363), .B(n_375), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_425), .B(n_71), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_387), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_401), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_SL g446 ( .A1(n_418), .A2(n_363), .B(n_218), .C(n_75), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_390), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_422), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_424), .B(n_72), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_381), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_381), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_411), .B(n_73), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_420), .B(n_150), .Y(n_453) );
INVx2_ASAP7_75t_SL g454 ( .A(n_378), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_378), .B(n_155), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_420), .B(n_162), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_409), .B(n_162), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_416), .A2(n_210), .B1(n_207), .B2(n_199), .Y(n_459) );
NAND2xp33_ASAP7_75t_L g460 ( .A(n_422), .B(n_210), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_392), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_423), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_423), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_412), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_410), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_395), .B(n_162), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_392), .B(n_141), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_410), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_395), .B(n_141), .Y(n_469) );
AOI21xp33_ASAP7_75t_L g470 ( .A1(n_400), .A2(n_141), .B(n_207), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_380), .B(n_207), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_382), .A2(n_207), .B1(n_188), .B2(n_167), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_396), .B(n_207), .Y(n_473) );
O2A1O1Ixp5_ASAP7_75t_L g474 ( .A1(n_415), .A2(n_169), .B(n_170), .C(n_171), .Y(n_474) );
XNOR2xp5_ASAP7_75t_L g475 ( .A(n_416), .B(n_185), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_377), .Y(n_476) );
AOI211xp5_ASAP7_75t_L g477 ( .A1(n_396), .A2(n_141), .B(n_185), .C(n_169), .Y(n_477) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_419), .A2(n_141), .B(n_170), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_377), .Y(n_479) );
XNOR2xp5_ASAP7_75t_L g480 ( .A(n_414), .B(n_170), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_405), .Y(n_481) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_386), .B(n_182), .Y(n_482) );
OAI31xp33_ASAP7_75t_L g483 ( .A1(n_419), .A2(n_182), .A3(n_178), .B(n_179), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_405), .Y(n_484) );
XNOR2x1_ASAP7_75t_L g485 ( .A(n_414), .B(n_182), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g486 ( .A1(n_393), .A2(n_141), .B1(n_190), .B2(n_165), .C(n_178), .Y(n_486) );
NOR2x1_ASAP7_75t_L g487 ( .A(n_386), .B(n_141), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_386), .A2(n_193), .B(n_178), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_407), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_397), .A2(n_179), .B(n_141), .C(n_190), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_383), .A2(n_165), .B(n_190), .C(n_389), .Y(n_491) );
NAND2xp33_ASAP7_75t_L g492 ( .A(n_397), .B(n_165), .Y(n_492) );
AOI21xp33_ASAP7_75t_SL g493 ( .A1(n_388), .A2(n_165), .B(n_404), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_404), .A2(n_165), .B1(n_407), .B2(n_384), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_426), .B(n_165), .C(n_427), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g496 ( .A1(n_407), .A2(n_408), .B(n_417), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_398), .B(n_402), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_391), .Y(n_498) );
OAI21xp33_ASAP7_75t_L g499 ( .A1(n_400), .A2(n_425), .B(n_421), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_385), .A2(n_373), .B1(n_380), .B2(n_400), .Y(n_500) );
OAI321xp33_ASAP7_75t_L g501 ( .A1(n_500), .A2(n_499), .A3(n_434), .B1(n_471), .B2(n_494), .C(n_442), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_429), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_482), .A2(n_475), .B1(n_496), .B2(n_448), .Y(n_503) );
XNOR2x1_ASAP7_75t_L g504 ( .A(n_464), .B(n_480), .Y(n_504) );
AOI21x1_ASAP7_75t_L g505 ( .A1(n_487), .A2(n_494), .B(n_445), .Y(n_505) );
OAI21xp33_ASAP7_75t_L g506 ( .A1(n_432), .A2(n_470), .B(n_433), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_498), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g508 ( .A(n_472), .B(n_477), .C(n_474), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g509 ( .A1(n_443), .A2(n_491), .B(n_433), .Y(n_509) );
OAI21xp5_ASAP7_75t_SL g510 ( .A1(n_459), .A2(n_493), .B(n_488), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_454), .A2(n_461), .B1(n_489), .B2(n_488), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_436), .A2(n_435), .B1(n_479), .B2(n_476), .C(n_431), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_437), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_447), .Y(n_514) );
NOR2x1p5_ASAP7_75t_L g515 ( .A(n_435), .B(n_465), .Y(n_515) );
OAI211xp5_ASAP7_75t_SL g516 ( .A1(n_483), .A2(n_460), .B(n_446), .C(n_492), .Y(n_516) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_460), .B(n_495), .Y(n_517) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_454), .A2(n_437), .B1(n_468), .B2(n_473), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_512), .B(n_503), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g520 ( .A1(n_506), .A2(n_446), .B1(n_463), .B2(n_462), .C(n_490), .Y(n_520) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_508), .Y(n_521) );
AOI21xp33_ASAP7_75t_L g522 ( .A1(n_501), .A2(n_449), .B(n_452), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_509), .A2(n_478), .B(n_497), .C(n_486), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_502), .Y(n_524) );
AOI221x1_ASAP7_75t_L g525 ( .A1(n_511), .A2(n_455), .B1(n_466), .B2(n_457), .C(n_453), .Y(n_525) );
AO22x2_ASAP7_75t_L g526 ( .A1(n_504), .A2(n_444), .B1(n_439), .B2(n_441), .Y(n_526) );
XNOR2x1_ASAP7_75t_L g527 ( .A(n_515), .B(n_485), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_507), .Y(n_528) );
OAI211xp5_ASAP7_75t_L g529 ( .A1(n_521), .A2(n_510), .B(n_508), .C(n_516), .Y(n_529) );
OAI22x1_ASAP7_75t_L g530 ( .A1(n_519), .A2(n_505), .B1(n_517), .B2(n_514), .Y(n_530) );
NAND4xp25_ASAP7_75t_L g531 ( .A(n_520), .B(n_469), .C(n_467), .D(n_428), .Y(n_531) );
NAND3xp33_ASAP7_75t_SL g532 ( .A(n_523), .B(n_469), .C(n_513), .Y(n_532) );
AOI221x1_ASAP7_75t_L g533 ( .A1(n_526), .A2(n_455), .B1(n_458), .B2(n_450), .C(n_451), .Y(n_533) );
OAI222xp33_ASAP7_75t_L g534 ( .A1(n_529), .A2(n_526), .B1(n_528), .B2(n_524), .C1(n_518), .C2(n_527), .Y(n_534) );
AND3x1_ASAP7_75t_L g535 ( .A(n_530), .B(n_522), .C(n_525), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_531), .A2(n_456), .B1(n_484), .B2(n_481), .Y(n_536) );
AOI322xp5_ASAP7_75t_L g537 ( .A1(n_534), .A2(n_532), .A3(n_533), .B1(n_440), .B2(n_438), .C1(n_428), .C2(n_430), .Y(n_537) );
XNOR2xp5_ASAP7_75t_L g538 ( .A(n_535), .B(n_440), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_538), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_539), .Y(n_540) );
XNOR2xp5_ASAP7_75t_L g541 ( .A(n_540), .B(n_536), .Y(n_541) );
AOI21xp33_ASAP7_75t_SL g542 ( .A1(n_541), .A2(n_537), .B(n_467), .Y(n_542) );
endmodule