module fake_jpeg_32012_n_165 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_73),
.B(n_49),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_80),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_64),
.B1(n_62),
.B2(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_85),
.B1(n_60),
.B2(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_50),
.B1(n_57),
.B2(n_47),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_54),
.B1(n_45),
.B2(n_57),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_97),
.B1(n_105),
.B2(n_4),
.Y(n_125)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_99),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_0),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_56),
.B1(n_51),
.B2(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_44),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_1),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_83),
.B(n_84),
.C(n_24),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_79),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_114),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_21),
.A3(n_43),
.B1(n_39),
.B2(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_116),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_125),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_96),
.C(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_11),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_2),
.C(n_3),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_123),
.C(n_7),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_95),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_3),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_4),
.B(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_20),
.B1(n_36),
.B2(n_35),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_121),
.B1(n_117),
.B2(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_13),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_140),
.B1(n_125),
.B2(n_17),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_133),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_7),
.B(n_9),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_136),
.B(n_14),
.Y(n_145)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_137),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_9),
.B(n_10),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_141),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_143),
.B(n_144),
.Y(n_148)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_16),
.C(n_19),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_150),
.C(n_140),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_26),
.C(n_28),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_155),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_142),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_148),
.C(n_151),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_158),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_149),
.C(n_128),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_153),
.C(n_127),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_131),
.B(n_135),
.Y(n_164)
);

OAI222xp33_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_135),
.B1(n_132),
.B2(n_30),
.C1(n_31),
.C2(n_32),
.Y(n_165)
);


endmodule