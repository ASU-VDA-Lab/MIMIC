module real_jpeg_25936_n_15 (n_108, n_8, n_0, n_111, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_106, n_11, n_14, n_110, n_7, n_3, n_5, n_4, n_102, n_105, n_109, n_101, n_1, n_13, n_103, n_15);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_106;
input n_11;
input n_14;
input n_110;
input n_7;
input n_3;
input n_5;
input n_4;
input n_102;
input n_105;
input n_109;
input n_101;
input n_1;
input n_13;
input n_103;

output n_15;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

BUFx10_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_2),
.B(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_3),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_5),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_5),
.B(n_56),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_6),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_8),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_8),
.B(n_74),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_9),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_9),
.B(n_90),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_11),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_13),
.B(n_36),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_29),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_28),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_24),
.B(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_26),
.B(n_97),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_27),
.B(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_27),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_94),
.B(n_99),
.Y(n_29)
);

OAI321xp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_84),
.A3(n_89),
.B1(n_92),
.B2(n_93),
.C(n_101),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_78),
.B(n_83),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_73),
.B(n_77),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_67),
.B(n_72),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B(n_66),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_59),
.B(n_65),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_55),
.B(n_58),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_49),
.B(n_54),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_79),
.B(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_98),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_102),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_103),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_104),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_105),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_106),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_107),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_108),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_109),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_110),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_111),
.Y(n_91)
);


endmodule