module fake_aes_7428_n_1405 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1405);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1405;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_1399;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_315;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1117;
wire n_1007;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1390;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g300 ( .A(n_247), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_250), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_79), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_115), .Y(n_303) );
INVxp33_ASAP7_75t_L g304 ( .A(n_133), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_75), .Y(n_305) );
INVxp33_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_173), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_176), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_242), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_83), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_11), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_169), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_76), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_77), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_24), .Y(n_315) );
NOR2xp67_ASAP7_75t_L g316 ( .A(n_51), .B(n_145), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_270), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_106), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_251), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_201), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_213), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_151), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_153), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_197), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_191), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_227), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_100), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_56), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_134), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_229), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_184), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_182), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_245), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_0), .Y(n_334) );
CKINVDCx14_ASAP7_75t_R g335 ( .A(n_266), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_243), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_240), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_78), .Y(n_338) );
INVxp33_ASAP7_75t_L g339 ( .A(n_136), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_67), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_224), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_158), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_84), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_122), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_126), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_157), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_53), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_190), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_155), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_154), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_15), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_253), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_293), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_238), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_119), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_12), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_63), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_172), .Y(n_358) );
CKINVDCx14_ASAP7_75t_R g359 ( .A(n_179), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_108), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_276), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_63), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_279), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_164), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_52), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_187), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_33), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_149), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_249), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_47), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_25), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_283), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_272), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_220), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_159), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_207), .Y(n_376) );
INVxp33_ASAP7_75t_SL g377 ( .A(n_105), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_257), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_81), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_160), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_121), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_79), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_194), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_156), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_222), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_271), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_264), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_236), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_167), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_297), .Y(n_390) );
INVxp33_ASAP7_75t_L g391 ( .A(n_123), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_58), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_55), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_108), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_268), .Y(n_395) );
INVxp67_ASAP7_75t_L g396 ( .A(n_43), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_84), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_41), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_287), .Y(n_399) );
BUFx5_ASAP7_75t_L g400 ( .A(n_234), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_178), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_202), .Y(n_402) );
INVxp33_ASAP7_75t_L g403 ( .A(n_274), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_53), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_22), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_130), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_2), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_168), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_24), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_260), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_77), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_7), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_41), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_54), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_128), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_44), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_228), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_36), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_16), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_241), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_12), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_129), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_137), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_237), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_165), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_69), .B(n_120), .Y(n_426) );
CKINVDCx14_ASAP7_75t_R g427 ( .A(n_132), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_186), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_58), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_290), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_269), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_138), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_42), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_56), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_212), .Y(n_435) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_13), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_215), .B(n_57), .Y(n_437) );
INVxp33_ASAP7_75t_SL g438 ( .A(n_278), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_235), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_69), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_289), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_265), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_32), .Y(n_443) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_117), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_127), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_38), .Y(n_446) );
INVxp33_ASAP7_75t_L g447 ( .A(n_226), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_91), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_67), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_11), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_175), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_221), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_3), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_21), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_163), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_211), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_440), .B(n_0), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_440), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_440), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_425), .B(n_1), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_300), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_375), .Y(n_462) );
NAND2xp33_ASAP7_75t_SL g463 ( .A(n_305), .B(n_1), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_300), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_301), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_301), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_323), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_323), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_425), .B(n_2), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_322), .Y(n_470) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_314), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_322), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_324), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_305), .B(n_4), .Y(n_474) );
INVxp33_ASAP7_75t_SL g475 ( .A(n_386), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_323), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_324), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_326), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_392), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_326), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_323), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_331), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_323), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_417), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_417), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_331), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_417), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_332), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_417), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_351), .B(n_5), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_332), .Y(n_491) );
OAI21x1_ASAP7_75t_L g492 ( .A1(n_352), .A2(n_114), .B(n_113), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_417), .Y(n_493) );
BUFx3_ASAP7_75t_L g494 ( .A(n_457), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_457), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_457), .Y(n_496) );
NAND3x1_ASAP7_75t_L g497 ( .A(n_474), .B(n_337), .C(n_333), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_467), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_460), .B(n_351), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_457), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_479), .B(n_335), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_460), .B(n_392), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_466), .A2(n_334), .B1(n_347), .B2(n_328), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_457), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_479), .B(n_359), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_457), .B(n_352), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_458), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_458), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
NOR2xp33_ASAP7_75t_SL g510 ( .A(n_466), .B(n_307), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_467), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_458), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_459), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_459), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_492), .Y(n_516) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_467), .Y(n_517) );
INVxp67_ASAP7_75t_L g518 ( .A(n_479), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_464), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_460), .B(n_427), .Y(n_520) );
INVx4_ASAP7_75t_L g521 ( .A(n_460), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_459), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_467), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_474), .A2(n_362), .B1(n_314), .B2(n_377), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_475), .B(n_304), .Y(n_525) );
AND2x6_ASAP7_75t_L g526 ( .A(n_460), .B(n_333), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_464), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_464), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_466), .A2(n_334), .B1(n_347), .B2(n_328), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_464), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_460), .B(n_442), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_470), .B(n_344), .C(n_337), .Y(n_532) );
OR2x2_ASAP7_75t_SL g533 ( .A(n_469), .B(n_356), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_470), .B(n_397), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_464), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_467), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_465), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_470), .B(n_346), .C(n_344), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_467), .Y(n_540) );
OR2x6_ASAP7_75t_L g541 ( .A(n_471), .B(n_406), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_472), .B(n_455), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_465), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_519), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_516), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_519), .Y(n_546) );
NOR2xp33_ASAP7_75t_R g547 ( .A(n_510), .B(n_462), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_539), .B(n_475), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_519), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_519), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_521), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_508), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_519), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_539), .B(n_461), .Y(n_554) );
BUFx3_ASAP7_75t_L g555 ( .A(n_526), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_539), .B(n_472), .Y(n_556) );
AO22x1_ASAP7_75t_L g557 ( .A1(n_526), .A2(n_438), .B1(n_377), .B2(n_383), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_510), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_525), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_526), .A2(n_463), .B1(n_473), .B2(n_472), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_525), .Y(n_561) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_494), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_501), .Y(n_563) );
BUFx3_ASAP7_75t_L g564 ( .A(n_526), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_501), .B(n_490), .Y(n_565) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_521), .B(n_465), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_530), .Y(n_567) );
INVx3_ASAP7_75t_L g568 ( .A(n_521), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_530), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_530), .Y(n_570) );
INVx3_ASAP7_75t_L g571 ( .A(n_521), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_508), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_518), .B(n_463), .C(n_490), .Y(n_573) );
BUFx3_ASAP7_75t_L g574 ( .A(n_526), .Y(n_574) );
OR2x6_ASAP7_75t_L g575 ( .A(n_521), .B(n_471), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_508), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_533), .A2(n_307), .B1(n_341), .B2(n_325), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_526), .A2(n_477), .B1(n_478), .B2(n_473), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_508), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_508), .Y(n_580) );
OR2x6_ASAP7_75t_L g581 ( .A(n_501), .B(n_492), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_530), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_518), .B(n_461), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_513), .Y(n_584) );
BUFx12f_ASAP7_75t_L g585 ( .A(n_533), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_513), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_513), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_513), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_516), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_513), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_542), .B(n_480), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_494), .Y(n_592) );
BUFx3_ASAP7_75t_L g593 ( .A(n_526), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_515), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_515), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_515), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_542), .B(n_480), .Y(n_597) );
NAND2x1p5_ASAP7_75t_L g598 ( .A(n_494), .B(n_465), .Y(n_598) );
BUFx5_ASAP7_75t_L g599 ( .A(n_526), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_526), .A2(n_477), .B1(n_478), .B2(n_473), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_530), .Y(n_601) );
BUFx3_ASAP7_75t_L g602 ( .A(n_526), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_505), .Y(n_603) );
OR2x2_ASAP7_75t_SL g604 ( .A(n_541), .B(n_362), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_505), .B(n_520), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_514), .Y(n_606) );
OR2x4_ASAP7_75t_L g607 ( .A(n_533), .B(n_477), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_505), .B(n_478), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_524), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_520), .A2(n_341), .B1(n_428), .B2(n_325), .Y(n_610) );
BUFx3_ASAP7_75t_L g611 ( .A(n_494), .Y(n_611) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_516), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_495), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_520), .A2(n_428), .B1(n_398), .B2(n_409), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_524), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_531), .B(n_482), .Y(n_616) );
BUFx3_ASAP7_75t_L g617 ( .A(n_500), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_496), .B(n_306), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_502), .B(n_482), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_531), .B(n_482), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_495), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_500), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_531), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_496), .B(n_504), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_522), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_502), .B(n_486), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_502), .B(n_486), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_495), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_507), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_500), .B(n_465), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_504), .B(n_339), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_502), .B(n_486), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_502), .B(n_488), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_534), .B(n_488), .Y(n_634) );
BUFx8_ASAP7_75t_L g635 ( .A(n_499), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_499), .B(n_391), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_509), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_495), .B(n_500), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_495), .Y(n_639) );
NOR2x1p5_ASAP7_75t_L g640 ( .A(n_541), .B(n_365), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_613), .Y(n_641) );
BUFx2_ASAP7_75t_L g642 ( .A(n_635), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_556), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_619), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_605), .B(n_499), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_619), .A2(n_499), .B1(n_534), .B2(n_541), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_605), .B(n_499), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_619), .Y(n_648) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_545), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_613), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_621), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_565), .A2(n_506), .B1(n_497), .B2(n_503), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_575), .A2(n_534), .B1(n_541), .B2(n_538), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_548), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_556), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_545), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_547), .Y(n_657) );
BUFx8_ASAP7_75t_SL g658 ( .A(n_575), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_565), .B(n_541), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_621), .Y(n_660) );
BUFx12f_ASAP7_75t_L g661 ( .A(n_604), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_638), .A2(n_516), .B(n_527), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_559), .A2(n_497), .B1(n_541), .B2(n_534), .Y(n_663) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_545), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_628), .Y(n_665) );
INVx3_ASAP7_75t_SL g666 ( .A(n_615), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_639), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_554), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_609), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_639), .Y(n_670) );
AND2x4_ASAP7_75t_L g671 ( .A(n_608), .B(n_534), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_568), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_639), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_565), .A2(n_529), .B1(n_503), .B2(n_541), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_608), .Y(n_675) );
CKINVDCx8_ASAP7_75t_R g676 ( .A(n_575), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_545), .B(n_527), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_598), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_609), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_598), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_566), .Y(n_681) );
BUFx3_ASAP7_75t_L g682 ( .A(n_599), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_563), .A2(n_491), .B(n_488), .C(n_529), .Y(n_683) );
BUFx12f_ASAP7_75t_L g684 ( .A(n_604), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_566), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_610), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_566), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_603), .B(n_365), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_634), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_628), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_591), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_626), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_627), .Y(n_693) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_545), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_638), .A2(n_535), .B(n_528), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_594), .Y(n_696) );
BUFx2_ASAP7_75t_L g697 ( .A(n_615), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_597), .B(n_509), .Y(n_698) );
OR2x6_ASAP7_75t_L g699 ( .A(n_575), .B(n_492), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_595), .Y(n_700) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_589), .Y(n_701) );
INVx3_ASAP7_75t_SL g702 ( .A(n_558), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_632), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_583), .B(n_512), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_614), .B(n_398), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_561), .A2(n_512), .B1(n_535), .B2(n_528), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_623), .B(n_537), .Y(n_707) );
INVx4_ASAP7_75t_L g708 ( .A(n_555), .Y(n_708) );
BUFx2_ASAP7_75t_L g709 ( .A(n_557), .Y(n_709) );
INVx3_ASAP7_75t_L g710 ( .A(n_571), .Y(n_710) );
BUFx3_ASAP7_75t_L g711 ( .A(n_599), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_555), .A2(n_532), .B1(n_538), .B2(n_537), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_633), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_607), .B(n_438), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_616), .Y(n_715) );
OR2x6_ASAP7_75t_L g716 ( .A(n_585), .B(n_394), .Y(n_716) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_589), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_577), .A2(n_491), .B1(n_416), .B2(n_409), .C(n_343), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_616), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_596), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_564), .A2(n_532), .B1(n_543), .B2(n_491), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_620), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_598), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_606), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_589), .B(n_543), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g726 ( .A1(n_585), .A2(n_416), .B1(n_436), .B2(n_338), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_625), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_589), .Y(n_728) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_589), .Y(n_729) );
BUFx3_ASAP7_75t_L g730 ( .A(n_599), .Y(n_730) );
NOR2xp67_ASAP7_75t_L g731 ( .A(n_573), .B(n_320), .Y(n_731) );
BUFx12f_ASAP7_75t_L g732 ( .A(n_640), .Y(n_732) );
BUFx2_ASAP7_75t_SL g733 ( .A(n_599), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_630), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_630), .Y(n_735) );
BUFx2_ASAP7_75t_L g736 ( .A(n_557), .Y(n_736) );
INVx3_ASAP7_75t_L g737 ( .A(n_571), .Y(n_737) );
OR2x2_ASAP7_75t_L g738 ( .A(n_560), .B(n_446), .Y(n_738) );
INVx2_ASAP7_75t_SL g739 ( .A(n_630), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_618), .B(n_340), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_564), .B(n_454), .Y(n_741) );
AOI21xp33_ASAP7_75t_L g742 ( .A1(n_551), .A2(n_447), .B(n_403), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_574), .B(n_316), .Y(n_743) );
AO22x1_ASAP7_75t_L g744 ( .A1(n_574), .A2(n_321), .B1(n_329), .B2(n_320), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_612), .B(n_321), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_629), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_612), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_637), .Y(n_748) );
BUFx3_ASAP7_75t_L g749 ( .A(n_599), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_593), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_631), .B(n_396), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_612), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_612), .Y(n_753) );
AND2x4_ASAP7_75t_L g754 ( .A(n_593), .B(n_394), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_607), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_544), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_612), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_602), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_544), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_567), .Y(n_760) );
CKINVDCx11_ASAP7_75t_R g761 ( .A(n_599), .Y(n_761) );
BUFx2_ASAP7_75t_L g762 ( .A(n_607), .Y(n_762) );
BUFx8_ASAP7_75t_L g763 ( .A(n_599), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_571), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_567), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_611), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g767 ( .A1(n_624), .A2(n_448), .B(n_449), .C(n_443), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_546), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_569), .Y(n_769) );
AND3x1_ASAP7_75t_SL g770 ( .A(n_569), .B(n_448), .C(n_443), .Y(n_770) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_611), .Y(n_771) );
INVx3_ASAP7_75t_L g772 ( .A(n_617), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_617), .B(n_449), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_636), .B(n_329), .Y(n_774) );
AND2x4_ASAP7_75t_SL g775 ( .A(n_578), .B(n_450), .Y(n_775) );
INVx6_ASAP7_75t_L g776 ( .A(n_581), .Y(n_776) );
INVx5_ASAP7_75t_L g777 ( .A(n_592), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_546), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_570), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_570), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_622), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_549), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_562), .B(n_336), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_581), .A2(n_536), .B(n_523), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_601), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_691), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_668), .B(n_600), .Y(n_787) );
BUFx4f_ASAP7_75t_SL g788 ( .A(n_732), .Y(n_788) );
INVx3_ASAP7_75t_L g789 ( .A(n_739), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_767), .B(n_581), .C(n_437), .Y(n_790) );
OR2x6_ASAP7_75t_L g791 ( .A(n_642), .B(n_622), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g792 ( .A1(n_657), .A2(n_581), .B1(n_433), .B2(n_397), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_773), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_674), .A2(n_592), .B1(n_551), .B2(n_572), .Y(n_794) );
OR2x6_ASAP7_75t_L g795 ( .A(n_716), .B(n_592), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_784), .A2(n_550), .B(n_549), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_773), .Y(n_797) );
INVx6_ASAP7_75t_L g798 ( .A(n_732), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_643), .B(n_552), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_657), .A2(n_433), .B1(n_345), .B2(n_361), .Y(n_800) );
OR2x2_ASAP7_75t_L g801 ( .A(n_654), .B(n_550), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_715), .B(n_576), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_661), .A2(n_345), .B1(n_361), .B2(n_336), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_696), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_646), .A2(n_584), .B1(n_586), .B2(n_580), .C(n_579), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_686), .A2(n_679), .B1(n_669), .B2(n_659), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_661), .A2(n_410), .B1(n_422), .B2(n_373), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_658), .Y(n_808) );
NAND3xp33_ASAP7_75t_L g809 ( .A(n_767), .B(n_426), .C(n_467), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_722), .B(n_587), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_684), .A2(n_410), .B1(n_422), .B2(n_373), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_696), .Y(n_812) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_678), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_662), .A2(n_590), .B(n_588), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_700), .Y(n_815) );
OR2x6_ASAP7_75t_L g816 ( .A(n_716), .B(n_553), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_686), .A2(n_582), .B1(n_553), .B2(n_310), .Y(n_817) );
AOI222xp33_ASAP7_75t_L g818 ( .A1(n_684), .A2(n_453), .B1(n_450), .B2(n_313), .C1(n_315), .C2(n_318), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_700), .Y(n_819) );
AND2x4_ASAP7_75t_L g820 ( .A(n_719), .B(n_582), .Y(n_820) );
OAI22xp5_ASAP7_75t_SL g821 ( .A1(n_676), .A2(n_441), .B1(n_453), .B2(n_311), .Y(n_821) );
INVxp67_ASAP7_75t_SL g822 ( .A(n_678), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_697), .A2(n_360), .B1(n_367), .B2(n_302), .Y(n_823) );
INVx3_ASAP7_75t_L g824 ( .A(n_739), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_773), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_675), .Y(n_826) );
INVx8_ASAP7_75t_L g827 ( .A(n_716), .Y(n_827) );
OAI22xp5_ASAP7_75t_SL g828 ( .A1(n_676), .A2(n_441), .B1(n_370), .B2(n_379), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_655), .B(n_371), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_705), .A2(n_404), .B1(n_405), .B2(n_382), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_671), .B(n_407), .Y(n_831) );
AO32x2_ASAP7_75t_L g832 ( .A1(n_652), .A2(n_483), .A3(n_467), .B1(n_468), .B2(n_481), .Y(n_832) );
BUFx2_ASAP7_75t_L g833 ( .A(n_680), .Y(n_833) );
INVx4_ASAP7_75t_SL g834 ( .A(n_776), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_688), .B(n_666), .Y(n_835) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_699), .A2(n_348), .B(n_346), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_645), .A2(n_412), .B1(n_413), .B2(n_411), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_724), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_641), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g840 ( .A1(n_677), .A2(n_536), .B(n_523), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_645), .A2(n_419), .B1(n_421), .B2(n_414), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_666), .B(n_429), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_727), .Y(n_843) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_663), .A2(n_357), .B1(n_393), .B2(n_327), .Y(n_844) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_649), .Y(n_845) );
INVx4_ASAP7_75t_L g846 ( .A(n_680), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_658), .Y(n_847) );
INVx1_ASAP7_75t_SL g848 ( .A(n_723), .Y(n_848) );
INVx3_ASAP7_75t_SL g849 ( .A(n_702), .Y(n_849) );
OAI22xp33_ASAP7_75t_L g850 ( .A1(n_718), .A2(n_357), .B1(n_393), .B2(n_327), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_646), .A2(n_342), .B1(n_363), .B2(n_355), .Y(n_851) );
INVx1_ASAP7_75t_SL g852 ( .A(n_723), .Y(n_852) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_681), .Y(n_853) );
AND2x4_ASAP7_75t_L g854 ( .A(n_685), .B(n_434), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_671), .B(n_418), .Y(n_855) );
INVx1_ASAP7_75t_SL g856 ( .A(n_687), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_746), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_748), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g859 ( .A1(n_709), .A2(n_418), .B1(n_374), .B2(n_369), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_671), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_734), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_699), .A2(n_349), .B(n_348), .Y(n_862) );
OAI21x1_ASAP7_75t_L g863 ( .A1(n_728), .A2(n_350), .B(n_349), .Y(n_863) );
NAND3xp33_ASAP7_75t_L g864 ( .A(n_699), .B(n_483), .C(n_467), .Y(n_864) );
OAI21xp5_ASAP7_75t_L g865 ( .A1(n_695), .A2(n_445), .B(n_350), .Y(n_865) );
BUFx6f_ASAP7_75t_L g866 ( .A(n_649), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_776), .A2(n_444), .B1(n_445), .B2(n_330), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_645), .B(n_303), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_755), .Y(n_869) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_649), .Y(n_870) );
BUFx3_ASAP7_75t_L g871 ( .A(n_735), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_720), .Y(n_872) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_751), .A2(n_408), .B1(n_309), .B2(n_312), .C(n_317), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_L g874 ( .A1(n_683), .A2(n_319), .B(n_353), .C(n_308), .Y(n_874) );
INVx3_ASAP7_75t_L g875 ( .A(n_763), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_776), .A2(n_364), .B1(n_366), .B2(n_354), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_647), .A2(n_368), .B1(n_376), .B2(n_372), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_641), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_736), .A2(n_358), .B1(n_400), .B2(n_380), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_647), .A2(n_378), .B1(n_384), .B2(n_381), .Y(n_880) );
NAND3xp33_ASAP7_75t_L g881 ( .A(n_714), .B(n_483), .C(n_387), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_647), .A2(n_385), .B1(n_390), .B2(n_389), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_754), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_754), .Y(n_884) );
OAI22xp33_ASAP7_75t_L g885 ( .A1(n_702), .A2(n_358), .B1(n_399), .B2(n_395), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_775), .A2(n_401), .B1(n_415), .B2(n_402), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_754), .Y(n_887) );
O2A1O1Ixp33_ASAP7_75t_L g888 ( .A1(n_740), .A2(n_420), .B(n_430), .C(n_423), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_653), .B(n_6), .Y(n_889) );
INVx3_ASAP7_75t_L g890 ( .A(n_763), .Y(n_890) );
OR2x6_ASAP7_75t_L g891 ( .A(n_733), .B(n_388), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_650), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_653), .B(n_432), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_650), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_741), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_714), .A2(n_439), .B1(n_456), .B2(n_435), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_644), .Y(n_897) );
INVx1_ASAP7_75t_SL g898 ( .A(n_775), .Y(n_898) );
OAI22xp33_ASAP7_75t_L g899 ( .A1(n_692), .A2(n_424), .B1(n_431), .B2(n_388), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_648), .Y(n_900) );
INVx2_ASAP7_75t_L g901 ( .A(n_651), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_738), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_693), .A2(n_451), .B1(n_400), .B2(n_452), .Y(n_903) );
INVx6_ASAP7_75t_L g904 ( .A(n_777), .Y(n_904) );
CKINVDCx14_ASAP7_75t_R g905 ( .A(n_762), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_726), .B(n_6), .Y(n_906) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_763), .A2(n_400), .B1(n_452), .B2(n_9), .Y(n_907) );
OAI22xp33_ASAP7_75t_L g908 ( .A1(n_703), .A2(n_452), .B1(n_9), .B2(n_7), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_713), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_689), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_698), .B(n_8), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_756), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_741), .A2(n_400), .B1(n_452), .B2(n_468), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_704), .A2(n_781), .B1(n_706), .B2(n_707), .Y(n_914) );
OAI22xp33_ASAP7_75t_L g915 ( .A1(n_758), .A2(n_13), .B1(n_8), .B2(n_10), .Y(n_915) );
OAI22xp5_ASAP7_75t_SL g916 ( .A1(n_774), .A2(n_15), .B1(n_10), .B2(n_14), .Y(n_916) );
OR2x6_ASAP7_75t_L g917 ( .A(n_744), .B(n_476), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_651), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_783), .B(n_14), .Y(n_919) );
NOR2xp67_ASAP7_75t_L g920 ( .A(n_731), .B(n_743), .Y(n_920) );
CKINVDCx16_ASAP7_75t_R g921 ( .A(n_743), .Y(n_921) );
INVx2_ASAP7_75t_SL g922 ( .A(n_743), .Y(n_922) );
INVx2_ASAP7_75t_SL g923 ( .A(n_777), .Y(n_923) );
AOI21xp33_ASAP7_75t_L g924 ( .A1(n_745), .A2(n_16), .B(n_17), .Y(n_924) );
AOI21xp5_ASAP7_75t_L g925 ( .A1(n_677), .A2(n_536), .B(n_523), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_759), .Y(n_926) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_649), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_760), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_758), .A2(n_484), .B1(n_485), .B2(n_481), .Y(n_929) );
OR2x6_ASAP7_75t_L g930 ( .A(n_708), .B(n_484), .Y(n_930) );
INVx2_ASAP7_75t_L g931 ( .A(n_660), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_781), .A2(n_484), .B1(n_487), .B2(n_485), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_660), .Y(n_933) );
INVx4_ASAP7_75t_SL g934 ( .A(n_771), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_765), .A2(n_485), .B1(n_489), .B2(n_487), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_742), .B(n_17), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_750), .B(n_18), .Y(n_937) );
OR2x6_ASAP7_75t_L g938 ( .A(n_708), .B(n_487), .Y(n_938) );
AOI21xp33_ASAP7_75t_L g939 ( .A1(n_745), .A2(n_18), .B(n_19), .Y(n_939) );
NAND2x1p5_ASAP7_75t_L g940 ( .A(n_708), .B(n_489), .Y(n_940) );
NOR2xp67_ASAP7_75t_SL g941 ( .A(n_771), .B(n_750), .Y(n_941) );
INVx3_ASAP7_75t_L g942 ( .A(n_771), .Y(n_942) );
OAI21x1_ASAP7_75t_L g943 ( .A1(n_796), .A2(n_747), .B(n_728), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_902), .B(n_785), .Y(n_944) );
INVx2_ASAP7_75t_SL g945 ( .A(n_827), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_898), .A2(n_771), .B1(n_690), .B2(n_665), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g947 ( .A1(n_898), .A2(n_770), .B1(n_664), .B2(n_694), .Y(n_947) );
AOI22xp33_ASAP7_75t_SL g948 ( .A1(n_827), .A2(n_770), .B1(n_711), .B2(n_730), .Y(n_948) );
OAI211xp5_ASAP7_75t_SL g949 ( .A1(n_818), .A2(n_493), .B(n_489), .C(n_667), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_786), .B(n_665), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_889), .A2(n_769), .B1(n_779), .B2(n_690), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_827), .B(n_768), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_914), .A2(n_772), .B1(n_766), .B2(n_768), .Y(n_953) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_830), .A2(n_721), .B1(n_712), .B2(n_670), .C(n_673), .Y(n_954) );
OR2x2_ASAP7_75t_L g955 ( .A(n_833), .B(n_778), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_790), .A2(n_778), .B1(n_782), .B2(n_777), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_838), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_843), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_909), .B(n_672), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g960 ( .A1(n_891), .A2(n_664), .B1(n_694), .B2(n_656), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_813), .B(n_782), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_790), .A2(n_777), .B1(n_710), .B2(n_737), .Y(n_962) );
OAI211xp5_ASAP7_75t_L g963 ( .A1(n_818), .A2(n_761), .B(n_710), .C(n_737), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_850), .A2(n_672), .B1(n_764), .B2(n_780), .C(n_725), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_916), .A2(n_761), .B1(n_711), .B2(n_730), .Y(n_965) );
AOI21x1_ASAP7_75t_L g966 ( .A1(n_864), .A2(n_725), .B(n_747), .Y(n_966) );
OR2x2_ASAP7_75t_L g967 ( .A(n_853), .B(n_19), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_873), .A2(n_749), .B1(n_682), .B2(n_752), .C(n_757), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_910), .Y(n_969) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_823), .A2(n_749), .B1(n_682), .B2(n_752), .C(n_757), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_857), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_856), .B(n_753), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_806), .A2(n_753), .B1(n_729), .B2(n_717), .C(n_701), .Y(n_973) );
OAI22xp5_ASAP7_75t_SL g974 ( .A1(n_847), .A2(n_664), .B1(n_694), .B2(n_656), .Y(n_974) );
NAND2xp5_ASAP7_75t_SL g975 ( .A(n_836), .B(n_656), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_804), .Y(n_976) );
AND2x4_ASAP7_75t_L g977 ( .A(n_846), .B(n_656), .Y(n_977) );
OAI221xp5_ASAP7_75t_L g978 ( .A1(n_896), .A2(n_717), .B1(n_701), .B2(n_694), .C(n_664), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_844), .A2(n_717), .B1(n_701), .B2(n_729), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_891), .A2(n_729), .B1(n_717), .B2(n_701), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_856), .B(n_729), .Y(n_981) );
OAI21x1_ASAP7_75t_L g982 ( .A1(n_864), .A2(n_493), .B(n_489), .Y(n_982) );
OAI21xp33_ASAP7_75t_L g983 ( .A1(n_907), .A2(n_493), .B(n_483), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_835), .B(n_20), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_921), .B(n_20), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_855), .A2(n_493), .B1(n_483), .B2(n_523), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g987 ( .A(n_860), .B(n_21), .Y(n_987) );
BUFx2_ASAP7_75t_L g988 ( .A(n_795), .Y(n_988) );
OAI21xp33_ASAP7_75t_L g989 ( .A1(n_936), .A2(n_483), .B(n_536), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_842), .A2(n_483), .B1(n_517), .B2(n_511), .Y(n_990) );
NOR2xp33_ASAP7_75t_SL g991 ( .A(n_788), .B(n_22), .Y(n_991) );
OAI22xp33_ASAP7_75t_L g992 ( .A1(n_891), .A2(n_483), .B1(n_25), .B2(n_26), .Y(n_992) );
OA21x2_ASAP7_75t_L g993 ( .A1(n_836), .A2(n_483), .B(n_498), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_893), .A2(n_540), .B1(n_517), .B2(n_511), .Y(n_994) );
INVx2_ASAP7_75t_L g995 ( .A(n_812), .Y(n_995) );
OAI221xp5_ASAP7_75t_L g996 ( .A1(n_837), .A2(n_540), .B1(n_517), .B2(n_511), .C(n_498), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_809), .A2(n_540), .B1(n_517), .B2(n_511), .Y(n_997) );
OA21x2_ASAP7_75t_L g998 ( .A1(n_862), .A2(n_540), .B(n_511), .Y(n_998) );
BUFx4f_ASAP7_75t_L g999 ( .A(n_795), .Y(n_999) );
OAI21xp33_ASAP7_75t_L g1000 ( .A1(n_862), .A2(n_511), .B(n_498), .Y(n_1000) );
BUFx6f_ASAP7_75t_L g1001 ( .A(n_845), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_858), .Y(n_1002) );
OR2x6_ASAP7_75t_L g1003 ( .A(n_795), .B(n_23), .Y(n_1003) );
AO21x2_ASAP7_75t_L g1004 ( .A1(n_865), .A2(n_511), .B(n_498), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_815), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_816), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_809), .A2(n_540), .B1(n_517), .B2(n_511), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_854), .B(n_27), .Y(n_1008) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_848), .B(n_28), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_908), .A2(n_540), .B1(n_517), .B2(n_498), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_852), .B(n_29), .Y(n_1011) );
A2O1A1Ixp33_ASAP7_75t_L g1012 ( .A1(n_888), .A2(n_540), .B(n_517), .C(n_498), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_816), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_906), .A2(n_540), .B1(n_517), .B2(n_498), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_792), .A2(n_498), .B1(n_31), .B2(n_32), .Y(n_1015) );
OAI21xp33_ASAP7_75t_L g1016 ( .A1(n_919), .A2(n_30), .B(n_33), .Y(n_1016) );
BUFx6f_ASAP7_75t_L g1017 ( .A(n_845), .Y(n_1017) );
AOI221xp5_ASAP7_75t_L g1018 ( .A1(n_841), .A2(n_34), .B1(n_35), .B2(n_36), .C(n_37), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1019 ( .A(n_846), .B(n_34), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_872), .Y(n_1020) );
A2O1A1Ixp33_ASAP7_75t_L g1021 ( .A1(n_874), .A2(n_35), .B(n_37), .C(n_38), .Y(n_1021) );
OAI221xp5_ASAP7_75t_L g1022 ( .A1(n_817), .A2(n_39), .B1(n_40), .B2(n_42), .C(n_43), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_852), .Y(n_1023) );
AOI222xp33_ASAP7_75t_L g1024 ( .A1(n_821), .A2(n_39), .B1(n_40), .B2(n_44), .C1(n_45), .C2(n_46), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_861), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_854), .B(n_45), .Y(n_1026) );
BUFx12f_ASAP7_75t_L g1027 ( .A(n_798), .Y(n_1027) );
AOI222xp33_ASAP7_75t_L g1028 ( .A1(n_828), .A2(n_46), .B1(n_47), .B2(n_48), .C1(n_49), .C2(n_50), .Y(n_1028) );
HB1xp67_ASAP7_75t_SL g1029 ( .A(n_808), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_819), .Y(n_1030) );
AOI21x1_ASAP7_75t_L g1031 ( .A1(n_941), .A2(n_118), .B(n_116), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_816), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_912), .Y(n_1033) );
AO31x2_ASAP7_75t_L g1034 ( .A1(n_935), .A2(n_51), .A3(n_52), .B(n_54), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_871), .B(n_55), .Y(n_1035) );
AOI21xp5_ASAP7_75t_L g1036 ( .A1(n_814), .A2(n_925), .B(n_840), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_822), .B(n_57), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_839), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_878), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_911), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_1040) );
NOR2x1_ASAP7_75t_SL g1041 ( .A(n_917), .B(n_62), .Y(n_1041) );
INVx2_ASAP7_75t_L g1042 ( .A(n_892), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_926), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_801), .B(n_64), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_895), .A2(n_65), .B1(n_66), .B2(n_68), .Y(n_1045) );
BUFx12f_ASAP7_75t_L g1046 ( .A(n_798), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_928), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_793), .A2(n_65), .B1(n_66), .B2(n_68), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_886), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_1049) );
OAI21x1_ASAP7_75t_L g1050 ( .A1(n_863), .A2(n_125), .B(n_124), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_826), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_797), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_1052) );
AND2x4_ASAP7_75t_L g1053 ( .A(n_875), .B(n_73), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_849), .B(n_73), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_829), .A2(n_831), .B1(n_859), .B2(n_899), .C(n_882), .Y(n_1055) );
AOI221xp5_ASAP7_75t_L g1056 ( .A1(n_877), .A2(n_74), .B1(n_75), .B2(n_76), .C(n_78), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_825), .A2(n_74), .B1(n_80), .B2(n_81), .Y(n_1057) );
OAI221xp5_ASAP7_75t_L g1058 ( .A1(n_880), .A2(n_80), .B1(n_82), .B2(n_83), .C(n_85), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_915), .A2(n_82), .B1(n_85), .B2(n_86), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_917), .A2(n_86), .B1(n_87), .B2(n_88), .Y(n_1060) );
AOI221x1_ASAP7_75t_SL g1061 ( .A1(n_885), .A2(n_87), .B1(n_88), .B2(n_89), .C(n_90), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_897), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_937), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_820), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_1064) );
AOI22xp33_ASAP7_75t_SL g1065 ( .A1(n_890), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_820), .A2(n_95), .B1(n_96), .B2(n_97), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_900), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_800), .B(n_95), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_894), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_803), .B(n_96), .Y(n_1070) );
OAI22xp33_ASAP7_75t_L g1071 ( .A1(n_917), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_810), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_794), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_1073) );
HB1xp67_ASAP7_75t_L g1074 ( .A(n_901), .Y(n_1074) );
INVx1_ASAP7_75t_SL g1075 ( .A(n_791), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_799), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_807), .B(n_101), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_811), .B(n_101), .Y(n_1078) );
AOI222xp33_ASAP7_75t_L g1079 ( .A1(n_868), .A2(n_787), .B1(n_851), .B2(n_869), .C1(n_802), .C2(n_884), .Y(n_1079) );
INVx2_ASAP7_75t_L g1080 ( .A(n_918), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_802), .A2(n_102), .B1(n_103), .B2(n_104), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_976), .B(n_931), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1025), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_1079), .A2(n_922), .B1(n_890), .B2(n_881), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_1003), .A2(n_881), .B1(n_883), .B2(n_887), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1072), .B(n_905), .Y(n_1086) );
INVx2_ASAP7_75t_L g1087 ( .A(n_993), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1088 ( .A1(n_1061), .A2(n_876), .B1(n_867), .B2(n_939), .C(n_924), .Y(n_1088) );
OAI33xp33_ASAP7_75t_L g1089 ( .A1(n_1071), .A2(n_935), .A3(n_932), .B1(n_933), .B2(n_920), .B3(n_110), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_1003), .A2(n_791), .B1(n_879), .B2(n_865), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_969), .Y(n_1091) );
NAND3xp33_ASAP7_75t_L g1092 ( .A(n_1028), .B(n_913), .C(n_903), .Y(n_1092) );
BUFx3_ASAP7_75t_L g1093 ( .A(n_1027), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_1076), .B(n_957), .Y(n_1094) );
INVx2_ASAP7_75t_L g1095 ( .A(n_993), .Y(n_1095) );
OAI21xp5_ASAP7_75t_L g1096 ( .A1(n_1012), .A2(n_929), .B(n_805), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_993), .Y(n_1097) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_1025), .Y(n_1098) );
OR2x2_ASAP7_75t_L g1099 ( .A(n_1023), .B(n_789), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_995), .B(n_789), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1033), .Y(n_1101) );
AOI222xp33_ASAP7_75t_L g1102 ( .A1(n_985), .A2(n_1055), .B1(n_991), .B2(n_999), .C1(n_1068), .C2(n_1078), .Y(n_1102) );
OA21x2_ASAP7_75t_L g1103 ( .A1(n_943), .A2(n_832), .B(n_923), .Y(n_1103) );
AOI222xp33_ASAP7_75t_L g1104 ( .A1(n_985), .A2(n_834), .B1(n_824), .B2(n_904), .C1(n_934), .C2(n_942), .Y(n_1104) );
AOI22xp33_ASAP7_75t_SL g1105 ( .A1(n_999), .A2(n_824), .B1(n_904), .B2(n_942), .Y(n_1105) );
OAI221xp5_ASAP7_75t_L g1106 ( .A1(n_1059), .A2(n_938), .B1(n_930), .B2(n_940), .C(n_870), .Y(n_1106) );
OAI33xp33_ASAP7_75t_L g1107 ( .A1(n_1071), .A2(n_105), .A3(n_106), .B1(n_107), .B2(n_109), .B3(n_110), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_1003), .A2(n_938), .B1(n_930), .B2(n_940), .Y(n_1108) );
AOI222xp33_ASAP7_75t_L g1109 ( .A1(n_1070), .A2(n_834), .B1(n_934), .B2(n_111), .C1(n_112), .C2(n_109), .Y(n_1109) );
INVx3_ASAP7_75t_L g1110 ( .A(n_977), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_958), .B(n_938), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_998), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_965), .A2(n_927), .B1(n_870), .B2(n_866), .Y(n_1113) );
OAI221xp5_ASAP7_75t_L g1114 ( .A1(n_1015), .A2(n_927), .B1(n_870), .B2(n_866), .C(n_845), .Y(n_1114) );
AOI22xp33_ASAP7_75t_SL g1115 ( .A1(n_1041), .A2(n_927), .B1(n_866), .B2(n_832), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1005), .B(n_832), .Y(n_1116) );
AOI22xp5_ASAP7_75t_L g1117 ( .A1(n_963), .A2(n_107), .B1(n_111), .B2(n_112), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_971), .B(n_131), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1043), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_1023), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_998), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_965), .A2(n_135), .B1(n_139), .B2(n_140), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_955), .Y(n_1123) );
BUFx3_ASAP7_75t_L g1124 ( .A(n_1046), .Y(n_1124) );
INVxp67_ASAP7_75t_SL g1125 ( .A(n_1074), .Y(n_1125) );
AOI22xp5_ASAP7_75t_L g1126 ( .A1(n_1019), .A2(n_141), .B1(n_142), .B2(n_143), .Y(n_1126) );
OA21x2_ASAP7_75t_L g1127 ( .A1(n_956), .A2(n_144), .B(n_146), .Y(n_1127) );
AOI31xp33_ASAP7_75t_L g1128 ( .A1(n_1024), .A2(n_147), .A3(n_148), .B(n_150), .Y(n_1128) );
INVx2_ASAP7_75t_SL g1129 ( .A(n_977), .Y(n_1129) );
OAI211xp5_ASAP7_75t_L g1130 ( .A1(n_1081), .A2(n_152), .B(n_161), .C(n_162), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1047), .Y(n_1131) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_992), .A2(n_166), .B1(n_170), .B2(n_171), .C(n_174), .Y(n_1132) );
AOI221xp5_ASAP7_75t_L g1133 ( .A1(n_992), .A2(n_177), .B1(n_180), .B2(n_181), .C(n_183), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1074), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1030), .B(n_185), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1038), .Y(n_1136) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_953), .A2(n_188), .B1(n_189), .B2(n_192), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_1077), .A2(n_193), .B1(n_195), .B2(n_196), .Y(n_1138) );
AO21x2_ASAP7_75t_L g1139 ( .A1(n_975), .A2(n_198), .B(n_199), .Y(n_1139) );
AOI21xp33_ASAP7_75t_L g1140 ( .A1(n_947), .A2(n_200), .B(n_203), .Y(n_1140) );
OAI211xp5_ASAP7_75t_L g1141 ( .A1(n_1081), .A2(n_204), .B(n_205), .C(n_206), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_1019), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1002), .B(n_299), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_961), .B(n_214), .Y(n_1144) );
AO21x2_ASAP7_75t_L g1145 ( .A1(n_975), .A2(n_216), .B(n_217), .Y(n_1145) );
OR2x6_ASAP7_75t_L g1146 ( .A(n_974), .B(n_218), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1020), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1044), .B(n_219), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1039), .B(n_223), .Y(n_1149) );
NOR2xp33_ASAP7_75t_L g1150 ( .A(n_945), .B(n_225), .Y(n_1150) );
INVx2_ASAP7_75t_L g1151 ( .A(n_998), .Y(n_1151) );
OAI221xp5_ASAP7_75t_L g1152 ( .A1(n_1015), .A2(n_230), .B1(n_231), .B2(n_233), .C(n_239), .Y(n_1152) );
AOI33xp33_ASAP7_75t_L g1153 ( .A1(n_1064), .A2(n_298), .A3(n_246), .B1(n_248), .B2(n_252), .B3(n_254), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1042), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_953), .A2(n_951), .B1(n_948), .B2(n_947), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1004), .Y(n_1156) );
AOI33xp33_ASAP7_75t_L g1157 ( .A1(n_1064), .A2(n_244), .A3(n_255), .B1(n_256), .B2(n_258), .B3(n_259), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_987), .A2(n_261), .B1(n_262), .B2(n_263), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1004), .Y(n_1159) );
INVxp67_ASAP7_75t_L g1160 ( .A(n_967), .Y(n_1160) );
BUFx3_ASAP7_75t_L g1161 ( .A(n_952), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1069), .Y(n_1162) );
BUFx2_ASAP7_75t_L g1163 ( .A(n_960), .Y(n_1163) );
AND2x4_ASAP7_75t_L g1164 ( .A(n_988), .B(n_267), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1080), .B(n_273), .Y(n_1165) );
OAI211xp5_ASAP7_75t_L g1166 ( .A1(n_1065), .A2(n_275), .B(n_277), .C(n_280), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1001), .Y(n_1167) );
OAI22xp33_ASAP7_75t_L g1168 ( .A1(n_1009), .A2(n_1022), .B1(n_1054), .B2(n_1058), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1062), .Y(n_1169) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1001), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_950), .B(n_281), .Y(n_1171) );
AO21x2_ASAP7_75t_L g1172 ( .A1(n_1036), .A2(n_282), .B(n_284), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_1053), .A2(n_285), .B1(n_286), .B2(n_288), .Y(n_1173) );
AOI21xp5_ASAP7_75t_L g1174 ( .A1(n_960), .A2(n_291), .B(n_292), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1075), .B(n_944), .Y(n_1175) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1001), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_1053), .A2(n_294), .B1(n_295), .B2(n_296), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_984), .A2(n_964), .B1(n_1073), .B2(n_951), .Y(n_1178) );
OAI211xp5_ASAP7_75t_L g1179 ( .A1(n_1063), .A2(n_1066), .B(n_1045), .C(n_1048), .Y(n_1179) );
INVxp67_ASAP7_75t_L g1180 ( .A(n_1035), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1067), .B(n_1034), .Y(n_1181) );
OAI211xp5_ASAP7_75t_L g1182 ( .A1(n_1063), .A2(n_1066), .B(n_1045), .C(n_1048), .Y(n_1182) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_1001), .Y(n_1183) );
AOI33xp33_ASAP7_75t_R g1184 ( .A1(n_1083), .A2(n_1006), .A3(n_1032), .B1(n_1013), .B2(n_1049), .B3(n_1060), .Y(n_1184) );
HB1xp67_ASAP7_75t_L g1185 ( .A(n_1098), .Y(n_1185) );
INVx3_ASAP7_75t_L g1186 ( .A(n_1087), .Y(n_1186) );
INVx1_ASAP7_75t_SL g1187 ( .A(n_1093), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1101), .Y(n_1188) );
BUFx2_ASAP7_75t_SL g1189 ( .A(n_1108), .Y(n_1189) );
HB1xp67_ASAP7_75t_L g1190 ( .A(n_1123), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_1090), .A2(n_1057), .B1(n_1052), .B2(n_1010), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1101), .Y(n_1192) );
NAND5xp2_ASAP7_75t_L g1193 ( .A(n_1102), .B(n_1018), .C(n_1056), .D(n_1052), .E(n_1057), .Y(n_1193) );
NAND4xp25_ASAP7_75t_SL g1194 ( .A(n_1109), .B(n_1008), .C(n_1026), .D(n_1037), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1119), .Y(n_1195) );
OAI21xp5_ASAP7_75t_L g1196 ( .A1(n_1128), .A2(n_1021), .B(n_1016), .Y(n_1196) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1112), .Y(n_1197) );
AOI33xp33_ASAP7_75t_L g1198 ( .A1(n_1131), .A2(n_1051), .A3(n_962), .B1(n_956), .B2(n_990), .B3(n_1010), .Y(n_1198) );
INVx2_ASAP7_75t_SL g1199 ( .A(n_1161), .Y(n_1199) );
OAI211xp5_ASAP7_75t_SL g1200 ( .A1(n_1160), .A2(n_1011), .B(n_962), .C(n_1040), .Y(n_1200) );
INVx2_ASAP7_75t_SL g1201 ( .A(n_1161), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1181), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_1155), .A2(n_949), .B1(n_983), .B2(n_954), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1181), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1134), .B(n_1034), .Y(n_1205) );
INVxp67_ASAP7_75t_L g1206 ( .A(n_1086), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1112), .Y(n_1207) );
AND2x4_ASAP7_75t_L g1208 ( .A(n_1110), .B(n_1034), .Y(n_1208) );
CKINVDCx16_ASAP7_75t_R g1209 ( .A(n_1093), .Y(n_1209) );
AND4x1_ASAP7_75t_L g1210 ( .A(n_1104), .B(n_1029), .C(n_990), .D(n_979), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1131), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1169), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1134), .B(n_1034), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1094), .B(n_959), .Y(n_1214) );
AND4x1_ASAP7_75t_L g1215 ( .A(n_1153), .B(n_979), .C(n_1014), .D(n_1000), .Y(n_1215) );
NAND4xp25_ASAP7_75t_L g1216 ( .A(n_1084), .B(n_1014), .C(n_986), .D(n_997), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1125), .B(n_972), .Y(n_1217) );
NAND3xp33_ASAP7_75t_L g1218 ( .A(n_1117), .B(n_986), .C(n_1007), .Y(n_1218) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1120), .B(n_981), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1136), .B(n_1017), .Y(n_1220) );
AND2x2_ASAP7_75t_SL g1221 ( .A(n_1163), .B(n_1017), .Y(n_1221) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1121), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1147), .B(n_946), .Y(n_1223) );
NAND3xp33_ASAP7_75t_L g1224 ( .A(n_1088), .B(n_1007), .C(n_997), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1091), .Y(n_1225) );
AOI21xp5_ASAP7_75t_L g1226 ( .A1(n_1114), .A2(n_980), .B(n_978), .Y(n_1226) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1121), .Y(n_1227) );
OAI31xp33_ASAP7_75t_L g1228 ( .A1(n_1179), .A2(n_973), .A3(n_989), .B(n_996), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1175), .B(n_968), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1175), .Y(n_1230) );
OAI211xp5_ASAP7_75t_L g1231 ( .A1(n_1182), .A2(n_970), .B(n_994), .C(n_1031), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1154), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1154), .B(n_1017), .Y(n_1233) );
OAI21xp5_ASAP7_75t_SL g1234 ( .A1(n_1105), .A2(n_994), .B(n_966), .Y(n_1234) );
AOI331xp33_ASAP7_75t_L g1235 ( .A1(n_1178), .A2(n_982), .A3(n_1050), .B1(n_1085), .B2(n_1162), .B3(n_1113), .C1(n_1173), .Y(n_1235) );
OAI21x1_ASAP7_75t_L g1236 ( .A1(n_1156), .A2(n_1159), .B(n_1151), .Y(n_1236) );
AO21x2_ASAP7_75t_L g1237 ( .A1(n_1156), .A2(n_1159), .B(n_1151), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1162), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1082), .B(n_1087), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1082), .B(n_1095), .Y(n_1240) );
OAI222xp33_ASAP7_75t_L g1241 ( .A1(n_1146), .A2(n_1106), .B1(n_1148), .B2(n_1163), .C1(n_1180), .C2(n_1111), .Y(n_1241) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1095), .Y(n_1242) );
HB1xp67_ASAP7_75t_L g1243 ( .A(n_1099), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1097), .Y(n_1244) );
BUFx2_ASAP7_75t_L g1245 ( .A(n_1146), .Y(n_1245) );
CKINVDCx16_ASAP7_75t_R g1246 ( .A(n_1124), .Y(n_1246) );
INVx2_ASAP7_75t_L g1247 ( .A(n_1097), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1116), .B(n_1110), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1116), .Y(n_1249) );
NAND2xp5_ASAP7_75t_SL g1250 ( .A(n_1115), .B(n_1153), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1148), .B(n_1168), .Y(n_1251) );
AND2x4_ASAP7_75t_L g1252 ( .A(n_1110), .B(n_1176), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1129), .B(n_1100), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1103), .Y(n_1254) );
NOR3xp33_ASAP7_75t_L g1255 ( .A(n_1107), .B(n_1089), .C(n_1092), .Y(n_1255) );
OAI32xp33_ASAP7_75t_L g1256 ( .A1(n_1171), .A2(n_1144), .A3(n_1140), .B1(n_1143), .B2(n_1118), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1100), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_1146), .A2(n_1126), .B1(n_1164), .B2(n_1142), .Y(n_1258) );
NAND4xp25_ASAP7_75t_L g1259 ( .A(n_1251), .B(n_1133), .C(n_1132), .D(n_1157), .Y(n_1259) );
INVx1_ASAP7_75t_SL g1260 ( .A(n_1187), .Y(n_1260) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1202), .B(n_1204), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1188), .Y(n_1262) );
NAND3xp33_ASAP7_75t_SL g1263 ( .A(n_1210), .B(n_1157), .C(n_1177), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1248), .B(n_1183), .Y(n_1264) );
OAI221xp5_ASAP7_75t_L g1265 ( .A1(n_1184), .A2(n_1122), .B1(n_1138), .B2(n_1129), .C(n_1146), .Y(n_1265) );
BUFx2_ASAP7_75t_L g1266 ( .A(n_1245), .Y(n_1266) );
NAND4xp25_ASAP7_75t_L g1267 ( .A(n_1193), .B(n_1158), .C(n_1150), .D(n_1164), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1248), .B(n_1239), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1230), .B(n_1171), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_1194), .A2(n_1164), .B1(n_1152), .B2(n_1096), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1192), .Y(n_1271) );
NAND4xp25_ASAP7_75t_SL g1272 ( .A(n_1209), .B(n_1130), .C(n_1141), .D(n_1166), .Y(n_1272) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1239), .B(n_1176), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1190), .B(n_1167), .Y(n_1274) );
INVx2_ASAP7_75t_L g1275 ( .A(n_1197), .Y(n_1275) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1222), .Y(n_1276) );
INVx3_ASAP7_75t_L g1277 ( .A(n_1186), .Y(n_1277) );
AND2x4_ASAP7_75t_SL g1278 ( .A(n_1199), .B(n_1170), .Y(n_1278) );
NOR2x1_ASAP7_75t_L g1279 ( .A(n_1245), .B(n_1127), .Y(n_1279) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1246), .B(n_1149), .Y(n_1280) );
INVx2_ASAP7_75t_SL g1281 ( .A(n_1201), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1240), .B(n_1170), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_1257), .B(n_1135), .Y(n_1283) );
AOI21xp5_ASAP7_75t_L g1284 ( .A1(n_1258), .A2(n_1127), .B(n_1174), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1195), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1240), .B(n_1127), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1249), .B(n_1205), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1225), .B(n_1149), .Y(n_1288) );
AOI22xp5_ASAP7_75t_L g1289 ( .A1(n_1191), .A2(n_1137), .B1(n_1165), .B2(n_1172), .Y(n_1289) );
INVx2_ASAP7_75t_L g1290 ( .A(n_1222), .Y(n_1290) );
OAI22xp33_ASAP7_75t_L g1291 ( .A1(n_1196), .A2(n_1165), .B1(n_1139), .B2(n_1145), .Y(n_1291) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1243), .B(n_1139), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1213), .B(n_1145), .Y(n_1293) );
OR2x2_ASAP7_75t_L g1294 ( .A(n_1213), .B(n_1145), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1208), .B(n_1186), .Y(n_1295) );
AND2x4_ASAP7_75t_L g1296 ( .A(n_1208), .B(n_1252), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1208), .B(n_1186), .Y(n_1297) );
NAND5xp2_ASAP7_75t_L g1298 ( .A(n_1255), .B(n_1203), .C(n_1228), .D(n_1234), .E(n_1231), .Y(n_1298) );
AND2x2_ASAP7_75t_SL g1299 ( .A(n_1221), .B(n_1189), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1211), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1217), .B(n_1185), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1207), .B(n_1244), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1212), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1232), .B(n_1238), .Y(n_1304) );
AND2x4_ASAP7_75t_L g1305 ( .A(n_1252), .B(n_1242), .Y(n_1305) );
NOR3xp33_ASAP7_75t_L g1306 ( .A(n_1200), .B(n_1241), .C(n_1224), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_1189), .A2(n_1216), .B1(n_1253), .B2(n_1218), .Y(n_1307) );
CKINVDCx16_ASAP7_75t_R g1308 ( .A(n_1253), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1227), .B(n_1247), .Y(n_1309) );
AND2x4_ASAP7_75t_L g1310 ( .A(n_1296), .B(n_1252), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1268), .B(n_1220), .Y(n_1311) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1298), .B(n_1206), .Y(n_1312) );
INVx2_ASAP7_75t_SL g1313 ( .A(n_1278), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1301), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1271), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1287), .B(n_1219), .Y(n_1316) );
NOR2x1_ASAP7_75t_L g1317 ( .A(n_1260), .B(n_1250), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1308), .B(n_1219), .Y(n_1318) );
INVx2_ASAP7_75t_SL g1319 ( .A(n_1278), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1285), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1261), .B(n_1229), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1285), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1295), .B(n_1247), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1264), .B(n_1220), .Y(n_1324) );
NAND4xp25_ASAP7_75t_L g1325 ( .A(n_1306), .B(n_1198), .C(n_1214), .D(n_1226), .Y(n_1325) );
NOR2xp33_ASAP7_75t_L g1326 ( .A(n_1267), .B(n_1256), .Y(n_1326) );
OAI22xp5_ASAP7_75t_SL g1327 ( .A1(n_1280), .A2(n_1235), .B1(n_1223), .B2(n_1215), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1300), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1273), .B(n_1237), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1303), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1273), .B(n_1237), .Y(n_1331) );
NAND3xp33_ASAP7_75t_L g1332 ( .A(n_1307), .B(n_1233), .C(n_1254), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1303), .B(n_1237), .Y(n_1333) );
OA22x2_ASAP7_75t_L g1334 ( .A1(n_1266), .A2(n_1236), .B1(n_1254), .B2(n_1256), .Y(n_1334) );
AO21x1_ASAP7_75t_L g1335 ( .A1(n_1284), .A2(n_1236), .B(n_1291), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_1263), .A2(n_1270), .B1(n_1259), .B2(n_1265), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1262), .Y(n_1337) );
A2O1A1Ixp33_ASAP7_75t_L g1338 ( .A1(n_1279), .A2(n_1299), .B(n_1266), .C(n_1289), .Y(n_1338) );
NAND4xp25_ASAP7_75t_L g1339 ( .A(n_1269), .B(n_1274), .C(n_1288), .D(n_1283), .Y(n_1339) );
NAND2x1_ASAP7_75t_L g1340 ( .A(n_1281), .B(n_1305), .Y(n_1340) );
XNOR2x2_ASAP7_75t_L g1341 ( .A(n_1317), .B(n_1304), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1337), .Y(n_1342) );
INVxp67_ASAP7_75t_L g1343 ( .A(n_1312), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1315), .Y(n_1344) );
OAI22xp33_ASAP7_75t_SL g1345 ( .A1(n_1340), .A2(n_1292), .B1(n_1294), .B2(n_1293), .Y(n_1345) );
XOR2x2_ASAP7_75t_L g1346 ( .A(n_1318), .B(n_1299), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1347 ( .A(n_1314), .B(n_1282), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1320), .Y(n_1348) );
NOR2xp33_ASAP7_75t_L g1349 ( .A(n_1325), .B(n_1296), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1311), .B(n_1295), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1322), .Y(n_1351) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_1313), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1321), .B(n_1282), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1316), .B(n_1329), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1339), .B(n_1302), .Y(n_1355) );
NOR2xp67_ASAP7_75t_L g1356 ( .A(n_1319), .B(n_1272), .Y(n_1356) );
AND3x1_ASAP7_75t_L g1357 ( .A(n_1336), .B(n_1297), .C(n_1286), .Y(n_1357) );
INVxp67_ASAP7_75t_SL g1358 ( .A(n_1331), .Y(n_1358) );
AND2x4_ASAP7_75t_L g1359 ( .A(n_1310), .B(n_1296), .Y(n_1359) );
XOR2x2_ASAP7_75t_L g1360 ( .A(n_1326), .B(n_1305), .Y(n_1360) );
OA21x2_ASAP7_75t_L g1361 ( .A1(n_1335), .A2(n_1294), .B(n_1276), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1328), .Y(n_1362) );
NOR2xp67_ASAP7_75t_L g1363 ( .A(n_1332), .B(n_1277), .Y(n_1363) );
CKINVDCx5p33_ASAP7_75t_R g1364 ( .A(n_1327), .Y(n_1364) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_1324), .B(n_1277), .Y(n_1365) );
A2O1A1Ixp33_ASAP7_75t_L g1366 ( .A1(n_1338), .A2(n_1277), .B(n_1309), .C(n_1275), .Y(n_1366) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1330), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1333), .Y(n_1368) );
AOI222xp33_ASAP7_75t_L g1369 ( .A1(n_1338), .A2(n_1275), .B1(n_1276), .B2(n_1290), .C1(n_1323), .C2(n_1310), .Y(n_1369) );
CKINVDCx20_ASAP7_75t_R g1370 ( .A(n_1364), .Y(n_1370) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1354), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1354), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1355), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1367), .Y(n_1374) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1367), .Y(n_1375) );
AOI22xp5_ASAP7_75t_L g1376 ( .A1(n_1364), .A2(n_1357), .B1(n_1343), .B2(n_1349), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1359), .B(n_1352), .Y(n_1377) );
AOI21xp5_ASAP7_75t_L g1378 ( .A1(n_1366), .A2(n_1356), .B(n_1369), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1368), .B(n_1342), .Y(n_1379) );
BUFx2_ASAP7_75t_L g1380 ( .A(n_1352), .Y(n_1380) );
XNOR2x1_ASAP7_75t_L g1381 ( .A(n_1346), .B(n_1360), .Y(n_1381) );
OAI21xp5_ASAP7_75t_L g1382 ( .A1(n_1378), .A2(n_1363), .B(n_1334), .Y(n_1382) );
AOI221x1_ASAP7_75t_L g1383 ( .A1(n_1378), .A2(n_1345), .B1(n_1368), .B2(n_1344), .C(n_1351), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1373), .B(n_1358), .Y(n_1384) );
OAI21xp33_ASAP7_75t_SL g1385 ( .A1(n_1381), .A2(n_1363), .B(n_1350), .Y(n_1385) );
HB1xp67_ASAP7_75t_L g1386 ( .A(n_1380), .Y(n_1386) );
OAI211xp5_ASAP7_75t_L g1387 ( .A1(n_1376), .A2(n_1361), .B(n_1341), .C(n_1365), .Y(n_1387) );
INVx2_ASAP7_75t_L g1388 ( .A(n_1374), .Y(n_1388) );
NAND2xp5_ASAP7_75t_SL g1389 ( .A(n_1370), .B(n_1359), .Y(n_1389) );
NAND3xp33_ASAP7_75t_L g1390 ( .A(n_1383), .B(n_1370), .C(n_1361), .Y(n_1390) );
AO22x2_ASAP7_75t_L g1391 ( .A1(n_1389), .A2(n_1372), .B1(n_1371), .B2(n_1377), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1386), .B(n_1379), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1384), .B(n_1375), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1387), .B(n_1361), .Y(n_1394) );
AO22x2_ASAP7_75t_L g1395 ( .A1(n_1390), .A2(n_1382), .B1(n_1388), .B2(n_1385), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1392), .Y(n_1396) );
OAI21xp5_ASAP7_75t_L g1397 ( .A1(n_1394), .A2(n_1359), .B(n_1353), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1397), .B(n_1391), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1396), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1395), .Y(n_1400) );
AOI22x1_ASAP7_75t_L g1401 ( .A1(n_1395), .A2(n_1391), .B1(n_1393), .B2(n_1347), .Y(n_1401) );
INVx2_ASAP7_75t_L g1402 ( .A(n_1401), .Y(n_1402) );
AOI22xp5_ASAP7_75t_L g1403 ( .A1(n_1402), .A2(n_1400), .B1(n_1398), .B2(n_1399), .Y(n_1403) );
INVx2_ASAP7_75t_L g1404 ( .A(n_1403), .Y(n_1404) );
AOI21xp5_ASAP7_75t_L g1405 ( .A1(n_1404), .A2(n_1348), .B(n_1362), .Y(n_1405) );
endmodule