module real_jpeg_30379_n_5 (n_4, n_0, n_1, n_2, n_3, n_5);

input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_5;

wire n_17;
wire n_12;
wire n_8;
wire n_18;
wire n_11;
wire n_10;
wire n_14;
wire n_6;
wire n_7;
wire n_16;
wire n_15;
wire n_13;
wire n_9;

INVx4_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

AOI211xp5_ASAP7_75t_L g10 ( 
.A1(n_1),
.A2(n_11),
.B(n_13),
.C(n_15),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_17),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_12),
.Y(n_14)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

OA22x2_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_L g5 ( 
.A1(n_6),
.A2(n_7),
.B1(n_10),
.B2(n_18),
.Y(n_5)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);


endmodule