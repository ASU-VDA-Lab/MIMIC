module fake_jpeg_17697_n_198 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_11),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_30),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_50),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_14),
.B1(n_27),
.B2(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_43),
.B1(n_52),
.B2(n_22),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_14),
.B1(n_27),
.B2(n_25),
.Y(n_43)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_28),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_30),
.A2(n_23),
.B1(n_15),
.B2(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_57),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_35),
.B1(n_32),
.B2(n_15),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_40),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_16),
.B(n_21),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_1),
.B(n_2),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_68),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_23),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_19),
.C(n_18),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_16),
.C(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_73),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_15),
.B1(n_21),
.B2(n_33),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_40),
.B1(n_47),
.B2(n_46),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_21),
.B(n_25),
.C(n_24),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_77),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_75),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_48),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_28),
.B(n_24),
.C(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_22),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_65),
.B1(n_70),
.B2(n_74),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_78),
.B1(n_56),
.B2(n_61),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_90),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_38),
.B(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_99),
.B1(n_47),
.B2(n_55),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_88),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_40),
.B(n_47),
.C(n_37),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_60),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_40),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_55),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_102),
.B1(n_59),
.B2(n_37),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_72),
.B(n_66),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_46),
.Y(n_120)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_54),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_114),
.B(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_111),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_90),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_55),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_120),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_92),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_88),
.B1(n_97),
.B2(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_59),
.B1(n_46),
.B2(n_19),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_125),
.B1(n_103),
.B2(n_18),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_19),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_19),
.B1(n_18),
.B2(n_17),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_82),
.B(n_99),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_126),
.A2(n_5),
.B(n_6),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_113),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_101),
.C(n_98),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_137),
.C(n_140),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_108),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_80),
.B(n_92),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_98),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_143),
.B1(n_144),
.B2(n_7),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_96),
.C(n_85),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_95),
.C(n_97),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_2),
.C(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_150),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_155),
.B(n_138),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_119),
.Y(n_150)
);

AOI221xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_111),
.B1(n_122),
.B2(n_123),
.C(n_105),
.Y(n_151)
);

OA21x2_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_156),
.B(n_139),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_140),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_2),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_142),
.Y(n_160)
);

AOI221xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_128),
.B(n_139),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_8),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_7),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_163),
.C(n_145),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g162 ( 
.A(n_155),
.B(n_144),
.C(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_166),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_134),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_139),
.B1(n_132),
.B2(n_152),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_168),
.B(n_141),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_175),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_153),
.B(n_129),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_171),
.B1(n_158),
.B2(n_11),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_130),
.B1(n_153),
.B2(n_145),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_174),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_143),
.B1(n_154),
.B2(n_9),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_177),
.C(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_163),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_10),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_182),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_171),
.B(n_160),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_184),
.C(n_170),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_178),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_186),
.Y(n_193)
);

NAND2x1_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_158),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_179),
.C(n_183),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_187),
.B(n_10),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_192),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_193),
.C(n_190),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_191),
.Y(n_197)
);


endmodule