module real_jpeg_19006_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_0),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_1),
.A2(n_54),
.B1(n_65),
.B2(n_72),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_54),
.Y(n_193)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_3),
.A2(n_65),
.B1(n_72),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_3),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_53),
.B1(n_55),
.B2(n_94),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_94),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_94),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_4),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_5),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_5),
.A2(n_53),
.B1(n_55),
.B2(n_73),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_73),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_73),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_6),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_6),
.A2(n_53),
.B(n_70),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_65),
.B1(n_72),
.B2(n_142),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_75),
.Y(n_190)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_6),
.A2(n_37),
.B(n_41),
.C(n_203),
.D(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_37),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_6),
.B(n_59),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_6),
.A2(n_25),
.B(n_218),
.Y(n_236)
);

A2O1A1O1Ixp25_ASAP7_75t_L g249 ( 
.A1(n_6),
.A2(n_55),
.B(n_56),
.C(n_151),
.D(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_6),
.B(n_55),
.Y(n_250)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_8),
.B(n_219),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_11),
.A2(n_65),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_11),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_11),
.A2(n_53),
.B1(n_55),
.B2(n_77),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_77),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_77),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_12),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_39),
.B1(n_53),
.B2(n_55),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_39),
.Y(n_145)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_15),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_20),
.B(n_102),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_85),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_21),
.A2(n_22),
.B1(n_78),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_23),
.B(n_51),
.C(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_24),
.B(n_35),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_25),
.A2(n_33),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_25),
.A2(n_81),
.B1(n_88),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_25),
.A2(n_81),
.B1(n_145),
.B2(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_25),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_25),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_26),
.A2(n_224),
.B(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_29),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_27),
.A2(n_43),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_29),
.B(n_42),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_29),
.B(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_31),
.A2(n_193),
.B(n_233),
.Y(n_257)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_36),
.A2(n_40),
.B1(n_48),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_38),
.B1(n_57),
.B2(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_37),
.B(n_57),
.Y(n_256)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_38),
.A2(n_58),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_40),
.A2(n_46),
.B1(n_48),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_40),
.A2(n_48),
.B1(n_215),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_40),
.A2(n_248),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_41),
.A2(n_44),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_41),
.B(n_167),
.Y(n_166)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_48),
.A2(n_90),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_48),
.B(n_168),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_48),
.A2(n_166),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_48),
.B(n_142),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B1(n_59),
.B2(n_61),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_57),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_55),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_56),
.A2(n_59),
.B1(n_61),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_74),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_65),
.A2(n_67),
.B(n_142),
.C(n_143),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_69),
.A2(n_93),
.B(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_74),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_80),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_82),
.Y(n_117)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_81),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_81),
.B(n_142),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_85),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.C(n_95),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_87),
.B(n_89),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_101),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_98),
.A2(n_148),
.B1(n_149),
.B2(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_98),
.A2(n_99),
.B(n_174),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_125),
.B2(n_126),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_114),
.B2(n_115),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_111),
.B(n_113),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_111),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_124),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_123),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_125),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_155),
.B(n_282),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_152),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_131),
.B(n_152),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_135),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_134),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_136),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.C(n_146),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_138),
.B1(n_146),
.B2(n_147),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B(n_150),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_195),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_178),
.B(n_194),
.Y(n_157)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_158),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_175),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_175),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.C(n_172),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_165),
.B1(n_172),
.B2(n_173),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_179),
.B(n_181),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_186),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_182),
.B(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_184),
.A2(n_186),
.B1(n_187),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_184),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_188),
.A2(n_189),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_190),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_280),
.C(n_281),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_274),
.B(n_279),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_260),
.B(n_273),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_242),
.B(n_259),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_220),
.B(n_241),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_209),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_201),
.B(n_209),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_205),
.B1(n_206),
.B2(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_216),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_217),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_219),
.B(n_225),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_230),
.B(n_240),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_222),
.B(n_228),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_235),
.B(n_239),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_244),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_253),
.B2(n_258),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_252),
.C(n_258),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_253),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_257),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_262),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_269),
.C(n_271),
.Y(n_275)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);


endmodule