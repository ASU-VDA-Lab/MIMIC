module real_aes_15800_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_953, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_953;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_905;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_298;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_947;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_617;
wire n_552;
wire n_402;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_0), .Y(n_197) );
AND2x4_ASAP7_75t_L g946 ( .A(n_1), .B(n_947), .Y(n_946) );
BUFx3_ASAP7_75t_L g242 ( .A(n_2), .Y(n_242) );
INVx1_ASAP7_75t_L g947 ( .A(n_3), .Y(n_947) );
AOI22xp5_ASAP7_75t_SL g913 ( .A1(n_4), .A2(n_914), .B1(n_915), .B2(n_916), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_4), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_5), .B(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_L g114 ( .A(n_6), .B(n_23), .Y(n_114) );
BUFx2_ASAP7_75t_L g940 ( .A(n_6), .Y(n_940) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_7), .Y(n_138) );
OAI22xp5_ASAP7_75t_R g910 ( .A1(n_8), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_8), .Y(n_911) );
CKINVDCx5p33_ASAP7_75t_R g928 ( .A(n_9), .Y(n_928) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_10), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g512 ( .A(n_11), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_11), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_12), .B(n_152), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_13), .B(n_157), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_14), .A2(n_84), .B1(n_152), .B2(n_166), .Y(n_251) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_15), .A2(n_36), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_16), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_17), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_18), .Y(n_557) );
AO32x1_ASAP7_75t_L g248 ( .A1(n_19), .A2(n_130), .A3(n_177), .B1(n_220), .B2(n_249), .Y(n_248) );
AO32x2_ASAP7_75t_L g283 ( .A1(n_19), .A2(n_130), .A3(n_177), .B1(n_220), .B2(n_249), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_20), .B(n_573), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_21), .B(n_177), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_22), .Y(n_662) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_23), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_24), .A2(n_43), .B1(n_140), .B2(n_150), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_25), .B(n_171), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_26), .A2(n_93), .B1(n_166), .B2(n_172), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_27), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_28), .B(n_212), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_29), .A2(n_64), .B1(n_172), .B2(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_30), .B(n_152), .Y(n_627) );
INVx2_ASAP7_75t_L g531 ( .A(n_31), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_32), .B(n_169), .Y(n_615) );
INVx1_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
BUFx3_ASAP7_75t_L g926 ( .A(n_33), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_34), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_35), .B(n_565), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_37), .Y(n_107) );
AND2x2_ASAP7_75t_L g564 ( .A(n_38), .B(n_565), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_39), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_40), .B(n_198), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_41), .B(n_573), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_42), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_44), .B(n_667), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_45), .A2(n_78), .B1(n_198), .B2(n_212), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_46), .A2(n_519), .B1(n_520), .B2(n_521), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_46), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_47), .B(n_264), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_48), .A2(n_141), .B(n_195), .C(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_49), .A2(n_80), .B1(n_152), .B2(n_166), .Y(n_238) );
INVx1_ASAP7_75t_L g132 ( .A(n_50), .Y(n_132) );
AND2x4_ASAP7_75t_L g154 ( .A(n_51), .B(n_155), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_52), .A2(n_53), .B1(n_150), .B2(n_172), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_54), .B(n_177), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_55), .B(n_565), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_56), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_57), .A2(n_105), .B1(n_936), .B2(n_950), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_58), .B(n_172), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_59), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_61), .B(n_177), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_62), .A2(n_195), .B(n_196), .C(n_199), .Y(n_194) );
NAND3xp33_ASAP7_75t_L g175 ( .A(n_63), .B(n_166), .C(n_174), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_65), .Y(n_638) );
OAI22xp5_ASAP7_75t_SL g521 ( .A1(n_66), .A2(n_88), .B1(n_522), .B2(n_523), .Y(n_521) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_66), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_66), .B(n_177), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_67), .B(n_562), .Y(n_571) );
AND2x2_ASAP7_75t_L g201 ( .A(n_68), .B(n_202), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_69), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_70), .A2(n_82), .B1(n_917), .B2(n_918), .Y(n_916) );
INVx1_ASAP7_75t_L g918 ( .A(n_70), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_71), .B(n_140), .C(n_169), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_72), .A2(n_96), .B1(n_152), .B2(n_198), .Y(n_229) );
INVx2_ASAP7_75t_L g143 ( .A(n_73), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_74), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_75), .B(n_562), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_76), .B(n_193), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_77), .B(n_152), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_79), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_81), .B(n_146), .Y(n_602) );
INVx1_ASAP7_75t_L g917 ( .A(n_82), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_83), .A2(n_92), .B1(n_573), .B2(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_85), .B(n_152), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_86), .B(n_174), .Y(n_173) );
NAND2xp33_ASAP7_75t_SL g588 ( .A(n_87), .B(n_168), .Y(n_588) );
INVx1_ASAP7_75t_L g522 ( .A(n_88), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_89), .B(n_137), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_90), .A2(n_103), .B1(n_150), .B2(n_172), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_91), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_94), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g907 ( .A(n_94), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_95), .B(n_157), .Y(n_222) );
NAND2xp33_ASAP7_75t_L g600 ( .A(n_97), .B(n_168), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_98), .B(n_565), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_99), .B(n_168), .C(n_193), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_100), .B(n_562), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_101), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_102), .B(n_573), .Y(n_576) );
OR2x6_ASAP7_75t_L g105 ( .A(n_106), .B(n_115), .Y(n_105) );
INVx1_ASAP7_75t_L g524 ( .A(n_106), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_106), .B(n_518), .Y(n_537) );
NOR2xp67_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .Y(n_106) );
CKINVDCx8_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
INVx5_ASAP7_75t_L g535 ( .A(n_109), .Y(n_535) );
AND2x6_ASAP7_75t_SL g109 ( .A(n_110), .B(n_113), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_112), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_113), .B(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2x1_ASAP7_75t_L g935 ( .A(n_114), .B(n_926), .Y(n_935) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_116), .B(n_538), .Y(n_115) );
AOI32xp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_118), .A3(n_515), .B1(n_525), .B2(n_536), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_512), .B(n_513), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NOR2xp33_ASAP7_75t_SL g513 ( .A(n_121), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g908 ( .A(n_121), .Y(n_908) );
NAND2x1p5_ASAP7_75t_L g121 ( .A(n_122), .B(n_386), .Y(n_121) );
AND5x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_312), .C(n_332), .D(n_348), .E(n_368), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_272), .Y(n_123) );
OAI21xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_178), .B(n_243), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g380 ( .A(n_126), .Y(n_380) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g366 ( .A(n_127), .Y(n_366) );
OR2x2_ASAP7_75t_L g403 ( .A(n_127), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g469 ( .A(n_127), .B(n_223), .Y(n_469) );
OR2x2_ASAP7_75t_L g478 ( .A(n_127), .B(n_297), .Y(n_478) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_160), .Y(n_127) );
BUFx2_ASAP7_75t_L g255 ( .A(n_128), .Y(n_255) );
INVx1_ASAP7_75t_L g271 ( .A(n_128), .Y(n_271) );
INVx2_ASAP7_75t_SL g330 ( .A(n_128), .Y(n_330) );
AND2x2_ASAP7_75t_L g351 ( .A(n_128), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g455 ( .A(n_128), .B(n_224), .Y(n_455) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B(n_156), .Y(n_128) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_129), .A2(n_133), .B(n_156), .Y(n_295) );
OAI21x1_ASAP7_75t_L g612 ( .A1(n_129), .A2(n_613), .B(n_621), .Y(n_612) );
OAI21x1_ASAP7_75t_L g623 ( .A1(n_129), .A2(n_624), .B(n_631), .Y(n_623) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_129), .A2(n_624), .B(n_631), .Y(n_645) );
OA21x2_ASAP7_75t_L g690 ( .A1(n_129), .A2(n_613), .B(n_621), .Y(n_690) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx4_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
INVx2_ASAP7_75t_SL g208 ( .A(n_130), .Y(n_208) );
BUFx3_ASAP7_75t_L g225 ( .A(n_130), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_130), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_130), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_SL g581 ( .A(n_130), .Y(n_581) );
AND2x4_ASAP7_75t_SL g605 ( .A(n_130), .B(n_153), .Y(n_605) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_144), .B(n_153), .Y(n_133) );
O2A1O1Ixp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_139), .C(n_141), .Y(n_134) );
O2A1O1Ixp5_ASAP7_75t_L g661 ( .A1(n_136), .A2(n_169), .B(n_662), .C(n_663), .Y(n_661) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_138), .Y(n_140) );
INVx1_ASAP7_75t_L g150 ( .A(n_138), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_138), .Y(n_152) );
INVx2_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
INVx1_ASAP7_75t_L g195 ( .A(n_138), .Y(n_195) );
INVx1_ASAP7_75t_L g198 ( .A(n_138), .Y(n_198) );
INVx3_ASAP7_75t_L g562 ( .A(n_138), .Y(n_562) );
INVx1_ASAP7_75t_L g574 ( .A(n_138), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_140), .A2(n_150), .B1(n_190), .B2(n_191), .Y(n_189) );
INVx2_ASAP7_75t_L g264 ( .A(n_140), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_141), .A2(n_169), .B1(n_250), .B2(n_251), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_141), .A2(n_571), .B(n_572), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_141), .A2(n_587), .B(n_588), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_141), .A2(n_599), .B(n_600), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_141), .A2(n_626), .B(n_627), .Y(n_625) );
BUFx4f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g148 ( .A(n_143), .Y(n_148) );
BUFx8_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
INVx1_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_147), .B1(n_149), .B2(n_151), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_146), .A2(n_665), .B(n_666), .Y(n_664) );
INVx2_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_147), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_601) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx3_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g218 ( .A(n_152), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_152), .A2(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g620 ( .A(n_152), .Y(n_620) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_153), .A2(n_164), .B(n_170), .Y(n_163) );
AOI31xp67_ASAP7_75t_L g235 ( .A1(n_153), .A2(n_236), .A3(n_237), .B(n_240), .Y(n_235) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_153), .A2(n_570), .B(n_575), .Y(n_569) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_153), .A2(n_583), .B(n_586), .Y(n_582) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_153), .A2(n_614), .B(n_617), .Y(n_613) );
OAI21x1_ASAP7_75t_L g624 ( .A1(n_153), .A2(n_625), .B(n_628), .Y(n_624) );
OAI21x1_ASAP7_75t_L g660 ( .A1(n_153), .A2(n_661), .B(n_664), .Y(n_660) );
BUFx10_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g200 ( .A(n_154), .Y(n_200) );
INVx1_ASAP7_75t_L g221 ( .A(n_154), .Y(n_221) );
AO31x2_ASAP7_75t_L g261 ( .A1(n_154), .A2(n_225), .A3(n_262), .B(n_266), .Y(n_261) );
BUFx10_ASAP7_75t_L g553 ( .A(n_154), .Y(n_553) );
INVx2_ASAP7_75t_L g186 ( .A(n_157), .Y(n_186) );
NOR2xp67_ASAP7_75t_SL g551 ( .A(n_157), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AO31x2_ASAP7_75t_L g632 ( .A1(n_158), .A2(n_553), .A3(n_633), .B(n_637), .Y(n_632) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g162 ( .A(n_159), .Y(n_162) );
INVx2_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
AND2x2_ASAP7_75t_L g311 ( .A(n_160), .B(n_295), .Y(n_311) );
AND2x2_ASAP7_75t_L g421 ( .A(n_160), .B(n_279), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_176), .Y(n_160) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_161), .A2(n_163), .B(n_176), .Y(n_258) );
OAI21x1_ASAP7_75t_L g568 ( .A1(n_161), .A2(n_569), .B(n_578), .Y(n_568) );
OAI21xp33_ASAP7_75t_SL g607 ( .A1(n_161), .A2(n_569), .B(n_578), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g659 ( .A1(n_161), .A2(n_660), .B(n_668), .Y(n_659) );
OAI21x1_ASAP7_75t_L g687 ( .A1(n_161), .A2(n_660), .B(n_668), .Y(n_687) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g565 ( .A(n_162), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_167), .B(n_169), .Y(n_164) );
INVx2_ASAP7_75t_SL g212 ( .A(n_166), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_166), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g667 ( .A(n_168), .Y(n_667) );
INVx6_ASAP7_75t_L g219 ( .A(n_169), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_169), .A2(n_219), .B1(n_238), .B2(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_169), .A2(n_629), .B(n_630), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_175), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_172), .A2(n_561), .B1(n_562), .B2(n_563), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_172), .A2(n_615), .B(n_616), .Y(n_614) );
INVx2_ASAP7_75t_L g635 ( .A(n_172), .Y(n_635) );
INVx2_ASAP7_75t_L g236 ( .A(n_177), .Y(n_236) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2x1_ASAP7_75t_L g179 ( .A(n_180), .B(n_204), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_182), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g355 ( .A(n_183), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_184), .Y(n_253) );
AND2x2_ASAP7_75t_L g285 ( .A(n_184), .B(n_261), .Y(n_285) );
INVx1_ASAP7_75t_L g289 ( .A(n_184), .Y(n_289) );
INVx1_ASAP7_75t_L g327 ( .A(n_184), .Y(n_327) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g268 ( .A(n_185), .Y(n_268) );
AOI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_201), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_194), .B(n_200), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_189), .B(n_192), .Y(n_188) );
AOI21x1_ASAP7_75t_L g617 ( .A1(n_192), .A2(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_SL g228 ( .A(n_193), .Y(n_228) );
INVx1_ASAP7_75t_L g603 ( .A(n_195), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx2_ASAP7_75t_L g214 ( .A(n_199), .Y(n_214) );
INVx2_ASAP7_75t_L g559 ( .A(n_199), .Y(n_559) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_203), .B(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_203), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_223), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_205), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g252 ( .A(n_206), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g281 ( .A(n_206), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g290 ( .A(n_206), .Y(n_290) );
INVx3_ASAP7_75t_L g302 ( .A(n_206), .Y(n_302) );
BUFx2_ASAP7_75t_L g340 ( .A(n_206), .Y(n_340) );
INVxp67_ASAP7_75t_L g360 ( .A(n_206), .Y(n_360) );
AND2x2_ASAP7_75t_L g383 ( .A(n_206), .B(n_283), .Y(n_383) );
INVx1_ASAP7_75t_L g397 ( .A(n_206), .Y(n_397) );
OR2x2_ASAP7_75t_L g418 ( .A(n_206), .B(n_282), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_206), .B(n_261), .Y(n_474) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OAI21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_222), .Y(n_207) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_215), .B(n_220), .Y(n_209) );
AOI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_213), .B(n_214), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_214), .A2(n_219), .B1(n_263), .B2(n_265), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_214), .A2(n_576), .B(n_577), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_219), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_219), .A2(n_227), .B1(n_228), .B2(n_229), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_219), .A2(n_559), .B1(n_634), .B2(n_636), .Y(n_633) );
INVx2_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_SL g230 ( .A(n_221), .Y(n_230) );
INVx1_ASAP7_75t_L g385 ( .A(n_223), .Y(n_385) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_233), .Y(n_223) );
AND2x2_ASAP7_75t_L g270 ( .A(n_224), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g297 ( .A(n_224), .Y(n_297) );
INVx2_ASAP7_75t_L g316 ( .A(n_224), .Y(n_316) );
AND2x2_ASAP7_75t_L g331 ( .A(n_224), .B(n_279), .Y(n_331) );
INVx1_ASAP7_75t_L g352 ( .A(n_224), .Y(n_352) );
AND2x2_ASAP7_75t_L g410 ( .A(n_224), .B(n_233), .Y(n_410) );
AND2x2_ASAP7_75t_L g420 ( .A(n_224), .B(n_295), .Y(n_420) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .A3(n_230), .B(n_231), .Y(n_224) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g257 ( .A(n_234), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g279 ( .A(n_235), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_242), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_254), .B1(n_259), .B2(n_269), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_244), .A2(n_472), .B1(n_476), .B2(n_477), .Y(n_471) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_252), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_245), .B(n_285), .Y(n_376) );
NAND2xp5_ASAP7_75t_R g395 ( .A(n_245), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g407 ( .A(n_247), .B(n_302), .Y(n_407) );
INVx1_ASAP7_75t_L g475 ( .A(n_247), .Y(n_475) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g303 ( .A(n_248), .B(n_261), .Y(n_303) );
OR2x2_ASAP7_75t_L g344 ( .A(n_248), .B(n_261), .Y(n_344) );
INVx1_ASAP7_75t_L g356 ( .A(n_248), .Y(n_356) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_252), .Y(n_498) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g313 ( .A(n_255), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_255), .B(n_331), .Y(n_347) );
INVx1_ASAP7_75t_L g409 ( .A(n_255), .Y(n_409) );
AND2x2_ASAP7_75t_L g269 ( .A(n_256), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_256), .B(n_351), .Y(n_500) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g317 ( .A(n_257), .Y(n_317) );
INVx1_ASAP7_75t_L g393 ( .A(n_257), .Y(n_393) );
OR2x2_ASAP7_75t_L g446 ( .A(n_257), .B(n_315), .Y(n_446) );
INVx2_ASAP7_75t_L g277 ( .A(n_258), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_259), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_259), .B(n_360), .Y(n_381) );
INVx1_ASAP7_75t_L g441 ( .A(n_259), .Y(n_441) );
OAI31xp33_ASAP7_75t_L g497 ( .A1(n_259), .A2(n_413), .A3(n_498), .B(n_499), .Y(n_497) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_268), .Y(n_259) );
AND2x4_ASAP7_75t_L g288 ( .A(n_260), .B(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g363 ( .A(n_260), .B(n_283), .Y(n_363) );
INVx1_ASAP7_75t_L g398 ( .A(n_260), .Y(n_398) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g326 ( .A(n_261), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g306 ( .A(n_268), .Y(n_306) );
INVx1_ASAP7_75t_L g362 ( .A(n_268), .Y(n_362) );
OR2x2_ASAP7_75t_L g436 ( .A(n_268), .B(n_356), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_268), .B(n_302), .Y(n_494) );
AND2x4_ASAP7_75t_L g274 ( .A(n_270), .B(n_275), .Y(n_274) );
OAI221xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_280), .B1(n_286), .B2(n_291), .C(n_300), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_276), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g415 ( .A(n_276), .B(n_316), .Y(n_415) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
INVx1_ASAP7_75t_L g309 ( .A(n_278), .Y(n_309) );
INVx1_ASAP7_75t_L g367 ( .A(n_278), .Y(n_367) );
AND2x2_ASAP7_75t_L g431 ( .A(n_278), .B(n_352), .Y(n_431) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g294 ( .A(n_279), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
AND2x2_ASAP7_75t_L g336 ( .A(n_281), .B(n_326), .Y(n_336) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g323 ( .A(n_283), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_284), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g319 ( .A(n_285), .Y(n_319) );
AND2x4_ASAP7_75t_L g406 ( .A(n_285), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g485 ( .A(n_285), .B(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_287), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx2_ASAP7_75t_L g426 ( .A(n_288), .Y(n_426) );
INVx1_ASAP7_75t_L g342 ( .A(n_289), .Y(n_342) );
AND2x2_ASAP7_75t_L g325 ( .A(n_290), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g400 ( .A(n_290), .B(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_290), .Y(n_435) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_290), .Y(n_486) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_294), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_294), .B(n_350), .Y(n_481) );
INVx1_ASAP7_75t_L g374 ( .A(n_295), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g350 ( .A(n_299), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_304), .B(n_307), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x2_ASAP7_75t_L g451 ( .A(n_302), .B(n_363), .Y(n_451) );
AND2x2_ASAP7_75t_L g304 ( .A(n_303), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_SL g401 ( .A(n_303), .Y(n_401) );
INVx1_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g371 ( .A(n_309), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g428 ( .A(n_309), .B(n_373), .Y(n_428) );
OR2x2_ASAP7_75t_L g510 ( .A(n_310), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI32xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_318), .A3(n_320), .B1(n_324), .B2(n_328), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_314), .A2(n_419), .B1(n_451), .B2(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx2_ASAP7_75t_L g379 ( .A(n_315), .Y(n_379) );
NAND4xp25_ASAP7_75t_L g389 ( .A(n_315), .B(n_319), .C(n_390), .D(n_391), .Y(n_389) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g444 ( .A(n_316), .B(n_397), .Y(n_444) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g324 ( .A(n_321), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g504 ( .A(n_323), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_325), .A2(n_431), .B(n_459), .C(n_460), .Y(n_458) );
BUFx2_ASAP7_75t_L g413 ( .A(n_326), .Y(n_413) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_330), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g467 ( .A(n_330), .Y(n_467) );
INVx2_ASAP7_75t_L g404 ( .A(n_331), .Y(n_404) );
AND2x4_ASAP7_75t_L g460 ( .A(n_331), .B(n_372), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_337), .B(n_345), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
AOI322xp5_ASAP7_75t_L g438 ( .A1(n_339), .A2(n_439), .A3(n_441), .B1(n_442), .B2(n_443), .C1(n_445), .C2(n_447), .Y(n_438) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g457 ( .A(n_340), .B(n_344), .Y(n_457) );
INVx1_ASAP7_75t_L g468 ( .A(n_341), .Y(n_468) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AND2x2_ASAP7_75t_L g462 ( .A(n_342), .B(n_383), .Y(n_462) );
AND2x2_ASAP7_75t_L g483 ( .A(n_343), .B(n_362), .Y(n_483) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g493 ( .A(n_344), .B(n_494), .Y(n_493) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI222xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B1(n_357), .B2(n_361), .C1(n_364), .C2(n_953), .Y(n_348) );
NOR2x1_ASAP7_75t_L g370 ( .A(n_349), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx2_ASAP7_75t_L g391 ( .A(n_350), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_351), .B(n_421), .Y(n_440) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g425 ( .A(n_360), .B(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_360), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_361), .Y(n_490) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx3_ASAP7_75t_L g437 ( .A(n_363), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_364), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_375), .B(n_377), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_372), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g459 ( .A(n_372), .Y(n_459) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI32xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .A3(n_381), .B1(n_382), .B2(n_384), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g480 ( .A(n_379), .B(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g390 ( .A(n_383), .Y(n_390) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_463), .Y(n_386) );
NOR3xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_422), .C(n_449), .Y(n_387) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .C(n_405), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_391), .B(n_409), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_399), .B2(n_402), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B(n_411), .Y(n_405) );
INVx1_ASAP7_75t_L g448 ( .A(n_407), .Y(n_448) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g511 ( .A(n_410), .Y(n_511) );
OAI21xp33_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_414), .B(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g495 ( .A(n_415), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx2_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
AND2x2_ASAP7_75t_L g453 ( .A(n_421), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_438), .Y(n_422) );
AOI22xp5_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_427), .B1(n_429), .B2(n_432), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_426), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g466 ( .A(n_431), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2x1p5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .C(n_458), .D(n_461), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_460), .B(n_462), .Y(n_461) );
NOR4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_479), .C(n_487), .D(n_496), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_468), .B1(n_469), .B2(n_470), .C(n_471), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g476 ( .A(n_469), .Y(n_476) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g505 ( .A(n_473), .Y(n_505) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g508 ( .A(n_475), .Y(n_508) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI21xp5_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_482), .B(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B(n_491), .C(n_495), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI31xp33_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_505), .A3(n_506), .B(n_509), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_524), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_524), .B(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_SL g536 ( .A(n_526), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_532), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g923 ( .A(n_531), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_531), .B(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_920), .B(n_927), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_909), .B1(n_910), .B2(n_919), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_904), .B1(n_905), .B2(n_908), .Y(n_540) );
OA22x2_ASAP7_75t_L g919 ( .A1(n_541), .A2(n_904), .B1(n_905), .B2(n_908), .Y(n_919) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_773), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_701), .C(n_744), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_544), .B(n_670), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_609), .B(n_639), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_590), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_546), .A2(n_861), .B1(n_864), .B2(n_867), .Y(n_860) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_547), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_566), .Y(n_547) );
AND2x2_ASAP7_75t_L g650 ( .A(n_548), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g718 ( .A(n_548), .Y(n_718) );
AND2x2_ASAP7_75t_L g772 ( .A(n_548), .B(n_699), .Y(n_772) );
NAND2xp5_ASAP7_75t_SL g796 ( .A(n_548), .B(n_643), .Y(n_796) );
AND2x2_ASAP7_75t_L g834 ( .A(n_548), .B(n_696), .Y(n_834) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g682 ( .A(n_549), .Y(n_682) );
AND2x2_ASAP7_75t_L g780 ( .A(n_549), .B(n_680), .Y(n_780) );
INVx2_ASAP7_75t_L g866 ( .A(n_549), .Y(n_866) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g608 ( .A(n_550), .Y(n_608) );
AND2x2_ASAP7_75t_L g706 ( .A(n_550), .B(n_580), .Y(n_706) );
AOI21x1_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_554), .B(n_564), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND3x2_ASAP7_75t_L g865 ( .A(n_566), .B(n_593), .C(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g887 ( .A(n_566), .B(n_888), .Y(n_887) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_579), .Y(n_566) );
OR2x2_ASAP7_75t_L g679 ( .A(n_567), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g705 ( .A(n_567), .Y(n_705) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g696 ( .A(n_568), .Y(n_696) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_579), .Y(n_727) );
INVxp67_ASAP7_75t_L g754 ( .A(n_579), .Y(n_754) );
OR2x2_ASAP7_75t_L g766 ( .A(n_579), .B(n_595), .Y(n_766) );
OR2x2_ASAP7_75t_L g833 ( .A(n_579), .B(n_658), .Y(n_833) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g654 ( .A(n_580), .Y(n_654) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_582), .B(n_589), .Y(n_580) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g852 ( .A(n_591), .B(n_753), .Y(n_852) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_606), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g719 ( .A(n_593), .B(n_680), .Y(n_719) );
AND2x2_ASAP7_75t_L g779 ( .A(n_593), .B(n_705), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g876 ( .A(n_593), .B(n_866), .Y(n_876) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g652 ( .A(n_594), .B(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g801 ( .A(n_594), .Y(n_801) );
NAND2x1_ASAP7_75t_L g814 ( .A(n_594), .B(n_795), .Y(n_814) );
AND2x2_ASAP7_75t_L g888 ( .A(n_594), .B(n_866), .Y(n_888) );
INVx4_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g677 ( .A(n_595), .Y(n_677) );
INVx1_ASAP7_75t_L g694 ( .A(n_595), .Y(n_694) );
AND2x2_ASAP7_75t_L g699 ( .A(n_595), .B(n_696), .Y(n_699) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_601), .B(n_605), .Y(n_597) );
AND2x2_ASAP7_75t_L g805 ( .A(n_606), .B(n_677), .Y(n_805) );
INVx1_ASAP7_75t_L g812 ( .A(n_606), .Y(n_812) );
AND2x2_ASAP7_75t_L g838 ( .A(n_606), .B(n_693), .Y(n_838) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g695 ( .A(n_608), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_622), .Y(n_610) );
INVx2_ASAP7_75t_L g786 ( .A(n_611), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_611), .B(n_643), .Y(n_868) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g647 ( .A(n_612), .Y(n_647) );
AND2x2_ASAP7_75t_L g685 ( .A(n_612), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g714 ( .A(n_612), .B(n_644), .Y(n_714) );
AND2x2_ASAP7_75t_L g764 ( .A(n_612), .B(n_632), .Y(n_764) );
AND2x2_ASAP7_75t_L g882 ( .A(n_612), .B(n_659), .Y(n_882) );
AND2x2_ASAP7_75t_L g721 ( .A(n_622), .B(n_697), .Y(n_721) );
BUFx2_ASAP7_75t_L g788 ( .A(n_622), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_622), .B(n_750), .Y(n_815) );
INVx1_ASAP7_75t_L g900 ( .A(n_622), .Y(n_900) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_632), .Y(n_622) );
AND2x2_ASAP7_75t_L g669 ( .A(n_623), .B(n_648), .Y(n_669) );
OR2x2_ASAP7_75t_L g712 ( .A(n_623), .B(n_632), .Y(n_712) );
INVx1_ASAP7_75t_L g739 ( .A(n_623), .Y(n_739) );
INVx1_ASAP7_75t_L g648 ( .A(n_632), .Y(n_648) );
AND2x2_ASAP7_75t_L g673 ( .A(n_632), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_632), .B(n_690), .Y(n_689) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_632), .Y(n_725) );
OR2x2_ASAP7_75t_L g741 ( .A(n_632), .B(n_690), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_649), .B(n_655), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2x1p5_ASAP7_75t_L g730 ( .A(n_641), .B(n_731), .Y(n_730) );
NAND2x1_ASAP7_75t_L g857 ( .A(n_641), .B(n_732), .Y(n_857) );
AND2x4_ASAP7_75t_L g641 ( .A(n_642), .B(n_646), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_642), .B(n_844), .Y(n_863) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g825 ( .A(n_644), .B(n_647), .Y(n_825) );
BUFx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g674 ( .A(n_645), .Y(n_674) );
AND2x2_ASAP7_75t_L g839 ( .A(n_646), .B(n_691), .Y(n_839) );
AND2x4_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g810 ( .A(n_652), .Y(n_810) );
OR2x2_ASAP7_75t_L g818 ( .A(n_652), .B(n_812), .Y(n_818) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g680 ( .A(n_654), .Y(n_680) );
AND2x2_ASAP7_75t_L g693 ( .A(n_654), .B(n_694), .Y(n_693) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_654), .Y(n_700) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_669), .Y(n_656) );
AND2x2_ASAP7_75t_L g756 ( .A(n_657), .B(n_693), .Y(n_756) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g769 ( .A(n_659), .B(n_690), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_669), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g845 ( .A(n_669), .Y(n_845) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_669), .B(n_862), .Y(n_861) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B1(n_683), .B2(n_692), .C1(n_697), .C2(n_698), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_672), .B(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g808 ( .A(n_673), .B(n_691), .Y(n_808) );
AND2x2_ASAP7_75t_L g856 ( .A(n_673), .B(n_769), .Y(n_856) );
AND2x2_ASAP7_75t_L g892 ( .A(n_673), .B(n_697), .Y(n_892) );
BUFx2_ASAP7_75t_L g771 ( .A(n_674), .Y(n_771) );
AND2x4_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x4_ASAP7_75t_L g703 ( .A(n_677), .B(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_677), .B(n_786), .Y(n_793) );
OR3x2_ASAP7_75t_L g846 ( .A(n_677), .B(n_679), .C(n_681), .Y(n_846) );
NOR2x1p5_ASAP7_75t_SL g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g743 ( .A(n_679), .Y(n_743) );
AND2x2_ASAP7_75t_L g873 ( .A(n_680), .B(n_695), .Y(n_873) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_688), .Y(n_683) );
INVx1_ASAP7_75t_L g895 ( .A(n_684), .Y(n_895) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g723 ( .A(n_685), .B(n_724), .Y(n_723) );
BUFx3_ASAP7_75t_L g691 ( .A(n_686), .Y(n_691) );
AND2x2_ASAP7_75t_L g697 ( .A(n_686), .B(n_690), .Y(n_697) );
INVxp67_ASAP7_75t_SL g733 ( .A(n_686), .Y(n_733) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_686), .Y(n_735) );
INVx1_ASAP7_75t_L g751 ( .A(n_686), .Y(n_751) );
INVx1_ASAP7_75t_L g844 ( .A(n_686), .Y(n_844) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_688), .B(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g830 ( .A(n_689), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_691), .B(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g869 ( .A(n_691), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_691), .B(n_764), .Y(n_877) );
NAND2xp5_ASAP7_75t_SL g884 ( .A(n_691), .B(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
AND2x2_ASAP7_75t_L g897 ( .A(n_693), .B(n_718), .Y(n_897) );
INVx2_ASAP7_75t_L g760 ( .A(n_695), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_695), .B(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g795 ( .A(n_696), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_697), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g728 ( .A(n_699), .Y(n_728) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_699), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_699), .B(n_780), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_729), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_707), .B(n_715), .Y(n_702) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g880 ( .A(n_705), .Y(n_880) );
INVx2_ASAP7_75t_L g784 ( .A(n_706), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_706), .B(n_801), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_713), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_711), .B(n_832), .C(n_834), .Y(n_831) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g804 ( .A(n_712), .B(n_750), .Y(n_804) );
INVx1_ASAP7_75t_L g885 ( .A(n_712), .Y(n_885) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x4_ASAP7_75t_L g851 ( .A(n_714), .B(n_735), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_720), .B1(n_722), .B2(n_726), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_723), .B(n_799), .Y(n_836) );
INVx1_ASAP7_75t_L g792 ( .A(n_724), .Y(n_792) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g797 ( .A(n_727), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_727), .B(n_880), .Y(n_879) );
NOR2x1_ASAP7_75t_SL g783 ( .A(n_728), .B(n_784), .Y(n_783) );
AO21x1_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_734), .B(n_742), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g763 ( .A(n_733), .B(n_764), .Y(n_763) );
NAND2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_736), .B(n_799), .Y(n_798) );
AND2x4_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_738), .Y(n_758) );
AND2x2_ASAP7_75t_L g855 ( .A(n_738), .B(n_764), .Y(n_855) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g822 ( .A(n_741), .Y(n_822) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_759), .B(n_761), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_755), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_750), .B(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
BUFx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OR2x2_ASAP7_75t_L g765 ( .A(n_760), .B(n_766), .Y(n_765) );
OAI21xp33_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_765), .B(n_767), .Y(n_761) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_772), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g781 ( .A(n_769), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_769), .B(n_770), .Y(n_871) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NOR2x1_ASAP7_75t_L g773 ( .A(n_774), .B(n_847), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_816), .Y(n_774) );
AOI211xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_787), .B(n_789), .C(n_806), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_781), .B1(n_782), .B2(n_785), .Y(n_776) );
INVx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x4_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
AND2x2_ASAP7_75t_L g893 ( .A(n_780), .B(n_801), .Y(n_893) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
OR2x6_ASAP7_75t_L g813 ( .A(n_784), .B(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND3xp33_ASAP7_75t_L g878 ( .A(n_788), .B(n_879), .C(n_881), .Y(n_878) );
NAND3xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_798), .C(n_802), .Y(n_789) );
NAND4xp25_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .C(n_794), .D(n_797), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx1_ASAP7_75t_SL g875 ( .A(n_795), .Y(n_875) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
OAI22xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_809), .B1(n_813), .B2(n_815), .Y(n_806) );
INVx3_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_808), .B(n_851), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g894 ( .A(n_813), .Y(n_894) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_835), .C(n_840), .Y(n_816) );
OAI211xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B(n_826), .C(n_831), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_823), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_846), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_845), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g903 ( .A(n_845), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g847 ( .A(n_848), .B(n_859), .C(n_890), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_853), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_850), .B(n_852), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_857), .B(n_858), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
INVx2_ASAP7_75t_L g889 ( .A(n_855), .Y(n_889) );
NOR3xp33_ASAP7_75t_SL g859 ( .A(n_860), .B(n_870), .C(n_883), .Y(n_859) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OR2x2_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
OAI221xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_874), .B2(n_877), .C(n_878), .Y(n_870) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g883 ( .A1(n_874), .A2(n_884), .B1(n_886), .B2(n_889), .Y(n_883) );
OR2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
BUFx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NAND2x1_ASAP7_75t_L g899 ( .A(n_882), .B(n_900), .Y(n_899) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_896), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_893), .B1(n_894), .B2(n_895), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_898), .B1(n_901), .B2(n_903), .Y(n_896) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx3_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
BUFx8_ASAP7_75t_SL g905 ( .A(n_906), .Y(n_905) );
AND2x2_ASAP7_75t_L g934 ( .A(n_906), .B(n_935), .Y(n_934) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
BUFx2_ASAP7_75t_L g949 ( .A(n_907), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx3_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx6_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AND2x6_ASAP7_75t_SL g922 ( .A(n_923), .B(n_924), .Y(n_922) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
BUFx6f_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
BUFx10_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
BUFx6f_ASAP7_75t_L g951 ( .A(n_936), .Y(n_951) );
INVx8_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
OR2x6_ASAP7_75t_L g937 ( .A(n_938), .B(n_943), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .Y(n_939) );
INVxp33_ASAP7_75t_SL g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
NOR3xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_948), .C(n_949), .Y(n_944) );
INVx2_ASAP7_75t_SL g945 ( .A(n_946), .Y(n_945) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
endmodule