module fake_jpeg_13919_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_0),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_20),
.C(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_4),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_23),
.B1(n_19),
.B2(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_36),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_20),
.B(n_17),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.C(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_31),
.B1(n_11),
.B2(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.C(n_33),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_8),
.B1(n_7),
.B2(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_34),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_44),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_38),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_27),
.C(n_32),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_4),
.C(n_5),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_42),
.B(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_6),
.B(n_45),
.C(n_46),
.Y(n_50)
);


endmodule