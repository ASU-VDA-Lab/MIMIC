module fake_netlist_1_8333_n_375 (n_107, n_103, n_52, n_50, n_7, n_3, n_34, n_25, n_9, n_96, n_72, n_77, n_90, n_99, n_43, n_73, n_62, n_97, n_33, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_66, n_88, n_46, n_108, n_37, n_18, n_65, n_87, n_5, n_81, n_85, n_102, n_47, n_109, n_1, n_16, n_78, n_95, n_40, n_68, n_105, n_36, n_11, n_15, n_71, n_70, n_94, n_2, n_17, n_58, n_20, n_84, n_12, n_56, n_80, n_67, n_22, n_19, n_26, n_39, n_101, n_98, n_38, n_104, n_100, n_24, n_35, n_91, n_32, n_93, n_48, n_63, n_54, n_41, n_55, n_29, n_60, n_10, n_30, n_13, n_92, n_75, n_82, n_53, n_64, n_69, n_83, n_23, n_0, n_57, n_51, n_106, n_45, n_42, n_21, n_86, n_27, n_89, n_28, n_79, n_49, n_14, n_31, n_375, n_948);
input n_107;
input n_103;
input n_52;
input n_50;
input n_7;
input n_3;
input n_34;
input n_25;
input n_9;
input n_96;
input n_72;
input n_77;
input n_90;
input n_99;
input n_43;
input n_73;
input n_62;
input n_97;
input n_33;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_66;
input n_88;
input n_46;
input n_108;
input n_37;
input n_18;
input n_65;
input n_87;
input n_5;
input n_81;
input n_85;
input n_102;
input n_47;
input n_109;
input n_1;
input n_16;
input n_78;
input n_95;
input n_40;
input n_68;
input n_105;
input n_36;
input n_11;
input n_15;
input n_71;
input n_70;
input n_94;
input n_2;
input n_17;
input n_58;
input n_20;
input n_84;
input n_12;
input n_56;
input n_80;
input n_67;
input n_22;
input n_19;
input n_26;
input n_39;
input n_101;
input n_98;
input n_38;
input n_104;
input n_100;
input n_24;
input n_35;
input n_91;
input n_32;
input n_93;
input n_48;
input n_63;
input n_54;
input n_41;
input n_55;
input n_29;
input n_60;
input n_10;
input n_30;
input n_13;
input n_92;
input n_75;
input n_82;
input n_53;
input n_64;
input n_69;
input n_83;
input n_23;
input n_0;
input n_57;
input n_51;
input n_106;
input n_45;
input n_42;
input n_21;
input n_86;
input n_27;
input n_89;
input n_28;
input n_79;
input n_49;
input n_14;
input n_31;
output n_375;
output n_948;
wire n_890;
wire n_646;
wire n_107;
wire n_759;
wire n_658;
wire n_673;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_944;
wire n_356;
wire n_895;
wire n_327;
wire n_25;
wire n_204;
wire n_592;
wire n_769;
wire n_929;
wire n_169;
wire n_370;
wire n_384;
wire n_439;
wire n_545;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_786;
wire n_831;
wire n_357;
wire n_74;
wire n_729;
wire n_308;
wire n_518;
wire n_394;
wire n_44;
wire n_189;
wire n_681;
wire n_226;
wire n_352;
wire n_447;
wire n_66;
wire n_379;
wire n_903;
wire n_535;
wire n_689;
wire n_886;
wire n_595;
wire n_875;
wire n_626;
wire n_316;
wire n_285;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_766;
wire n_475;
wire n_744;
wire n_850;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_942;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_805;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_557;
wire n_288;
wire n_176;
wire n_753;
wire n_859;
wire n_438;
wire n_900;
wire n_869;
wire n_931;
wire n_935;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_723;
wire n_223;
wire n_833;
wire n_405;
wire n_830;
wire n_562;
wire n_19;
wire n_409;
wire n_482;
wire n_838;
wire n_534;
wire n_569;
wire n_707;
wire n_526;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_709;
wire n_303;
wire n_502;
wire n_821;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_301;
wire n_340;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_752;
wire n_246;
wire n_676;
wire n_823;
wire n_191;
wire n_143;
wire n_780;
wire n_864;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_876;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_494;
wire n_553;
wire n_343;
wire n_555;
wire n_135;
wire n_481;
wire n_621;
wire n_817;
wire n_776;
wire n_315;
wire n_397;
wire n_53;
wire n_880;
wire n_213;
wire n_196;
wire n_293;
wire n_797;
wire n_836;
wire n_127;
wire n_312;
wire n_742;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_751;
wire n_887;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_164;
wire n_433;
wire n_660;
wire n_120;
wire n_392;
wire n_650;
wire n_806;
wire n_155;
wire n_162;
wire n_114;
wire n_772;
wire n_50;
wire n_816;
wire n_789;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_882;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_884;
wire n_9;
wire n_737;
wire n_428;
wire n_178;
wire n_478;
wire n_814;
wire n_652;
wire n_678;
wire n_708;
wire n_229;
wire n_97;
wire n_133;
wire n_442;
wire n_324;
wire n_422;
wire n_192;
wire n_699;
wire n_857;
wire n_329;
wire n_6;
wire n_8;
wire n_578;
wire n_928;
wire n_883;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_801;
wire n_441;
wire n_868;
wire n_628;
wire n_425;
wire n_912;
wire n_920;
wire n_314;
wire n_824;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_736;
wire n_172;
wire n_905;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_934;
wire n_653;
wire n_351;
wire n_1;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_755;
wire n_716;
wire n_228;
wire n_863;
wire n_671;
wire n_892;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_765;
wire n_829;
wire n_599;
wire n_715;
wire n_849;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_721;
wire n_362;
wire n_617;
wire n_688;
wire n_837;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_720;
wire n_152;
wire n_851;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_855;
wire n_17;
wire n_322;
wire n_911;
wire n_506;
wire n_221;
wire n_328;
wire n_317;
wire n_711;
wire n_491;
wire n_800;
wire n_388;
wire n_773;
wire n_266;
wire n_763;
wire n_80;
wire n_632;
wire n_793;
wire n_906;
wire n_679;
wire n_522;
wire n_546;
wire n_615;
wire n_684;
wire n_701;
wire n_532;
wire n_326;
wire n_756;
wire n_635;
wire n_544;
wire n_888;
wire n_879;
wire n_576;
wire n_275;
wire n_691;
wire n_622;
wire n_661;
wire n_909;
wire n_493;
wire n_274;
wire n_910;
wire n_150;
wire n_235;
wire n_690;
wire n_38;
wire n_533;
wire n_272;
wire n_686;
wire n_299;
wire n_100;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_757;
wire n_844;
wire n_695;
wire n_193;
wire n_344;
wire n_232;
wire n_878;
wire n_812;
wire n_783;
wire n_147;
wire n_185;
wire n_367;
wire n_795;
wire n_267;
wire n_687;
wire n_171;
wire n_638;
wire n_873;
wire n_899;
wire n_450;
wire n_585;
wire n_140;
wire n_644;
wire n_111;
wire n_779;
wire n_212;
wire n_746;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_704;
wire n_435;
wire n_728;
wire n_583;
wire n_841;
wire n_64;
wire n_69;
wire n_248;
wire n_866;
wire n_407;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_262;
wire n_921;
wire n_119;
wire n_667;
wire n_503;
wire n_856;
wire n_927;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_748;
wire n_79;
wire n_129;
wire n_904;
wire n_611;
wire n_521;
wire n_157;
wire n_774;
wire n_103;
wire n_808;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_273;
wire n_325;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_743;
wire n_163;
wire n_348;
wire n_96;
wire n_669;
wire n_685;
wire n_72;
wire n_77;
wire n_90;
wire n_594;
wire n_762;
wire n_214;
wire n_787;
wire n_740;
wire n_770;
wire n_167;
wire n_861;
wire n_809;
wire n_364;
wire n_33;
wire n_908;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_609;
wire n_946;
wire n_121;
wire n_286;
wire n_206;
wire n_408;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_860;
wire n_413;
wire n_537;
wire n_65;
wire n_710;
wire n_525;
wire n_560;
wire n_5;
wire n_496;
wire n_393;
wire n_843;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_733;
wire n_846;
wire n_290;
wire n_217;
wire n_201;
wire n_791;
wire n_792;
wire n_277;
wire n_932;
wire n_259;
wire n_885;
wire n_612;
wire n_244;
wire n_666;
wire n_771;
wire n_827;
wire n_276;
wire n_297;
wire n_225;
wire n_631;
wire n_350;
wire n_747;
wire n_208;
wire n_616;
wire n_815;
wire n_523;
wire n_854;
wire n_901;
wire n_528;
wire n_419;
wire n_252;
wire n_922;
wire n_519;
wire n_168;
wire n_839;
wire n_271;
wire n_693;
wire n_785;
wire n_896;
wire n_739;
wire n_94;
wire n_194;
wire n_858;
wire n_758;
wire n_825;
wire n_282;
wire n_58;
wire n_775;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_321;
wire n_302;
wire n_538;
wire n_703;
wire n_811;
wire n_116;
wire n_734;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_597;
wire n_554;
wire n_698;
wire n_705;
wire n_257;
wire n_741;
wire n_828;
wire n_722;
wire n_26;
wire n_203;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_714;
wire n_146;
wire n_337;
wire n_32;
wire n_637;
wire n_641;
wire n_726;
wire n_531;
wire n_872;
wire n_539;
wire n_93;
wire n_847;
wire n_406;
wire n_372;
wire n_842;
wire n_820;
wire n_713;
wire n_467;
wire n_923;
wire n_702;
wire n_41;
wire n_760;
wire n_826;
wire n_918;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_898;
wire n_647;
wire n_445;
wire n_500;
wire n_732;
wire n_926;
wire n_845;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_818;
wire n_82;
wire n_75;
wire n_183;
wire n_731;
wire n_550;
wire n_132;
wire n_643;
wire n_761;
wire n_778;
wire n_582;
wire n_784;
wire n_170;
wire n_925;
wire n_205;
wire n_158;
wire n_915;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_834;
wire n_510;
wire n_360;
wire n_363;
wire n_749;
wire n_427;
wire n_724;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_835;
wire n_437;
wire n_871;
wire n_620;
wire n_89;
wire n_480;
wire n_939;
wire n_940;
wire n_130;
wire n_310;
wire n_341;
wire n_700;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_727;
wire n_136;
wire n_260;
wire n_891;
wire n_580;
wire n_610;
wire n_938;
wire n_222;
wire n_657;
wire n_822;
wire n_381;
wire n_142;
wire n_34;
wire n_853;
wire n_754;
wire n_385;
wire n_798;
wire n_395;
wire n_227;
wire n_454;
wire n_943;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_190;
wire n_606;
wire n_62;
wire n_712;
wire n_777;
wire n_4;
wire n_565;
wire n_323;
wire n_59;
wire n_781;
wire n_914;
wire n_945;
wire n_852;
wire n_376;
wire n_902;
wire n_694;
wire n_240;
wire n_459;
wire n_768;
wire n_568;
wire n_88;
wire n_46;
wire n_174;
wire n_717;
wire n_807;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_802;
wire n_865;
wire n_672;
wire n_867;
wire n_87;
wire n_466;
wire n_349;
wire n_207;
wire n_197;
wire n_541;
wire n_572;
wire n_81;
wire n_298;
wire n_112;
wire n_630;
wire n_735;
wire n_649;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_919;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_810;
wire n_36;
wire n_416;
wire n_916;
wire n_870;
wire n_889;
wire n_432;
wire n_913;
wire n_917;
wire n_465;
wire n_414;
wire n_730;
wire n_680;
wire n_369;
wire n_469;
wire n_361;
wire n_767;
wire n_237;
wire n_881;
wire n_654;
wire n_15;
wire n_520;
wire n_633;
wire n_429;
wire n_803;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_804;
wire n_796;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_907;
wire n_591;
wire n_391;
wire n_209;
wire n_241;
wire n_874;
wire n_84;
wire n_20;
wire n_782;
wire n_449;
wire n_832;
wire n_12;
wire n_412;
wire n_56;
wire n_455;
wire n_67;
wire n_504;
wire n_618;
wire n_790;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_877;
wire n_383;
wire n_813;
wire n_202;
wire n_319;
wire n_542;
wire n_725;
wire n_819;
wire n_862;
wire n_930;
wire n_39;
wire n_101;
wire n_941;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_933;
wire n_508;
wire n_764;
wire n_719;
wire n_486;
wire n_788;
wire n_24;
wire n_35;
wire n_655;
wire n_472;
wire n_490;
wire n_540;
wire n_947;
wire n_840;
wire n_400;
wire n_794;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_563;
wire n_513;
wire n_55;
wire n_718;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_893;
wire n_173;
wire n_488;
wire n_556;
wire n_648;
wire n_382;
wire n_799;
wire n_894;
wire n_138;
wire n_60;
wire n_936;
wire n_937;
wire n_462;
wire n_536;
wire n_573;
wire n_474;
wire n_924;
wire n_745;
wire n_305;
wire n_505;
wire n_430;
wire n_418;
wire n_495;
wire n_358;
wire n_313;
wire n_333;
wire n_627;
wire n_92;
wire n_706;
wire n_750;
wire n_589;
wire n_175;
wire n_897;
wire n_128;
wire n_306;
wire n_31;
wire n_697;
wire n_0;
wire n_512;
wire n_258;
wire n_619;
wire n_642;
wire n_675;
wire n_607;
wire n_234;
wire n_848;
wire n_184;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_144;
wire n_403;
wire n_625;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_738;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_436;
wire n_415;
INVx1_ASAP7_75t_L g110 ( .A(n_48), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_84), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_45), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_69), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_49), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_94), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_97), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_15), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_1), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_96), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_87), .Y(n_120) );
BUFx8_ASAP7_75t_SL g121 ( .A(n_46), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_64), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_22), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_68), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_71), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_99), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_58), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_7), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_74), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_40), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_103), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g132 ( .A(n_105), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_8), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_80), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_6), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_104), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_85), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_9), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_29), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_76), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_21), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_82), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_108), .Y(n_143) );
BUFx10_ASAP7_75t_L g144 ( .A(n_7), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_36), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_102), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_39), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_86), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_32), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_38), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_109), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_13), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_23), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_37), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_67), .Y(n_155) );
NOR2xp33_ASAP7_75t_SL g156 ( .A(n_134), .B(n_42), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_127), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_110), .B(n_112), .Y(n_159) );
INVx5_ASAP7_75t_L g160 ( .A(n_127), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_110), .B(n_0), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_112), .B(n_0), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_137), .B(n_1), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_143), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_117), .B(n_2), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_117), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_128), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_121), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_133), .B(n_138), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_111), .B(n_2), .Y(n_178) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_175), .A2(n_123), .B1(n_141), .B2(n_152), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_178), .A2(n_111), .B1(n_132), .B2(n_153), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_163), .A2(n_154), .B1(n_139), .B2(n_147), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_175), .A2(n_123), .B1(n_135), .B2(n_154), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_178), .A2(n_132), .B1(n_118), .B2(n_150), .Y(n_183) );
NAND3x1_ASAP7_75t_L g184 ( .A(n_178), .B(n_139), .C(n_145), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_175), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_163), .A2(n_145), .B1(n_147), .B2(n_134), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_175), .B(n_144), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_170), .A2(n_130), .B1(n_149), .B2(n_126), .Y(n_189) );
OAI22xp33_ASAP7_75t_SL g190 ( .A1(n_170), .A2(n_144), .B1(n_155), .B2(n_148), .Y(n_190) );
BUFx10_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_162), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
OA22x2_ASAP7_75t_L g196 ( .A1(n_163), .A2(n_124), .B1(n_114), .B2(n_142), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_170), .A2(n_151), .B1(n_113), .B2(n_140), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_162), .B(n_115), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
AO22x2_ASAP7_75t_L g201 ( .A1(n_165), .A2(n_144), .B1(n_121), .B2(n_5), .Y(n_201) );
OAI22xp33_ASAP7_75t_SL g202 ( .A1(n_159), .A2(n_136), .B1(n_131), .B2(n_129), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_178), .A2(n_125), .B1(n_122), .B2(n_120), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_176), .B(n_171), .Y(n_204) );
AO22x2_ASAP7_75t_L g205 ( .A1(n_165), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_205) );
AO22x2_ASAP7_75t_L g206 ( .A1(n_165), .A2(n_3), .B1(n_4), .B2(n_6), .Y(n_206) );
AO22x2_ASAP7_75t_L g207 ( .A1(n_165), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g208 ( .A1(n_171), .A2(n_119), .B1(n_116), .B2(n_12), .Y(n_208) );
CKINVDCx6p67_ASAP7_75t_R g209 ( .A(n_162), .Y(n_209) );
OAI22xp33_ASAP7_75t_R g210 ( .A1(n_176), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_165), .A2(n_11), .B1(n_13), .B2(n_14), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g212 ( .A1(n_171), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_213) );
OR2x6_ASAP7_75t_L g214 ( .A(n_165), .B(n_17), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_174), .Y(n_217) );
OAI22xp33_ASAP7_75t_SL g218 ( .A1(n_159), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_218) );
AO22x2_ASAP7_75t_L g219 ( .A1(n_174), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_156), .B(n_22), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_174), .A2(n_23), .B1(n_24), .B2(n_25), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_162), .A2(n_24), .B1(n_25), .B2(n_26), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_214), .B(n_162), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_204), .B(n_162), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_195), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_195), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_187), .B(n_162), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_197), .Y(n_231) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_215), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_185), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_197), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_188), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_192), .Y(n_236) );
XOR2xp5_ASAP7_75t_L g237 ( .A(n_179), .B(n_26), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_217), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_181), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_181), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_181), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_191), .Y(n_242) );
XOR2xp5_ASAP7_75t_L g243 ( .A(n_179), .B(n_27), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_185), .B(n_162), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_191), .Y(n_245) );
INVx3_ASAP7_75t_R g246 ( .A(n_199), .Y(n_246) );
XOR2xp5_ASAP7_75t_L g247 ( .A(n_201), .B(n_27), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_186), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_180), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_198), .B(n_162), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_182), .B(n_176), .Y(n_251) );
INVxp67_ASAP7_75t_L g252 ( .A(n_201), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_214), .B(n_161), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_186), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_186), .B(n_161), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_214), .B(n_161), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_198), .B(n_199), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_182), .B(n_167), .Y(n_258) );
XNOR2xp5_ASAP7_75t_L g259 ( .A(n_201), .B(n_28), .Y(n_259) );
INVxp33_ASAP7_75t_SL g260 ( .A(n_183), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_203), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_190), .B(n_202), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_194), .B(n_167), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_205), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_209), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_196), .B(n_167), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_206), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_222), .B(n_167), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_216), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_196), .B(n_189), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_206), .Y(n_274) );
XOR2xp5_ASAP7_75t_L g275 ( .A(n_189), .B(n_28), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_193), .Y(n_276) );
NOR2xp33_ASAP7_75t_SL g277 ( .A(n_222), .B(n_156), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_220), .B(n_167), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_200), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_207), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_211), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_213), .Y(n_283) );
NOR2xp67_ASAP7_75t_L g284 ( .A(n_225), .B(n_167), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_207), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_207), .B(n_167), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_221), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_223), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_219), .B(n_169), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_220), .A2(n_169), .B(n_158), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_219), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_271), .B(n_184), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_238), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_271), .B(n_219), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_227), .B(n_169), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_226), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_227), .B(n_169), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_289), .B(n_169), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_238), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_253), .B(n_169), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_289), .B(n_169), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_226), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_226), .B(n_224), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_226), .B(n_224), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_258), .B(n_160), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_258), .B(n_160), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_235), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_268), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_235), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_253), .B(n_208), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_235), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_253), .B(n_208), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_253), .B(n_212), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_268), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_233), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_256), .B(n_212), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_276), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_239), .B(n_160), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_256), .B(n_218), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_268), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_228), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_236), .B(n_164), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_244), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_286), .B(n_160), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_239), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_286), .B(n_160), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_236), .B(n_164), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_273), .B(n_164), .Y(n_328) );
AND2x6_ASAP7_75t_L g329 ( .A(n_240), .B(n_164), .Y(n_329) );
INVxp33_ASAP7_75t_L g330 ( .A(n_263), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_257), .B(n_156), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_255), .B(n_164), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_228), .Y(n_333) );
INVx11_ASAP7_75t_L g334 ( .A(n_246), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_255), .B(n_164), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_240), .B(n_160), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_230), .B(n_164), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_267), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_251), .B(n_247), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_241), .B(n_160), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_257), .B(n_164), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_276), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_241), .B(n_160), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_274), .B(n_160), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_267), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_246), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_284), .B(n_269), .Y(n_347) );
OR2x6_ASAP7_75t_SL g348 ( .A(n_339), .B(n_291), .Y(n_348) );
NOR2x1_ASAP7_75t_L g349 ( .A(n_338), .B(n_291), .Y(n_349) );
NOR2x1p5_ASAP7_75t_L g350 ( .A(n_296), .B(n_262), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_293), .B(n_251), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_293), .Y(n_352) );
OR2x6_ASAP7_75t_L g353 ( .A(n_303), .B(n_274), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_293), .B(n_262), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_296), .B(n_252), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_299), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_307), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_299), .B(n_264), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_303), .B(n_230), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_315), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_307), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_299), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_315), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_307), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_302), .Y(n_366) );
BUFx2_ASAP7_75t_SL g367 ( .A(n_302), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_339), .B(n_247), .Y(n_368) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_302), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_315), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_310), .B(n_260), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_302), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_300), .B(n_242), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_334), .Y(n_374) );
UNKNOWN g375 ( );
AND2x4_ASAP7_75t_L g376 ( .A(n_300), .B(n_242), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_303), .B(n_244), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_303), .B(n_285), .Y(n_378) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_329), .B(n_277), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_308), .B(n_277), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_321), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_302), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_357), .Y(n_383) );
INVx6_ASAP7_75t_L g384 ( .A(n_369), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_357), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_352), .B(n_294), .Y(n_386) );
INVx4_ASAP7_75t_L g387 ( .A(n_358), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_364), .Y(n_388) );
INVx4_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_357), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_369), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_357), .Y(n_392) );
INVx5_ASAP7_75t_L g393 ( .A(n_369), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
INVx4_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_369), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_358), .Y(n_398) );
INVx8_ASAP7_75t_L g399 ( .A(n_353), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_377), .B(n_304), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_358), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_362), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_358), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_358), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_362), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_365), .Y(n_406) );
BUFx12f_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
BUFx3_ASAP7_75t_L g409 ( .A(n_358), .Y(n_409) );
INVx2_ASAP7_75t_SL g410 ( .A(n_365), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_365), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_377), .B(n_304), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_358), .Y(n_413) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_388), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_397), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_392), .Y(n_416) );
INVx4_ASAP7_75t_L g417 ( .A(n_393), .Y(n_417) );
BUFx2_ASAP7_75t_SL g418 ( .A(n_393), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_407), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_392), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_392), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_399), .A2(n_353), .B1(n_259), .B2(n_339), .Y(n_422) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_393), .A2(n_368), .B1(n_339), .B2(n_353), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_393), .A2(n_368), .B1(n_353), .B2(n_364), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_400), .B(n_371), .Y(n_426) );
BUFx4f_ASAP7_75t_SL g427 ( .A(n_391), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_399), .A2(n_371), .B1(n_259), .B2(n_368), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_388), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_400), .B(n_316), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_399), .A2(n_210), .B1(n_353), .B2(n_330), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_393), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_397), .Y(n_433) );
INVx8_ASAP7_75t_L g434 ( .A(n_393), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_383), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_399), .A2(n_353), .B1(n_243), .B2(n_237), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_393), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_393), .A2(n_353), .B1(n_313), .B2(n_348), .Y(n_438) );
INVx6_ASAP7_75t_L g439 ( .A(n_393), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_405), .Y(n_440) );
INVx6_ASAP7_75t_L g441 ( .A(n_393), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_383), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g443 ( .A1(n_399), .A2(n_370), .B1(n_361), .B2(n_294), .Y(n_443) );
AOI22xp33_ASAP7_75t_SL g444 ( .A1(n_399), .A2(n_370), .B1(n_361), .B2(n_294), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_383), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_393), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_383), .Y(n_447) );
BUFx4_ASAP7_75t_R g448 ( .A(n_393), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_391), .A2(n_283), .B1(n_282), .B2(n_249), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_385), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_385), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_392), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_393), .Y(n_453) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_399), .A2(n_313), .B1(n_348), .B2(n_312), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g455 ( .A1(n_399), .A2(n_294), .B1(n_304), .B2(n_379), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_407), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_400), .A2(n_275), .B1(n_237), .B2(n_243), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_399), .A2(n_304), .B1(n_275), .B2(n_377), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_426), .B(n_400), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_422), .A2(n_399), .B1(n_384), .B2(n_391), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_449), .B(n_261), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_414), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_431), .A2(n_412), .B1(n_400), .B2(n_360), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_423), .A2(n_412), .B1(n_360), .B2(n_384), .Y(n_464) );
OAI21xp5_ASAP7_75t_SL g465 ( .A1(n_457), .A2(n_396), .B(n_391), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_416), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_424), .A2(n_412), .B1(n_360), .B2(n_384), .Y(n_467) );
OAI21xp5_ASAP7_75t_SL g468 ( .A1(n_457), .A2(n_396), .B(n_391), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_428), .A2(n_310), .B1(n_312), .B2(n_316), .C1(n_313), .C2(n_375), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_430), .B(n_412), .Y(n_470) );
OAI21xp5_ASAP7_75t_SL g471 ( .A1(n_436), .A2(n_396), .B(n_316), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_448), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_417), .B(n_385), .Y(n_475) );
OAI21xp5_ASAP7_75t_SL g476 ( .A1(n_438), .A2(n_396), .B(n_266), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_435), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_454), .A2(n_284), .B(n_331), .Y(n_478) );
OAI222xp33_ASAP7_75t_L g479 ( .A1(n_417), .A2(n_396), .B1(n_387), .B2(n_389), .C1(n_395), .C2(n_403), .Y(n_479) );
OAI22xp33_ASAP7_75t_L g480 ( .A1(n_427), .A2(n_419), .B1(n_417), .B2(n_434), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_416), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_442), .B(n_385), .Y(n_482) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_418), .A2(n_384), .B1(n_396), .B2(n_395), .Y(n_483) );
NOR2x1_ASAP7_75t_R g484 ( .A(n_414), .B(n_407), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_442), .B(n_412), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_434), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_434), .Y(n_487) );
OAI222xp33_ASAP7_75t_L g488 ( .A1(n_443), .A2(n_396), .B1(n_387), .B2(n_395), .C1(n_389), .C2(n_403), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_455), .A2(n_384), .B1(n_378), .B2(n_350), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_445), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_445), .Y(n_491) );
NOR2x1p5_ASAP7_75t_L g492 ( .A(n_432), .B(n_396), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_434), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_458), .A2(n_384), .B1(n_348), .B2(n_410), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_447), .Y(n_495) );
BUFx5_ASAP7_75t_L g496 ( .A(n_447), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_450), .Y(n_497) );
OAI222xp33_ASAP7_75t_L g498 ( .A1(n_444), .A2(n_403), .B1(n_389), .B2(n_395), .C1(n_387), .C2(n_410), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_434), .Y(n_499) );
BUFx12f_ASAP7_75t_L g500 ( .A(n_456), .Y(n_500) );
BUFx4f_ASAP7_75t_SL g501 ( .A(n_429), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_420), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_450), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_451), .B(n_390), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_418), .A2(n_384), .B1(n_395), .B2(n_387), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_439), .A2(n_384), .B1(n_378), .B2(n_441), .Y(n_506) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_439), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_419), .A2(n_384), .B1(n_405), .B2(n_410), .Y(n_508) );
OAI21xp5_ASAP7_75t_SL g509 ( .A1(n_432), .A2(n_266), .B(n_264), .Y(n_509) );
BUFx2_ASAP7_75t_L g510 ( .A(n_425), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_451), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_415), .B(n_390), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_439), .A2(n_378), .B1(n_350), .B2(n_355), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_415), .B(n_390), .Y(n_514) );
BUFx12f_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
OAI21xp5_ASAP7_75t_SL g516 ( .A1(n_432), .A2(n_279), .B(n_270), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_439), .A2(n_350), .B1(n_355), .B2(n_270), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_441), .A2(n_355), .B1(n_281), .B2(n_279), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_441), .A2(n_355), .B1(n_281), .B2(n_319), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_433), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_453), .B(n_319), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_433), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_441), .A2(n_355), .B1(n_319), .B2(n_351), .Y(n_523) );
AOI222xp33_ASAP7_75t_L g524 ( .A1(n_453), .A2(n_292), .B1(n_351), .B2(n_347), .C1(n_386), .C2(n_332), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_446), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_420), .B(n_390), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_437), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_421), .B(n_394), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_446), .A2(n_395), .B1(n_403), .B2(n_389), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_421), .B(n_394), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_446), .A2(n_292), .B1(n_347), .B2(n_386), .C1(n_332), .C2(n_335), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_452), .B(n_394), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_471), .A2(n_437), .B1(n_355), .B2(n_440), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_482), .B(n_452), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_494), .A2(n_440), .B1(n_386), .B2(n_395), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_460), .A2(n_403), .B1(n_389), .B2(n_395), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_482), .B(n_394), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_465), .A2(n_405), .B1(n_410), .B2(n_411), .Y(n_538) );
AOI222xp33_ASAP7_75t_L g539 ( .A1(n_463), .A2(n_292), .B1(n_347), .B2(n_335), .C1(n_177), .C2(n_172), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_468), .A2(n_177), .B1(n_173), .B2(n_172), .C(n_300), .Y(n_540) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_507), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_489), .A2(n_405), .B1(n_410), .B2(n_411), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_501), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_467), .A2(n_464), .B1(n_478), .B2(n_472), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_469), .A2(n_331), .B1(n_356), .B2(n_363), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_472), .A2(n_389), .B1(n_387), .B2(n_403), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_472), .A2(n_389), .B1(n_387), .B2(n_403), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_482), .B(n_406), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_475), .A2(n_389), .B1(n_387), .B2(n_403), .Y(n_549) );
OAI222xp33_ASAP7_75t_L g550 ( .A1(n_508), .A2(n_387), .B1(n_406), .B2(n_411), .C1(n_408), .C2(n_392), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g551 ( .A(n_461), .B(n_328), .C(n_337), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_513), .A2(n_411), .B1(n_408), .B2(n_406), .Y(n_552) );
AOI22xp5_ASAP7_75t_SL g553 ( .A1(n_462), .A2(n_408), .B1(n_406), .B2(n_374), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_476), .A2(n_408), .B1(n_402), .B2(n_363), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_487), .A2(n_407), .B1(n_379), .B2(n_413), .Y(n_555) );
OAI211xp5_ASAP7_75t_SL g556 ( .A1(n_524), .A2(n_328), .B(n_349), .C(n_323), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_487), .A2(n_402), .B1(n_356), .B2(n_352), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_504), .B(n_402), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_475), .A2(n_349), .B1(n_367), .B2(n_352), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_504), .B(n_402), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_475), .A2(n_367), .B1(n_356), .B2(n_363), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_487), .A2(n_402), .B1(n_248), .B2(n_254), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_531), .A2(n_367), .B1(n_248), .B2(n_254), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_523), .A2(n_382), .B1(n_381), .B2(n_413), .Y(n_564) );
OAI221xp5_ASAP7_75t_SL g565 ( .A1(n_480), .A2(n_306), .B1(n_305), .B2(n_323), .C(n_341), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_486), .A2(n_407), .B1(n_381), .B2(n_409), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_506), .A2(n_382), .B1(n_381), .B2(n_413), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_485), .B(n_354), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_521), .A2(n_382), .B1(n_409), .B2(n_413), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_459), .A2(n_382), .B1(n_409), .B2(n_413), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_470), .A2(n_409), .B1(n_401), .B2(n_398), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_486), .A2(n_409), .B1(n_401), .B2(n_398), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_486), .A2(n_401), .B1(n_398), .B2(n_404), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_492), .A2(n_401), .B1(n_398), .B2(n_376), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_483), .A2(n_366), .B1(n_359), .B2(n_354), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_529), .B(n_168), .C(n_164), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_474), .B(n_404), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_505), .A2(n_493), .B1(n_499), .B2(n_517), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_493), .A2(n_366), .B1(n_359), .B2(n_398), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_499), .A2(n_401), .B1(n_373), .B2(n_376), .Y(n_580) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_509), .A2(n_346), .B1(n_173), .B2(n_177), .C(n_172), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_477), .B(n_404), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_519), .A2(n_376), .B1(n_373), .B2(n_380), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_496), .A2(n_376), .B1(n_373), .B2(n_380), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_518), .A2(n_404), .B1(n_376), .B2(n_373), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_496), .A2(n_376), .B1(n_373), .B2(n_404), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_496), .A2(n_373), .B1(n_404), .B2(n_372), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_496), .A2(n_404), .B1(n_372), .B2(n_306), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_496), .A2(n_404), .B1(n_372), .B2(n_306), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_510), .A2(n_404), .B1(n_300), .B2(n_306), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_510), .A2(n_404), .B1(n_372), .B2(n_341), .Y(n_591) );
INVx4_ASAP7_75t_L g592 ( .A(n_496), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_520), .B(n_164), .C(n_166), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_496), .A2(n_404), .B1(n_372), .B2(n_305), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g595 ( .A1(n_462), .A2(n_515), .B1(n_500), .B2(n_484), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_525), .A2(n_404), .B1(n_372), .B2(n_305), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_525), .A2(n_507), .B1(n_500), .B2(n_515), .Y(n_597) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_341), .B1(n_302), .B2(n_346), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_490), .B(n_172), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g600 ( .A1(n_507), .A2(n_300), .B1(n_305), .B2(n_344), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_516), .A2(n_300), .B1(n_333), .B2(n_321), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_507), .A2(n_168), .B1(n_166), .B2(n_164), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_507), .A2(n_168), .B1(n_166), .B2(n_172), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_527), .A2(n_168), .B1(n_166), .B2(n_172), .Y(n_604) );
NAND2xp33_ASAP7_75t_L g605 ( .A(n_473), .B(n_329), .Y(n_605) );
OA21x2_ASAP7_75t_L g606 ( .A1(n_498), .A2(n_322), .B(n_327), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_466), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_520), .A2(n_168), .B1(n_166), .B2(n_172), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g609 ( .A1(n_522), .A2(n_158), .B(n_166), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_477), .A2(n_491), .B1(n_511), .B2(n_503), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_491), .A2(n_168), .B1(n_166), .B2(n_172), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_503), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_495), .B(n_172), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_497), .B(n_172), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_528), .A2(n_300), .B1(n_333), .B2(n_321), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_511), .B(n_528), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_532), .B(n_166), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_512), .A2(n_166), .B1(n_168), .B2(n_177), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_514), .A2(n_166), .B1(n_168), .B2(n_177), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_466), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g621 ( .A1(n_532), .A2(n_530), .B1(n_526), .B2(n_488), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_481), .B(n_172), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_479), .A2(n_173), .B1(n_177), .B2(n_168), .C(n_166), .Y(n_623) );
AOI222xp33_ASAP7_75t_L g624 ( .A1(n_481), .A2(n_173), .B1(n_177), .B2(n_168), .C1(n_344), .C2(n_298), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_502), .A2(n_168), .B1(n_173), .B2(n_177), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_502), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_494), .A2(n_173), .B1(n_177), .B2(n_325), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_494), .A2(n_173), .B1(n_177), .B2(n_325), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_494), .A2(n_173), .B1(n_177), .B2(n_344), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_474), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_482), .B(n_173), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_482), .B(n_173), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_494), .A2(n_173), .B1(n_344), .B2(n_302), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_460), .A2(n_307), .B1(n_342), .B2(n_309), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_616), .B(n_29), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_621), .A2(n_298), .B(n_301), .Y(n_636) );
OAI21xp33_ASAP7_75t_SL g637 ( .A1(n_592), .A2(n_250), .B(n_334), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_540), .B(n_158), .C(n_160), .Y(n_638) );
AND4x1_ASAP7_75t_L g639 ( .A(n_597), .B(n_30), .C(n_31), .D(n_32), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_554), .A2(n_333), .B1(n_298), .B2(n_301), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_612), .B(n_30), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_612), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_577), .B(n_158), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_630), .B(n_31), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_630), .B(n_33), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_578), .A2(n_250), .B(n_329), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_544), .A2(n_158), .B1(n_318), .B2(n_337), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_592), .B(n_158), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_556), .A2(n_158), .B1(n_160), .B2(n_295), .C(n_297), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_577), .B(n_158), .Y(n_650) );
AOI221x1_ASAP7_75t_SL g651 ( .A1(n_538), .A2(n_33), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_623), .B(n_158), .C(n_160), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_582), .B(n_158), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_582), .B(n_158), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_610), .B(n_34), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_620), .B(n_35), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_553), .A2(n_301), .B1(n_298), .B2(n_345), .Y(n_657) );
AND2x2_ASAP7_75t_SL g658 ( .A(n_592), .B(n_302), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_620), .B(n_37), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_607), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_581), .B(n_322), .C(n_295), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_576), .B(n_322), .C(n_327), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_631), .B(n_343), .C(n_340), .Y(n_663) );
OAI221xp5_ASAP7_75t_SL g664 ( .A1(n_533), .A2(n_301), .B1(n_295), .B2(n_324), .C(n_326), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_533), .A2(n_324), .B(n_326), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_632), .B(n_343), .C(n_340), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_537), .B(n_38), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_548), .B(n_39), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_607), .B(n_40), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_626), .B(n_41), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_617), .B(n_41), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g672 ( .A1(n_550), .A2(n_324), .B(n_326), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_617), .B(n_336), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_609), .B(n_309), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_536), .B(n_336), .C(n_343), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_543), .B(n_43), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_558), .B(n_336), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_560), .B(n_336), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_545), .B(n_340), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_549), .B(n_343), .C(n_340), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_545), .B(n_309), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_565), .A2(n_345), .B1(n_338), .B2(n_297), .C(n_302), .Y(n_682) );
OA21x2_ASAP7_75t_L g683 ( .A1(n_609), .A2(n_342), .B(n_309), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_534), .B(n_311), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_535), .B(n_311), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_626), .B(n_44), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_568), .B(n_311), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_599), .B(n_311), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_613), .B(n_317), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_614), .B(n_317), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_626), .B(n_47), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_552), .B(n_317), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_626), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_579), .B(n_317), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_542), .B(n_342), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_626), .B(n_50), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_590), .B(n_342), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_601), .A2(n_345), .B1(n_338), .B2(n_334), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_615), .B(n_324), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_615), .B(n_326), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_557), .B(n_561), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_595), .B(n_345), .C(n_338), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_606), .B(n_51), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_606), .B(n_52), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_586), .B(n_318), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_563), .B(n_318), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_606), .B(n_53), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_575), .B(n_318), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_606), .B(n_54), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_601), .B(n_591), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_546), .B(n_318), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_633), .A2(n_334), .B1(n_302), .B2(n_318), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_547), .B(n_318), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_541), .B(n_55), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_584), .B(n_329), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_629), .B(n_329), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_541), .B(n_56), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_608), .B(n_288), .C(n_287), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_627), .B(n_329), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g720 ( .A(n_628), .B(n_229), .C(n_234), .D(n_231), .Y(n_720) );
OAI21xp5_ASAP7_75t_SL g721 ( .A1(n_555), .A2(n_267), .B(n_320), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_541), .B(n_57), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_541), .B(n_59), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_541), .B(n_60), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_593), .B(n_288), .C(n_287), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_587), .B(n_329), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_588), .B(n_329), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_589), .B(n_329), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_594), .B(n_329), .Y(n_729) );
AND2x2_ASAP7_75t_SL g730 ( .A(n_605), .B(n_314), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_571), .B(n_61), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_622), .B(n_329), .Y(n_732) );
OAI221xp5_ASAP7_75t_SL g733 ( .A1(n_583), .A2(n_229), .B1(n_231), .B2(n_234), .C(n_232), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_551), .B(n_329), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_618), .B(n_314), .C(n_308), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_564), .B(n_62), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_585), .A2(n_276), .B1(n_280), .B2(n_320), .C(n_278), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_570), .B(n_63), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_572), .B(n_65), .Y(n_739) );
OR2x2_ASAP7_75t_L g740 ( .A(n_660), .B(n_634), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_642), .B(n_559), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_647), .A2(n_539), .B1(n_600), .B2(n_624), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_658), .B(n_574), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_642), .B(n_543), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_658), .B(n_569), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_710), .A2(n_562), .B1(n_605), .B2(n_580), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_660), .Y(n_747) );
AOI221x1_ASAP7_75t_SL g748 ( .A1(n_635), .A2(n_566), .B1(n_598), .B2(n_573), .C(n_619), .Y(n_748) );
INVxp67_ASAP7_75t_SL g749 ( .A(n_648), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_643), .B(n_567), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_643), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_650), .B(n_596), .Y(n_752) );
NAND3xp33_ASAP7_75t_L g753 ( .A(n_639), .B(n_604), .C(n_611), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_669), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_650), .B(n_625), .Y(n_755) );
NOR2x1_ASAP7_75t_L g756 ( .A(n_721), .B(n_320), .Y(n_756) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_655), .B(n_320), .C(n_280), .Y(n_757) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_639), .B(n_603), .C(n_602), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_669), .Y(n_759) );
OR2x2_ASAP7_75t_L g760 ( .A(n_653), .B(n_66), .Y(n_760) );
OA211x2_ASAP7_75t_L g761 ( .A1(n_646), .A2(n_70), .B(n_72), .C(n_73), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_701), .B(n_75), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_649), .A2(n_314), .B1(n_308), .B2(n_320), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_654), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_654), .B(n_684), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_651), .A2(n_280), .B1(n_320), .B2(n_308), .C(n_314), .Y(n_766) );
NAND4xp75_ASAP7_75t_L g767 ( .A(n_730), .B(n_77), .C(n_78), .D(n_79), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_636), .A2(n_314), .B1(n_308), .B2(n_245), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_693), .Y(n_769) );
AOI22xp33_ASAP7_75t_SL g770 ( .A1(n_730), .A2(n_308), .B1(n_314), .B2(n_267), .Y(n_770) );
OAI211xp5_ASAP7_75t_SL g771 ( .A1(n_657), .A2(n_245), .B(n_290), .C(n_265), .Y(n_771) );
AO21x2_ASAP7_75t_L g772 ( .A1(n_641), .A2(n_81), .B(n_83), .Y(n_772) );
AOI211xp5_ASAP7_75t_L g773 ( .A1(n_637), .A2(n_314), .B(n_308), .C(n_90), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_656), .B(n_88), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_659), .B(n_89), .Y(n_775) );
BUFx3_ASAP7_75t_L g776 ( .A(n_676), .Y(n_776) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_637), .B(n_648), .C(n_667), .Y(n_777) );
INVx2_ASAP7_75t_SL g778 ( .A(n_670), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_659), .B(n_91), .Y(n_779) );
NAND4xp75_ASAP7_75t_L g780 ( .A(n_703), .B(n_92), .C(n_93), .D(n_95), .Y(n_780) );
AO21x2_ASAP7_75t_L g781 ( .A1(n_644), .A2(n_98), .B(n_100), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_693), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_670), .B(n_101), .Y(n_783) );
NOR2xp33_ASAP7_75t_SL g784 ( .A(n_664), .B(n_308), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_672), .A2(n_308), .B1(n_314), .B2(n_272), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_668), .B(n_308), .C(n_314), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_645), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_686), .B(n_106), .Y(n_788) );
AO21x2_ASAP7_75t_L g789 ( .A1(n_703), .A2(n_107), .B(n_314), .Y(n_789) );
AND2x2_ASAP7_75t_L g790 ( .A(n_686), .B(n_272), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_671), .A2(n_272), .B1(n_665), .B2(n_733), .C(n_682), .Y(n_791) );
NAND3xp33_ASAP7_75t_L g792 ( .A(n_704), .B(n_707), .C(n_709), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_681), .B(n_687), .Y(n_793) );
NAND3xp33_ASAP7_75t_L g794 ( .A(n_704), .B(n_707), .C(n_709), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_694), .Y(n_795) );
AND2x4_ASAP7_75t_L g796 ( .A(n_691), .B(n_696), .Y(n_796) );
AOI211xp5_ASAP7_75t_L g797 ( .A1(n_698), .A2(n_674), .B(n_675), .C(n_702), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_679), .B(n_711), .Y(n_798) );
NAND4xp75_ASAP7_75t_L g799 ( .A(n_674), .B(n_731), .C(n_738), .D(n_739), .Y(n_799) );
INVxp67_ASAP7_75t_L g800 ( .A(n_683), .Y(n_800) );
NAND4xp75_ASAP7_75t_L g801 ( .A(n_731), .B(n_738), .C(n_739), .D(n_640), .Y(n_801) );
AO21x2_ASAP7_75t_L g802 ( .A1(n_691), .A2(n_696), .B(n_714), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_673), .B(n_678), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_680), .B(n_708), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g805 ( .A1(n_725), .A2(n_662), .B(n_735), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_714), .B(n_722), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_717), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_692), .Y(n_808) );
NOR3xp33_ASAP7_75t_L g809 ( .A(n_720), .B(n_638), .C(n_652), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_685), .Y(n_810) );
AO21x2_ASAP7_75t_L g811 ( .A1(n_717), .A2(n_724), .B(n_723), .Y(n_811) );
NAND3xp33_ASAP7_75t_L g812 ( .A(n_737), .B(n_734), .C(n_736), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_640), .A2(n_697), .B1(n_663), .B2(n_666), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g814 ( .A1(n_677), .A2(n_661), .B1(n_713), .B2(n_712), .C(n_705), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_695), .B(n_688), .Y(n_815) );
NAND4xp75_ASAP7_75t_L g816 ( .A(n_683), .B(n_722), .C(n_724), .D(n_723), .Y(n_816) );
NOR3xp33_ASAP7_75t_L g817 ( .A(n_718), .B(n_706), .C(n_699), .Y(n_817) );
NAND3xp33_ASAP7_75t_SL g818 ( .A(n_726), .B(n_715), .C(n_728), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_700), .B(n_689), .Y(n_819) );
AOI22xp33_ASAP7_75t_SL g820 ( .A1(n_683), .A2(n_727), .B1(n_729), .B2(n_690), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_732), .A2(n_422), .B1(n_428), .B2(n_423), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_747), .B(n_719), .Y(n_822) );
XOR2x2_ASAP7_75t_L g823 ( .A(n_801), .B(n_716), .Y(n_823) );
XNOR2xp5_ASAP7_75t_L g824 ( .A(n_744), .B(n_748), .Y(n_824) );
NAND4xp75_ASAP7_75t_L g825 ( .A(n_756), .B(n_805), .C(n_761), .D(n_762), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_787), .B(n_810), .Y(n_826) );
NAND4xp75_ASAP7_75t_SL g827 ( .A(n_804), .B(n_762), .C(n_743), .D(n_745), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_808), .B(n_795), .Y(n_828) );
NOR3xp33_ASAP7_75t_SL g829 ( .A(n_812), .B(n_799), .C(n_813), .Y(n_829) );
XNOR2xp5_ASAP7_75t_L g830 ( .A(n_744), .B(n_776), .Y(n_830) );
NAND4xp75_ASAP7_75t_L g831 ( .A(n_814), .B(n_785), .C(n_804), .D(n_768), .Y(n_831) );
AND2x4_ASAP7_75t_L g832 ( .A(n_778), .B(n_811), .Y(n_832) );
NAND4xp75_ASAP7_75t_L g833 ( .A(n_791), .B(n_766), .C(n_755), .D(n_783), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_754), .B(n_759), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_747), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_751), .Y(n_836) );
NAND4xp75_ASAP7_75t_L g837 ( .A(n_741), .B(n_750), .C(n_815), .D(n_793), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_764), .B(n_749), .Y(n_838) );
NAND4xp75_ASAP7_75t_L g839 ( .A(n_798), .B(n_774), .C(n_775), .D(n_779), .Y(n_839) );
XNOR2xp5_ASAP7_75t_L g840 ( .A(n_803), .B(n_752), .Y(n_840) );
INVx3_ASAP7_75t_L g841 ( .A(n_816), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_749), .B(n_819), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_802), .B(n_811), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_792), .A2(n_794), .B1(n_777), .B2(n_746), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_802), .B(n_807), .Y(n_845) );
OR2x2_ASAP7_75t_L g846 ( .A(n_765), .B(n_740), .Y(n_846) );
NOR4xp25_ASAP7_75t_L g847 ( .A(n_818), .B(n_746), .C(n_771), .D(n_786), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_769), .B(n_782), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_806), .B(n_796), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_800), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_800), .Y(n_851) );
BUFx2_ASAP7_75t_L g852 ( .A(n_796), .Y(n_852) );
NAND3xp33_ASAP7_75t_L g853 ( .A(n_820), .B(n_797), .C(n_773), .Y(n_853) );
INVx2_ASAP7_75t_SL g854 ( .A(n_789), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_820), .B(n_789), .Y(n_855) );
AND2x2_ASAP7_75t_L g856 ( .A(n_817), .B(n_757), .Y(n_856) );
NAND4xp75_ASAP7_75t_SL g857 ( .A(n_788), .B(n_784), .C(n_790), .D(n_780), .Y(n_857) );
NAND3xp33_ASAP7_75t_L g858 ( .A(n_809), .B(n_817), .C(n_757), .Y(n_858) );
XNOR2x2_ASAP7_75t_L g859 ( .A(n_767), .B(n_753), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_818), .Y(n_860) );
XNOR2xp5_ASAP7_75t_L g861 ( .A(n_742), .B(n_821), .Y(n_861) );
NOR2x1_ASAP7_75t_L g862 ( .A(n_772), .B(n_781), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_821), .B(n_809), .Y(n_863) );
INVx1_ASAP7_75t_SL g864 ( .A(n_760), .Y(n_864) );
NAND3xp33_ASAP7_75t_SL g865 ( .A(n_770), .B(n_742), .C(n_758), .Y(n_865) );
NAND4xp75_ASAP7_75t_L g866 ( .A(n_771), .B(n_756), .C(n_805), .D(n_761), .Y(n_866) );
OAI22xp33_ASAP7_75t_L g867 ( .A1(n_763), .A2(n_792), .B1(n_794), .B2(n_777), .Y(n_867) );
BUFx3_ASAP7_75t_L g868 ( .A(n_763), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_747), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_747), .Y(n_870) );
NOR2xp33_ASAP7_75t_SL g871 ( .A(n_776), .B(n_595), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_871), .B(n_861), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_846), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_846), .Y(n_874) );
INVx2_ASAP7_75t_SL g875 ( .A(n_830), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_867), .B(n_844), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_850), .Y(n_877) );
INVxp67_ASAP7_75t_L g878 ( .A(n_824), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_851), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_869), .Y(n_880) );
XOR2x2_ASAP7_75t_L g881 ( .A(n_861), .B(n_824), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_870), .Y(n_882) );
AND2x2_ASAP7_75t_L g883 ( .A(n_845), .B(n_843), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_838), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_848), .Y(n_885) );
OR2x2_ASAP7_75t_L g886 ( .A(n_835), .B(n_834), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_828), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_848), .Y(n_888) );
XNOR2x2_ASAP7_75t_L g889 ( .A(n_858), .B(n_865), .Y(n_889) );
OAI22xp33_ASAP7_75t_SL g890 ( .A1(n_841), .A2(n_860), .B1(n_852), .B2(n_832), .Y(n_890) );
INVx1_ASAP7_75t_SL g891 ( .A(n_830), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_845), .B(n_843), .Y(n_892) );
XNOR2x1_ASAP7_75t_L g893 ( .A(n_863), .B(n_827), .Y(n_893) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_836), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_826), .Y(n_895) );
XOR2x2_ASAP7_75t_L g896 ( .A(n_863), .B(n_823), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_822), .Y(n_897) );
OAI22xp33_ASAP7_75t_L g898 ( .A1(n_841), .A2(n_853), .B1(n_852), .B2(n_842), .Y(n_898) );
AOI22x1_ASAP7_75t_L g899 ( .A1(n_878), .A2(n_841), .B1(n_856), .B2(n_855), .Y(n_899) );
INVx2_ASAP7_75t_SL g900 ( .A(n_894), .Y(n_900) );
XNOR2xp5_ASAP7_75t_L g901 ( .A(n_881), .B(n_829), .Y(n_901) );
INVx1_ASAP7_75t_SL g902 ( .A(n_891), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_875), .A2(n_837), .B1(n_840), .B2(n_832), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_872), .A2(n_856), .B1(n_833), .B2(n_831), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_896), .A2(n_833), .B1(n_831), .B2(n_868), .Y(n_905) );
AO22x2_ASAP7_75t_L g906 ( .A1(n_875), .A2(n_855), .B1(n_854), .B2(n_832), .Y(n_906) );
INVx2_ASAP7_75t_SL g907 ( .A(n_873), .Y(n_907) );
OA22x2_ASAP7_75t_L g908 ( .A1(n_876), .A2(n_840), .B1(n_854), .B2(n_849), .Y(n_908) );
BUFx2_ASAP7_75t_L g909 ( .A(n_874), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_889), .B(n_825), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_888), .Y(n_911) );
HB1xp67_ASAP7_75t_L g912 ( .A(n_880), .Y(n_912) );
AOI22x1_ASAP7_75t_SL g913 ( .A1(n_889), .A2(n_859), .B1(n_864), .B2(n_857), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_893), .A2(n_866), .B1(n_825), .B2(n_862), .Y(n_914) );
INVxp33_ASAP7_75t_SL g915 ( .A(n_902), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_909), .Y(n_916) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_902), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_912), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_911), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_907), .Y(n_920) );
XOR2x2_ASAP7_75t_L g921 ( .A(n_901), .B(n_881), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_900), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_906), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_923), .A2(n_910), .B1(n_898), .B2(n_906), .C(n_903), .Y(n_924) );
INVx1_ASAP7_75t_SL g925 ( .A(n_917), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g926 ( .A1(n_915), .A2(n_905), .B1(n_904), .B2(n_893), .Y(n_926) );
NAND4xp25_ASAP7_75t_L g927 ( .A(n_915), .B(n_905), .C(n_904), .D(n_914), .Y(n_927) );
INVxp67_ASAP7_75t_L g928 ( .A(n_922), .Y(n_928) );
A2O1A1Ixp33_ASAP7_75t_SL g929 ( .A1(n_926), .A2(n_916), .B(n_918), .C(n_921), .Y(n_929) );
OAI211xp5_ASAP7_75t_L g930 ( .A1(n_927), .A2(n_899), .B(n_921), .C(n_920), .Y(n_930) );
INVxp67_ASAP7_75t_SL g931 ( .A(n_928), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_930), .A2(n_913), .B1(n_924), .B2(n_925), .Y(n_932) );
AO22x2_ASAP7_75t_L g933 ( .A1(n_931), .A2(n_919), .B1(n_896), .B2(n_892), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_929), .B(n_890), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_932), .A2(n_933), .B1(n_934), .B2(n_908), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_932), .B(n_887), .Y(n_936) );
NOR3xp33_ASAP7_75t_SL g937 ( .A(n_936), .B(n_866), .C(n_919), .Y(n_937) );
AND4x1_ASAP7_75t_L g938 ( .A(n_935), .B(n_847), .C(n_892), .D(n_883), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_938), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_937), .Y(n_940) );
AO22x2_ASAP7_75t_L g941 ( .A1(n_940), .A2(n_895), .B1(n_883), .B2(n_884), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_941), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_942), .A2(n_939), .B1(n_897), .B2(n_859), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_943), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_944), .A2(n_897), .B1(n_885), .B2(n_839), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_945), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_946), .A2(n_882), .B1(n_880), .B2(n_877), .C(n_879), .Y(n_947) );
AOI211xp5_ASAP7_75t_L g948 ( .A1(n_947), .A2(n_886), .B(n_885), .C(n_882), .Y(n_948) );
endmodule