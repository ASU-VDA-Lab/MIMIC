module fake_jpeg_26721_n_341 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_14),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_32),
.B1(n_23),
.B2(n_27),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_67),
.Y(n_78)
);

NAND2x1_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_17),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_17),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_43),
.B1(n_49),
.B2(n_45),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_70),
.A2(n_113),
.B1(n_83),
.B2(n_73),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_43),
.B1(n_40),
.B2(n_46),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_71),
.A2(n_77),
.B1(n_84),
.B2(n_96),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_73),
.B(n_83),
.Y(n_140)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_46),
.B1(n_32),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_86),
.B1(n_93),
.B2(n_108),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_32),
.B1(n_33),
.B2(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_90),
.Y(n_119)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_33),
.B1(n_27),
.B2(n_42),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_85),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_33),
.B1(n_44),
.B2(n_14),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_28),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_29),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_97),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_29),
.B1(n_28),
.B2(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_26),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_103),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_21),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_0),
.C(n_1),
.Y(n_135)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_25),
.B1(n_15),
.B2(n_30),
.Y(n_133)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_65),
.A2(n_18),
.B1(n_28),
.B2(n_31),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_65),
.A2(n_18),
.B1(n_31),
.B2(n_22),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_41),
.B1(n_15),
.B2(n_22),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_25),
.B1(n_30),
.B2(n_21),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_64),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_64),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_130),
.B1(n_148),
.B2(n_91),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_38),
.B1(n_36),
.B2(n_18),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_129),
.B1(n_143),
.B2(n_97),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_71),
.A2(n_38),
.B1(n_36),
.B2(n_19),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_36),
.B1(n_38),
.B2(n_15),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_76),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_137),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_138),
.B(n_78),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_48),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g144 ( 
.A1(n_99),
.A2(n_48),
.B1(n_47),
.B2(n_35),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_47),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_30),
.B1(n_47),
.B2(n_48),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_90),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_140),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_117),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_154),
.A2(n_171),
.B1(n_118),
.B2(n_35),
.Y(n_214)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_157),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_156),
.A2(n_159),
.B(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_161),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_179),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_164),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_151),
.B(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_170),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_100),
.C(n_92),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_180),
.C(n_128),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_101),
.B1(n_80),
.B2(n_88),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_149),
.B1(n_115),
.B2(n_123),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_103),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_150),
.B(n_136),
.Y(n_189)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_174),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_122),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_74),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_134),
.B(n_12),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_114),
.B(n_94),
.C(n_98),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_35),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_137),
.A2(n_87),
.B(n_85),
.C(n_106),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_185),
.B(n_72),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_183),
.Y(n_196)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_159),
.B(n_176),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_128),
.B1(n_146),
.B2(n_132),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_168),
.B1(n_154),
.B2(n_162),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_117),
.B(n_150),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_193),
.A2(n_213),
.B(n_182),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_206),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_203),
.B1(n_208),
.B2(n_214),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_123),
.B1(n_149),
.B2(n_146),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_132),
.B1(n_125),
.B2(n_142),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_142),
.B1(n_147),
.B2(n_118),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_216),
.B1(n_162),
.B2(n_174),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_21),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_180),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_156),
.A2(n_20),
.B1(n_19),
.B2(n_107),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_155),
.B(n_11),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_217),
.B(n_182),
.Y(n_246)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_232),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_173),
.B(n_165),
.C(n_181),
.D(n_179),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_221),
.A2(n_235),
.B(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_163),
.Y(n_223)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_234),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_227),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_243),
.B1(n_186),
.B2(n_200),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_170),
.Y(n_228)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_152),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_206),
.C(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_153),
.B(n_175),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_204),
.A2(n_195),
.B1(n_199),
.B2(n_216),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_184),
.B(n_185),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_188),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_188),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_203),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_220),
.A2(n_195),
.B1(n_199),
.B2(n_194),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_249),
.B1(n_251),
.B2(n_230),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_220),
.A2(n_232),
.B1(n_219),
.B2(n_235),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_194),
.B1(n_204),
.B2(n_193),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_225),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_260),
.A2(n_186),
.B1(n_191),
.B2(n_172),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_222),
.C(n_227),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_268),
.C(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_200),
.C(n_198),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_269),
.A2(n_238),
.B1(n_223),
.B2(n_228),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_270),
.A2(n_274),
.B1(n_279),
.B2(n_263),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_275),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_276),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_229),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_278),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_221),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_233),
.B1(n_197),
.B2(n_205),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_207),
.C(n_191),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_253),
.C(n_262),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_209),
.B(n_207),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_282),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_196),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_251),
.B(n_224),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_285),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_288),
.B1(n_253),
.B2(n_264),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_247),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_0),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_292),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_303),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_260),
.B1(n_261),
.B2(n_255),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_272),
.B1(n_279),
.B2(n_266),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_271),
.C(n_282),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_301),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_256),
.C(n_255),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_270),
.B(n_256),
.CI(n_259),
.CON(n_302),
.SN(n_302)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_302),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_248),
.C(n_264),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_298),
.A2(n_273),
.B1(n_278),
.B2(n_284),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_309),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_299),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_20),
.B(n_19),
.C(n_3),
.Y(n_308)
);

OAI321xp33_ASAP7_75t_L g322 ( 
.A1(n_308),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_20),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_312),
.C(n_298),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_289),
.A2(n_1),
.B(n_2),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_1),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_316),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_296),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_319),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_299),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_321),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_302),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_305),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_300),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_4),
.B(n_6),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_324),
.B(n_293),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_293),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_4),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_331),
.A2(n_332),
.B(n_333),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_319),
.B(n_308),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_328),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_334),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_325),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

OAI31xp33_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_308),
.A3(n_290),
.B(n_324),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_308),
.B1(n_309),
.B2(n_9),
.Y(n_341)
);


endmodule