module fake_jpeg_5841_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_23),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_51),
.Y(n_84)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_35),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_52),
.B(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_22),
.B1(n_26),
.B2(n_31),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_67),
.B1(n_29),
.B2(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_22),
.B1(n_26),
.B2(n_31),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_28),
.B1(n_33),
.B2(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_29),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_23),
.C(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_22),
.B1(n_24),
.B2(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_73),
.B(n_76),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_45),
.B1(n_19),
.B2(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_68),
.Y(n_96)
);

OAI22x1_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_29),
.B1(n_63),
.B2(n_27),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_43),
.B(n_36),
.C(n_29),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_21),
.B1(n_18),
.B2(n_30),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_90),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_54),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_99),
.B1(n_102),
.B2(n_117),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_84),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_91),
.B(n_86),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_101),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_70),
.B1(n_68),
.B2(n_55),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_60),
.B1(n_59),
.B2(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_113),
.Y(n_134)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_66),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_51),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_51),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_58),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_90),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_79),
.A2(n_64),
.B1(n_63),
.B2(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_78),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_113),
.A2(n_79),
.B1(n_94),
.B2(n_76),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_123),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_116),
.A2(n_94),
.B1(n_81),
.B2(n_72),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_127),
.B(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_132),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_36),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_72),
.B1(n_83),
.B2(n_89),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_114),
.B1(n_103),
.B2(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_43),
.A3(n_36),
.B1(n_72),
.B2(n_94),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_81),
.B(n_71),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_140),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_139),
.B(n_110),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_43),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_99),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_96),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_100),
.B1(n_98),
.B2(n_114),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_139),
.B(n_137),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_150),
.B(n_125),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_164),
.B1(n_120),
.B2(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_156),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_138),
.A2(n_109),
.B(n_97),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_133),
.B(n_126),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_95),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_165),
.C(n_167),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_160),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_105),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_95),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_117),
.B1(n_86),
.B2(n_78),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_71),
.C(n_106),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_152),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_20),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_182),
.B1(n_165),
.B2(n_145),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_132),
.B1(n_135),
.B2(n_141),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_173),
.B(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_179),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_127),
.B(n_136),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_127),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_180),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_190)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_163),
.B1(n_166),
.B2(n_147),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_133),
.B1(n_124),
.B2(n_143),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_145),
.A2(n_124),
.B1(n_21),
.B2(n_30),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_188),
.A2(n_186),
.B(n_179),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_197),
.B1(n_199),
.B2(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_172),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_192),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_201),
.B(n_204),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_150),
.B1(n_153),
.B2(n_167),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_144),
.B1(n_150),
.B2(n_154),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_20),
.C(n_21),
.Y(n_200)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_2),
.C(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_30),
.B1(n_18),
.B2(n_20),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_171),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_168),
.A2(n_20),
.B1(n_0),
.B2(n_3),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_187),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_206),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_173),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_175),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_208),
.C(n_210),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_187),
.C(n_174),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_193),
.B(n_201),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_170),
.C(n_176),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_170),
.C(n_0),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_217),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_2),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_190),
.CI(n_198),
.CON(n_218),
.SN(n_218)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_222),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_211),
.B1(n_206),
.B2(n_212),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_188),
.B(n_194),
.C(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_191),
.B(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_204),
.Y(n_223)
);

OAI221xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_7),
.C(n_11),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_217),
.B(n_4),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_231),
.C(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_208),
.C(n_207),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_213),
.B1(n_9),
.B2(n_11),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_232),
.A2(n_7),
.B(n_11),
.C(n_12),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_7),
.C(n_9),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_221),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_218),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_236),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_222),
.B1(n_218),
.B2(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_225),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_12),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_225),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_231),
.C(n_238),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_16),
.C(n_13),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_239),
.B(n_14),
.C(n_15),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_13),
.B(n_14),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

OAI311xp33_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_241),
.A3(n_246),
.B1(n_247),
.C1(n_13),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_15),
.B(n_16),
.Y(n_250)
);


endmodule