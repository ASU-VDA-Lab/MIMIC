module real_jpeg_24166_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_0),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_0),
.A2(n_34),
.B1(n_61),
.B2(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_0),
.A2(n_34),
.B1(n_55),
.B2(n_56),
.Y(n_351)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_61),
.B1(n_65),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_2),
.A2(n_39),
.B1(n_41),
.B2(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_70),
.B1(n_84),
.B2(n_130),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_84),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_5),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_6),
.A2(n_61),
.B1(n_65),
.B2(n_72),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_6),
.A2(n_39),
.B1(n_41),
.B2(n_72),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_72),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_7),
.A2(n_48),
.B1(n_61),
.B2(n_65),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_7),
.A2(n_48),
.B1(n_130),
.B2(n_131),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_8),
.A2(n_70),
.B1(n_71),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_8),
.A2(n_61),
.B1(n_65),
.B2(n_160),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_8),
.A2(n_39),
.B1(n_41),
.B2(n_160),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_160),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_9),
.A2(n_55),
.B1(n_71),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_9),
.A2(n_61),
.B1(n_65),
.B2(n_106),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_9),
.A2(n_39),
.B1(n_41),
.B2(n_106),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_106),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_11),
.A2(n_58),
.B1(n_61),
.B2(n_65),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_11),
.A2(n_39),
.B1(n_41),
.B2(n_58),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_58),
.Y(n_222)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_13),
.B(n_70),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_13),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_13),
.B(n_60),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_13),
.B(n_39),
.C(n_80),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_13),
.A2(n_61),
.B1(n_65),
.B2(n_213),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_13),
.B(n_121),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_13),
.A2(n_39),
.B1(n_41),
.B2(n_213),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_13),
.B(n_26),
.C(n_44),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_13),
.A2(n_25),
.B(n_272),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_38),
.B1(n_61),
.B2(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_38),
.B1(n_56),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_16),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_347),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_334),
.B(n_346),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_134),
.A3(n_150),
.B(n_331),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_110),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_21),
.B(n_110),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_22),
.A2(n_75),
.B1(n_76),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_22),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_23),
.A2(n_24),
.B(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_24),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_25),
.A2(n_30),
.B1(n_33),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_25),
.A2(n_96),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_25),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_25),
.A2(n_189),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_25),
.B(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_25),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_27),
.B1(n_44),
.B2(n_45),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_27),
.B(n_297),
.Y(n_296)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_29),
.Y(n_170)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_29),
.Y(n_299)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_37),
.A2(n_42),
.B1(n_49),
.B2(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g41 ( 
.A(n_39),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_39),
.A2(n_41),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_39),
.B(n_279),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_42),
.A2(n_49),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_42),
.B(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_42),
.A2(n_49),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_46),
.A2(n_87),
.B1(n_100),
.B2(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_46),
.A2(n_172),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_46),
.A2(n_209),
.B(n_245),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_46),
.B(n_213),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_49),
.B(n_210),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_59),
.B(n_67),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_54),
.A2(n_59),
.B1(n_107),
.B2(n_129),
.Y(n_128)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_63),
.B1(n_66),
.B2(n_70),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_56),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_59),
.A2(n_107),
.B1(n_129),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_59),
.A2(n_67),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_60),
.A2(n_73),
.B1(n_105),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_60),
.A2(n_73),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_60),
.A2(n_73),
.B1(n_342),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_65),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_61),
.B(n_66),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_61),
.B(n_238),
.Y(n_237)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g183 ( 
.A1(n_63),
.A2(n_65),
.A3(n_71),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_73),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_73),
.A2(n_109),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_90),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_85),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_78),
.A2(n_79),
.B1(n_123),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_78),
.A2(n_179),
.B(n_181),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_78),
.A2(n_181),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_79),
.A2(n_102),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_79),
.A2(n_163),
.B(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_87),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_87),
.A2(n_260),
.B(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_89),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_91),
.A2(n_92),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_101),
.C(n_103),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_93),
.A2(n_94),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_95),
.A2(n_97),
.B1(n_98),
.B2(n_174),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_95),
.Y(n_174)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_101),
.B(n_103),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B(n_108),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_113),
.C(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_128),
.B2(n_133),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_125),
.C(n_128),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_120),
.A2(n_121),
.B1(n_180),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_120),
.A2(n_121),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_121),
.B(n_164),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_125),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_125),
.B(n_141),
.C(n_147),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_128),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_133),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_128),
.B(n_137),
.C(n_140),
.Y(n_335)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_135),
.A2(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_149),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_136),
.B(n_149),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_142),
.Y(n_341)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_148),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_324),
.B(n_330),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_198),
.B(n_323),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_191),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_153),
.B(n_191),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_173),
.C(n_175),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_154),
.A2(n_155),
.B1(n_173),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_161),
.C(n_165),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_171),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_187),
.B1(n_188),
.B2(n_190),
.Y(n_186)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_170),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_173),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_175),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_176),
.B(n_178),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_182),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_186),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_187),
.A2(n_283),
.B1(n_285),
.B2(n_287),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_193),
.B(n_194),
.C(n_197),
.Y(n_329)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_230),
.B(n_317),
.C(n_322),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_224),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_224),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_215),
.C(n_216),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_201),
.A2(n_202),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_211),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_207),
.C(n_211),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_213),
.B(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_215),
.B(n_216),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.C(n_221),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_311),
.B(n_316),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_261),
.B(n_310),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_250),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_235),
.B(n_250),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_243),
.C(n_247),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_236),
.B(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_243),
.A2(n_247),
.B1(n_248),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_243),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_251),
.B(n_257),
.C(n_258),
.Y(n_315)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_304),
.B(n_309),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_280),
.B(n_303),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_274),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_274),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_269),
.C(n_270),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_290),
.B(n_302),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_288),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_286),
.B(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_295),
.B(n_301),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_293),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_300),
.Y(n_295)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_308),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_329),
.Y(n_330)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_345),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_340),
.B1(n_343),
.B2(n_344),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_338),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_340),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_343),
.C(n_345),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_352),
.Y(n_353)
);


endmodule