module fake_jpeg_7510_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_19),
.B1(n_30),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_27),
.B1(n_26),
.B2(n_23),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_17),
.B1(n_33),
.B2(n_34),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_57),
.B1(n_69),
.B2(n_27),
.Y(n_97)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_21),
.B1(n_30),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_21),
.B1(n_30),
.B2(n_28),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_28),
.B(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_65),
.Y(n_78)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_67),
.Y(n_84)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_31),
.B1(n_20),
.B2(n_22),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_73),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_42),
.B1(n_31),
.B2(n_22),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_76),
.B1(n_64),
.B2(n_56),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_43),
.C(n_40),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_44),
.C(n_62),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_22),
.B1(n_31),
.B2(n_34),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_39),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_26),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_85),
.Y(n_124)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_88),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_58),
.B1(n_19),
.B2(n_24),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_96),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_33),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_98),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_24),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_24),
.B1(n_19),
.B2(n_25),
.Y(n_127)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_0),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_72),
.B1(n_73),
.B2(n_89),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_105),
.B(n_114),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_125),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_40),
.C(n_44),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_118),
.C(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_115),
.B(n_120),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_44),
.C(n_16),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_44),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_99),
.B(n_103),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_71),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_79),
.A2(n_34),
.B1(n_33),
.B2(n_17),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_129),
.A2(n_96),
.B1(n_77),
.B2(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_138),
.B1(n_136),
.B2(n_145),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_142),
.B1(n_156),
.B2(n_160),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_131),
.A2(n_97),
.B1(n_76),
.B2(n_74),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_152),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_78),
.B(n_81),
.C(n_103),
.D(n_101),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_122),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_82),
.B1(n_102),
.B2(n_86),
.Y(n_142)
);

BUFx8_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_149),
.B(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_161),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_150),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_99),
.B(n_80),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_81),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_99),
.B(n_92),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_98),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_25),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_162),
.B(n_146),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_25),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_105),
.C(n_114),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_123),
.B1(n_107),
.B2(n_110),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_93),
.B1(n_89),
.B2(n_86),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_158),
.B1(n_164),
.B2(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_90),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_121),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_88),
.B1(n_34),
.B2(n_33),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

OAI21x1_ASAP7_75t_SL g162 ( 
.A1(n_119),
.A2(n_32),
.B(n_17),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_165),
.B(n_167),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_118),
.B(n_111),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_168),
.B(n_179),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_108),
.B(n_119),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_185),
.C(n_14),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_129),
.B1(n_122),
.B2(n_112),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_174),
.A2(n_197),
.B1(n_198),
.B2(n_5),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_181),
.B1(n_143),
.B2(n_14),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_154),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_112),
.B(n_120),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_184),
.Y(n_223)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_124),
.C(n_121),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_194),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_32),
.B(n_17),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_32),
.B(n_3),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_124),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_199),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_138),
.A2(n_83),
.B1(n_3),
.B2(n_4),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_155),
.A2(n_83),
.B1(n_3),
.B2(n_4),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_189),
.A2(n_141),
.B1(n_133),
.B2(n_150),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_205),
.A2(n_214),
.B1(n_221),
.B2(n_198),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_15),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_215),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_176),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_133),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_170),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_196),
.B1(n_180),
.B2(n_195),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_220),
.C(n_173),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_184),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_14),
.C(n_13),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_171),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_228),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_13),
.B1(n_12),
.B2(n_7),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_225),
.B1(n_226),
.B2(n_192),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_5),
.C(n_6),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_175),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_172),
.A2(n_197),
.B1(n_174),
.B2(n_187),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_SL g261 ( 
.A1(n_229),
.A2(n_230),
.B(n_232),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_202),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_235),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_169),
.B1(n_172),
.B2(n_165),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_243),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_166),
.B(n_179),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_240),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_200),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_237),
.B(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_242),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_224),
.A2(n_168),
.B(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_244),
.C(n_248),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_188),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_188),
.C(n_193),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_205),
.A2(n_199),
.B1(n_180),
.B2(n_9),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_246),
.A2(n_249),
.B1(n_217),
.B2(n_225),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_7),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_221),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_11),
.C(n_8),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_220),
.C(n_211),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_253),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_213),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_255),
.B(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_SL g264 ( 
.A(n_236),
.B(n_218),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_246),
.B(n_238),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_268),
.C(n_271),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_207),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_240),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_274),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_207),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_241),
.B(n_212),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_273),
.C(n_252),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_204),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_230),
.Y(n_274)
);

BUFx12_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_287),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_232),
.B1(n_242),
.B2(n_251),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_282),
.B(n_283),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_256),
.B(n_204),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_214),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_285),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_249),
.B1(n_216),
.B2(n_201),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_233),
.C(n_206),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_290),
.B(n_239),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_263),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_259),
.B(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_273),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_258),
.C(n_263),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_297),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_277),
.A2(n_280),
.B(n_279),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_278),
.B(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_290),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_302),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_268),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_258),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_271),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_298),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_291),
.B(n_281),
.Y(n_307)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_275),
.B(n_304),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_287),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_309),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_267),
.B1(n_275),
.B2(n_276),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_310),
.A2(n_8),
.B1(n_11),
.B2(n_307),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_315),
.B1(n_300),
.B2(n_292),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_213),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_316),
.C(n_11),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_302),
.C(n_10),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_272),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_293),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_321),
.C(n_322),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_324),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_310),
.B1(n_308),
.B2(n_314),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_301),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_323),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_328),
.B(n_323),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_317),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_331),
.B(n_332),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_327),
.A2(n_321),
.B(n_322),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_325),
.B1(n_326),
.B2(n_314),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_325),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_11),
.Y(n_337)
);


endmodule