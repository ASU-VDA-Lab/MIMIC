module fake_jpeg_4288_n_216 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_40),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_0),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_53),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_33),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_16),
.B1(n_30),
.B2(n_28),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_37),
.B1(n_28),
.B2(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_64),
.Y(n_75)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_69),
.A2(n_76),
.B1(n_31),
.B2(n_17),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_30),
.B1(n_16),
.B2(n_39),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_39),
.B1(n_41),
.B2(n_21),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_74),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_19),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_82),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_34),
.B(n_29),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_40),
.B1(n_26),
.B2(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_89),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_17),
.C(n_31),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_97),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_70),
.B1(n_17),
.B2(n_55),
.Y(n_128)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_61),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_103),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_105),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_67),
.B(n_77),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_60),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_47),
.B1(n_34),
.B2(n_55),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_104),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_33),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_44),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_65),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_17),
.B1(n_19),
.B2(n_24),
.Y(n_150)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_79),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_65),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_60),
.B(n_90),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_81),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_68),
.Y(n_144)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_127),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_44),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_87),
.C(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_95),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_91),
.B1(n_98),
.B2(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_150),
.B1(n_120),
.B2(n_127),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_88),
.C(n_91),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_143),
.C(n_145),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_36),
.B(n_60),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_148),
.B(n_149),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_139),
.B(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_70),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_68),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_112),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_155),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_160),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_124),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_130),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_166),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_110),
.C(n_111),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_129),
.B1(n_110),
.B2(n_121),
.Y(n_161)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_141),
.B(n_149),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_165),
.B(n_134),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_123),
.B(n_114),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_128),
.C(n_123),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_134),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_173),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_145),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_178),
.C(n_151),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_179),
.B(n_36),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_180),
.B(n_19),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_157),
.Y(n_178)
);

AO221x1_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_86),
.B1(n_147),
.B2(n_144),
.C(n_82),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_159),
.B(n_143),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_184),
.C(n_186),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_166),
.B1(n_160),
.B2(n_158),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_151),
.C(n_153),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_168),
.B(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_82),
.C(n_66),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_189),
.C(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_66),
.C(n_36),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_189),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_173),
.B1(n_171),
.B2(n_167),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_197),
.B(n_188),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_174),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_198),
.A2(n_184),
.B(n_182),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_66),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_200),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_204),
.B(n_4),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_203),
.C(n_205),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_11),
.B(n_14),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_195),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_8),
.C2(n_5),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_13),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_4),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_208),
.C(n_7),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_206),
.C(n_6),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_211),
.A2(n_212),
.B(n_213),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_5),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_6),
.B(n_8),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_8),
.Y(n_216)
);


endmodule