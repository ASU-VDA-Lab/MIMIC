module fake_jpeg_24745_n_348 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_8),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_44),
.B(n_48),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_39),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_20),
.B1(n_22),
.B2(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_0),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_61),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_65),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_67),
.B1(n_40),
.B2(n_22),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_23),
.B1(n_21),
.B2(n_36),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_23),
.B1(n_21),
.B2(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_64),
.Y(n_104)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_23),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_17),
.B1(n_34),
.B2(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_75),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_74),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_76),
.B(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_84),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_52),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_97),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_27),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_86),
.B1(n_92),
.B2(n_93),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_46),
.B1(n_29),
.B2(n_31),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_87),
.Y(n_124)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_46),
.B1(n_29),
.B2(n_31),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_96),
.B1(n_32),
.B2(n_18),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_27),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_48),
.B1(n_35),
.B2(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_48),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_106),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_37),
.B(n_25),
.C(n_29),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_29),
.C(n_19),
.Y(n_114)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

BUFx4f_ASAP7_75t_SL g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_51),
.B(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_68),
.B1(n_49),
.B2(n_50),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_118),
.B1(n_128),
.B2(n_129),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_120),
.B(n_99),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_19),
.B(n_31),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_102),
.B(n_81),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_49),
.B1(n_61),
.B2(n_69),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_71),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_16),
.C(n_13),
.Y(n_158)
);

NOR2x1_ASAP7_75t_R g120 ( 
.A(n_84),
.B(n_39),
.Y(n_120)
);

OA22x2_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_39),
.B1(n_71),
.B2(n_28),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_121),
.A2(n_106),
.B(n_82),
.C(n_18),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_39),
.Y(n_123)
);

NAND2x1_ASAP7_75t_SL g159 ( 
.A(n_123),
.B(n_101),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_35),
.B1(n_71),
.B2(n_28),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_93),
.A2(n_28),
.B1(n_26),
.B2(n_34),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_105),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_24),
.C(n_28),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_102),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_90),
.B1(n_78),
.B2(n_76),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_137),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_139),
.B(n_141),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_88),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_159),
.B(n_120),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_121),
.B1(n_114),
.B2(n_136),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_164),
.B1(n_167),
.B2(n_128),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_151),
.Y(n_181)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_88),
.A3(n_96),
.B1(n_102),
.B2(n_77),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_32),
.B(n_18),
.C(n_25),
.D(n_11),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_89),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_133),
.C(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_155),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_165),
.B(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_161),
.B1(n_162),
.B2(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

AO21x2_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_74),
.B(n_91),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_119),
.A2(n_73),
.B(n_80),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_32),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_100),
.B1(n_32),
.B2(n_18),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_179),
.B1(n_182),
.B2(n_190),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_169),
.A2(n_188),
.B(n_189),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_172),
.C(n_175),
.Y(n_220)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_124),
.C(n_116),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_130),
.C(n_126),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_129),
.B1(n_108),
.B2(n_126),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_201),
.B1(n_9),
.B2(n_14),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_178),
.B(n_185),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_134),
.B1(n_125),
.B2(n_117),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_197),
.B(n_198),
.Y(n_203)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_187),
.B(n_196),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_125),
.B(n_135),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_154),
.A2(n_74),
.B(n_117),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_74),
.B1(n_117),
.B2(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_24),
.Y(n_193)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_24),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_138),
.B(n_24),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_164),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_25),
.B(n_2),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_7),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_143),
.B(n_164),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_204),
.A2(n_206),
.B(n_232),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_227),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_164),
.B(n_153),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_1),
.Y(n_211)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_216),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_219),
.B1(n_15),
.B2(n_232),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_223),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_171),
.A2(n_3),
.B1(n_4),
.B2(n_15),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_231),
.B1(n_177),
.B2(n_173),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_4),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_181),
.B(n_6),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_230),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_191),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_229),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_7),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_168),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_183),
.A2(n_9),
.B(n_13),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_194),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_234),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_170),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_172),
.C(n_175),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_237),
.C(n_241),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_188),
.B1(n_169),
.B2(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_195),
.C(n_197),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_209),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_221),
.C(n_206),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_207),
.A2(n_216),
.B1(n_223),
.B2(n_224),
.Y(n_243)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_198),
.C(n_199),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_203),
.C(n_219),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_208),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_247),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_205),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_192),
.B1(n_202),
.B2(n_14),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_249),
.A2(n_258),
.B1(n_252),
.B2(n_238),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_229),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_254),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_230),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_213),
.A2(n_15),
.B1(n_226),
.B2(n_204),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_245),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_267),
.C(n_270),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_221),
.C(n_203),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_209),
.C(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_278),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_212),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_276),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_249),
.B1(n_242),
.B2(n_255),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_240),
.B(n_214),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_275),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_236),
.B(n_217),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_227),
.C(n_228),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_252),
.C(n_242),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_240),
.B(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_239),
.B1(n_256),
.B2(n_258),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_283),
.A2(n_287),
.B1(n_259),
.B2(n_278),
.Y(n_304)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_237),
.B1(n_256),
.B2(n_243),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_246),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_272),
.Y(n_306)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_295),
.B1(n_297),
.B2(n_280),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_294),
.C(n_296),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_257),
.C(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_257),
.C(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_274),
.Y(n_299)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_265),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_282),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_283),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_298),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_309),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_289),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_263),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_307),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_308),
.B(n_312),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_288),
.B(n_259),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_264),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_313),
.B(n_285),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_267),
.B(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_316),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_285),
.B(n_293),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_324),
.Y(n_329)
);

AO22x1_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_301),
.B1(n_303),
.B2(n_295),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_311),
.B(n_297),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_330),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_331),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_322),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_300),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_325),
.A2(n_290),
.B(n_306),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_332),
.A2(n_330),
.B(n_326),
.Y(n_340)
);

AOI31xp33_ASAP7_75t_L g334 ( 
.A1(n_316),
.A2(n_281),
.A3(n_290),
.B(n_317),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_324),
.B(n_327),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_314),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_335),
.B(n_339),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_333),
.A2(n_320),
.B1(n_315),
.B2(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_340),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_342),
.B(n_343),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_345),
.A2(n_341),
.B(n_338),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_337),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_337),
.Y(n_348)
);


endmodule