module real_aes_17979_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_887;
wire n_599;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_552;
wire n_590;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1250;
wire n_1095;
wire n_360;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_315;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1129;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1163;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1162;
wire n_762;
wire n_325;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_832;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_974;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_304;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_244;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1252;
wire n_269;
wire n_430;
wire n_1132;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_338;
wire n_698;
wire n_371;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_0), .A2(n_179), .B1(n_1000), .B2(n_1002), .Y(n_1052) );
OAI22xp33_ASAP7_75t_SL g358 ( .A1(n_1), .A2(n_105), .B1(n_359), .B2(n_362), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g395 ( .A1(n_1), .A2(n_22), .B1(n_396), .B2(n_397), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_2), .A2(n_24), .B1(n_352), .B2(n_750), .Y(n_879) );
OAI22xp5_ASAP7_75t_SL g887 ( .A1(n_2), .A2(n_110), .B1(n_375), .B2(n_396), .Y(n_887) );
INVx1_ASAP7_75t_L g722 ( .A(n_3), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_4), .A2(n_54), .B1(n_1000), .B2(n_1002), .Y(n_1020) );
OAI22xp33_ASAP7_75t_L g959 ( .A1(n_5), .A2(n_160), .B1(n_352), .B2(n_362), .Y(n_959) );
OAI22xp33_ASAP7_75t_SL g969 ( .A1(n_5), .A2(n_160), .B1(n_396), .B2(n_754), .Y(n_969) );
INVx1_ASAP7_75t_L g576 ( .A(n_6), .Y(n_576) );
OAI211xp5_ASAP7_75t_L g581 ( .A1(n_6), .A2(n_582), .B(n_583), .C(n_584), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_7), .Y(n_882) );
INVx1_ASAP7_75t_L g776 ( .A(n_8), .Y(n_776) );
OAI211xp5_ASAP7_75t_L g898 ( .A1(n_9), .A2(n_333), .B(n_488), .C(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g909 ( .A(n_9), .Y(n_909) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_10), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_11), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g329 ( .A(n_11), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_12), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_13), .A2(n_186), .B1(n_543), .B2(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_13), .A2(n_186), .B1(n_676), .B2(n_678), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_14), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_15), .Y(n_276) );
INVx1_ASAP7_75t_L g505 ( .A(n_16), .Y(n_505) );
INVx1_ASAP7_75t_L g915 ( .A(n_17), .Y(n_915) );
INVx2_ASAP7_75t_L g992 ( .A(n_18), .Y(n_992) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_18), .B(n_91), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_18), .B(n_993), .Y(n_1007) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_19), .A2(n_225), .B1(n_788), .B2(n_791), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_19), .A2(n_23), .B1(n_814), .B2(n_819), .Y(n_826) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_20), .A2(n_130), .B1(n_539), .B2(n_540), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_20), .A2(n_130), .B1(n_547), .B2(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g836 ( .A(n_21), .Y(n_836) );
OAI22xp33_ASAP7_75t_SL g351 ( .A1(n_22), .A2(n_215), .B1(n_352), .B2(n_355), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_23), .A2(n_162), .B1(n_793), .B2(n_798), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_24), .B(n_373), .Y(n_886) );
AO22x2_ASAP7_75t_L g933 ( .A1(n_25), .A2(n_934), .B1(n_974), .B2(n_975), .Y(n_933) );
INVx1_ASAP7_75t_L g974 ( .A(n_25), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g1029 ( .A1(n_25), .A2(n_35), .B1(n_1005), .B2(n_1006), .Y(n_1029) );
INVx1_ASAP7_75t_L g773 ( .A(n_26), .Y(n_773) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_27), .A2(n_140), .B1(n_362), .B2(n_455), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_27), .A2(n_227), .B1(n_396), .B2(n_397), .Y(n_457) );
INVx1_ASAP7_75t_L g479 ( .A(n_28), .Y(n_479) );
XOR2xp5_ASAP7_75t_L g239 ( .A(n_29), .B(n_240), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_29), .A2(n_104), .B1(n_1005), .B2(n_1006), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_30), .A2(n_157), .B1(n_362), .B2(n_543), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_30), .A2(n_157), .B1(n_397), .B2(n_840), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_31), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g751 ( .A1(n_32), .A2(n_127), .B1(n_352), .B2(n_666), .Y(n_751) );
OAI22xp33_ASAP7_75t_SL g753 ( .A1(n_32), .A2(n_127), .B1(n_396), .B2(n_754), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_33), .Y(n_867) );
INVx1_ASAP7_75t_L g939 ( .A(n_34), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_36), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_37), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_38), .A2(n_89), .B1(n_1000), .B2(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g712 ( .A(n_39), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g1026 ( .A1(n_40), .A2(n_86), .B1(n_1000), .B2(n_1017), .Y(n_1026) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_41), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_42), .A2(n_154), .B1(n_362), .B2(n_543), .Y(n_542) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_42), .A2(n_154), .B1(n_559), .B2(n_561), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_43), .Y(n_415) );
INVx1_ASAP7_75t_L g606 ( .A(n_44), .Y(n_606) );
XOR2x2_ASAP7_75t_L g783 ( .A(n_45), .B(n_784), .Y(n_783) );
XNOR2xp5_ASAP7_75t_L g471 ( .A(n_46), .B(n_472), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_47), .Y(n_864) );
INVx1_ASAP7_75t_L g832 ( .A(n_48), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g897 ( .A1(n_49), .A2(n_109), .B1(n_455), .B2(n_750), .Y(n_897) );
OAI22xp33_ASAP7_75t_L g910 ( .A1(n_49), .A2(n_55), .B1(n_375), .B2(n_397), .Y(n_910) );
INVx1_ASAP7_75t_L g748 ( .A(n_50), .Y(n_748) );
INVx1_ASAP7_75t_L g257 ( .A(n_51), .Y(n_257) );
INVx1_ASAP7_75t_L g263 ( .A(n_51), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_52), .A2(n_122), .B1(n_561), .B2(n_676), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g707 ( .A1(n_52), .A2(n_122), .B1(n_362), .B2(n_543), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_53), .A2(n_114), .B1(n_1000), .B2(n_1017), .Y(n_1016) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_55), .A2(n_184), .B1(n_352), .B2(n_666), .Y(n_902) );
INVx1_ASAP7_75t_L g650 ( .A(n_56), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_57), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_58), .A2(n_94), .B1(n_455), .B2(n_967), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g973 ( .A1(n_58), .A2(n_94), .B1(n_373), .B2(n_375), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_59), .A2(n_199), .B1(n_1005), .B2(n_1006), .Y(n_1091) );
INVx1_ASAP7_75t_L g644 ( .A(n_60), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_61), .A2(n_176), .B1(n_1212), .B2(n_1223), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_61), .A2(n_185), .B1(n_1236), .B2(n_1240), .Y(n_1242) );
INVx1_ASAP7_75t_L g487 ( .A(n_62), .Y(n_487) );
INVx1_ASAP7_75t_L g981 ( .A(n_63), .Y(n_981) );
INVx2_ASAP7_75t_L g250 ( .A(n_64), .Y(n_250) );
XNOR2x2_ASAP7_75t_L g635 ( .A(n_65), .B(n_636), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_66), .A2(n_200), .B1(n_540), .B2(n_589), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_66), .A2(n_200), .B1(n_570), .B2(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g901 ( .A(n_67), .Y(n_901) );
INVx1_ASAP7_75t_L g645 ( .A(n_68), .Y(n_645) );
INVx1_ASAP7_75t_L g918 ( .A(n_69), .Y(n_918) );
INVx1_ASAP7_75t_L g613 ( .A(n_70), .Y(n_613) );
OAI222xp33_ASAP7_75t_L g1205 ( .A1(n_71), .A2(n_95), .B1(n_213), .B2(n_377), .C1(n_1206), .C2(n_1207), .Y(n_1205) );
OAI222xp33_ASAP7_75t_L g1251 ( .A1(n_71), .A2(n_95), .B1(n_213), .B2(n_488), .C1(n_587), .C2(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g768 ( .A(n_72), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_73), .A2(n_232), .B1(n_1218), .B2(n_1220), .Y(n_1217) );
AOI22xp33_ASAP7_75t_SL g1243 ( .A1(n_73), .A2(n_120), .B1(n_1244), .B2(n_1245), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_74), .A2(n_120), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
AOI22xp33_ASAP7_75t_SL g1235 ( .A1(n_74), .A2(n_232), .B1(n_1236), .B2(n_1240), .Y(n_1235) );
INVx1_ASAP7_75t_L g747 ( .A(n_75), .Y(n_747) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_76), .A2(n_189), .B1(n_798), .B2(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_76), .A2(n_78), .B1(n_279), .B2(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g341 ( .A(n_77), .Y(n_341) );
OAI211xp5_ASAP7_75t_SL g376 ( .A1(n_77), .A2(n_377), .B(n_382), .C(n_392), .Y(n_376) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_78), .A2(n_152), .B1(n_788), .B2(n_791), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_79), .A2(n_107), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_80), .A2(n_93), .B1(n_1000), .B2(n_1002), .Y(n_1037) );
XOR2x2_ASAP7_75t_L g741 ( .A(n_81), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g640 ( .A(n_82), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g667 ( .A1(n_83), .A2(n_527), .B(n_668), .C(n_672), .Y(n_667) );
INVx1_ASAP7_75t_L g683 ( .A(n_83), .Y(n_683) );
INVx1_ASAP7_75t_L g494 ( .A(n_84), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_85), .A2(n_153), .B1(n_455), .B2(n_750), .Y(n_749) );
OAI22xp33_ASAP7_75t_L g761 ( .A1(n_85), .A2(n_153), .B1(n_373), .B2(n_375), .Y(n_761) );
INVx1_ASAP7_75t_L g718 ( .A(n_87), .Y(n_718) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_88), .Y(n_983) );
AND2x2_ASAP7_75t_L g990 ( .A(n_88), .B(n_981), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_90), .A2(n_158), .B1(n_548), .B2(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_90), .A2(n_158), .B1(n_540), .B2(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g993 ( .A(n_91), .Y(n_993) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_91), .B(n_992), .Y(n_1001) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_92), .A2(n_148), .B1(n_1005), .B2(n_1006), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_96), .Y(n_423) );
INVx1_ASAP7_75t_L g949 ( .A(n_97), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_98), .A2(n_204), .B1(n_1203), .B2(n_1204), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_98), .A2(n_204), .B1(n_355), .B2(n_589), .Y(n_1250) );
INVx2_ASAP7_75t_L g249 ( .A(n_99), .Y(n_249) );
INVx1_ASAP7_75t_L g293 ( .A(n_99), .Y(n_293) );
INVx1_ASAP7_75t_L g575 ( .A(n_100), .Y(n_575) );
INVx1_ASAP7_75t_L g921 ( .A(n_101), .Y(n_921) );
INVx1_ASAP7_75t_L g766 ( .A(n_102), .Y(n_766) );
INVx1_ASAP7_75t_L g534 ( .A(n_103), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_105), .A2(n_215), .B1(n_373), .B2(n_375), .Y(n_372) );
OAI22xp33_ASAP7_75t_SL g884 ( .A1(n_106), .A2(n_110), .B1(n_455), .B2(n_666), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_106), .A2(n_119), .B1(n_387), .B2(n_388), .Y(n_891) );
INVx1_ASAP7_75t_L g1199 ( .A(n_108), .Y(n_1199) );
OAI22xp5_ASAP7_75t_SL g904 ( .A1(n_109), .A2(n_184), .B1(n_373), .B2(n_396), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_111), .A2(n_218), .B1(n_1005), .B2(n_1006), .Y(n_1038) );
INVx1_ASAP7_75t_L g726 ( .A(n_112), .Y(n_726) );
INVx1_ASAP7_75t_L g924 ( .A(n_113), .Y(n_924) );
INVx1_ASAP7_75t_L g962 ( .A(n_115), .Y(n_962) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_116), .A2(n_118), .B1(n_1000), .B2(n_1002), .Y(n_999) );
INVx1_ASAP7_75t_L g775 ( .A(n_117), .Y(n_775) );
INVx1_ASAP7_75t_L g883 ( .A(n_119), .Y(n_883) );
INVx1_ASAP7_75t_L g598 ( .A(n_121), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_123), .A2(n_126), .B1(n_1005), .B2(n_1006), .Y(n_1019) );
AOI222xp33_ASAP7_75t_L g1193 ( .A1(n_123), .A2(n_1194), .B1(n_1254), .B2(n_1258), .C1(n_1262), .C2(n_1264), .Y(n_1193) );
XOR2xp5_ASAP7_75t_L g1195 ( .A(n_123), .B(n_1196), .Y(n_1195) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_124), .Y(n_449) );
INVx1_ASAP7_75t_L g604 ( .A(n_125), .Y(n_604) );
INVx1_ASAP7_75t_L g922 ( .A(n_128), .Y(n_922) );
INVx1_ASAP7_75t_L g948 ( .A(n_129), .Y(n_948) );
BUFx3_ASAP7_75t_L g255 ( .A(n_131), .Y(n_255) );
OAI211xp5_ASAP7_75t_SL g880 ( .A1(n_132), .A2(n_332), .B(n_333), .C(n_881), .Y(n_880) );
OAI211xp5_ASAP7_75t_SL g888 ( .A1(n_132), .A2(n_392), .B(n_889), .C(n_890), .Y(n_888) );
INVx1_ASAP7_75t_L g916 ( .A(n_133), .Y(n_916) );
INVx1_ASAP7_75t_L g711 ( .A(n_134), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g1027 ( .A1(n_135), .A2(n_137), .B1(n_1005), .B2(n_1006), .Y(n_1027) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_136), .Y(n_430) );
INVx1_ASAP7_75t_L g642 ( .A(n_138), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g1030 ( .A1(n_139), .A2(n_203), .B1(n_1000), .B2(n_1002), .Y(n_1030) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_140), .A2(n_231), .B1(n_373), .B2(n_375), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_141), .Y(n_425) );
INVx1_ASAP7_75t_L g537 ( .A(n_142), .Y(n_537) );
OAI211xp5_ASAP7_75t_SL g549 ( .A1(n_142), .A2(n_392), .B(n_550), .C(n_552), .Y(n_549) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_143), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_144), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_145), .A2(n_182), .B1(n_559), .B2(n_578), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_145), .A2(n_182), .B1(n_352), .B2(n_362), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_146), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_147), .A2(n_185), .B1(n_1212), .B2(n_1216), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_147), .A2(n_176), .B1(n_1232), .B2(n_1234), .Y(n_1231) );
XOR2x2_ASAP7_75t_L g894 ( .A(n_148), .B(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g946 ( .A(n_149), .Y(n_946) );
INVx1_ASAP7_75t_L g716 ( .A(n_150), .Y(n_716) );
INVx1_ASAP7_75t_L g941 ( .A(n_151), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_152), .A2(n_189), .B1(n_808), .B2(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g694 ( .A(n_155), .Y(n_694) );
INVx1_ASAP7_75t_L g648 ( .A(n_156), .Y(n_648) );
OA22x2_ASAP7_75t_L g566 ( .A1(n_159), .A2(n_567), .B1(n_630), .B2(n_631), .Y(n_566) );
INVxp67_ASAP7_75t_L g631 ( .A(n_159), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_161), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_162), .A2(n_225), .B1(n_814), .B2(n_819), .Y(n_813) );
INVx1_ASAP7_75t_L g834 ( .A(n_163), .Y(n_834) );
INVx1_ASAP7_75t_L g502 ( .A(n_164), .Y(n_502) );
INVx1_ASAP7_75t_L g925 ( .A(n_165), .Y(n_925) );
INVx1_ASAP7_75t_L g595 ( .A(n_166), .Y(n_595) );
OAI211xp5_ASAP7_75t_SL g692 ( .A1(n_167), .A2(n_392), .B(n_680), .C(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g703 ( .A(n_167), .Y(n_703) );
INVx1_ASAP7_75t_L g963 ( .A(n_168), .Y(n_963) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_169), .Y(n_288) );
OAI211xp5_ASAP7_75t_L g571 ( .A1(n_170), .A2(n_462), .B(n_572), .C(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g585 ( .A(n_170), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_171), .Y(n_417) );
OAI211xp5_ASAP7_75t_L g331 ( .A1(n_172), .A2(n_332), .B(n_333), .C(n_340), .Y(n_331) );
INVx1_ASAP7_75t_L g391 ( .A(n_172), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g696 ( .A1(n_173), .A2(n_223), .B1(n_570), .B2(n_685), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_173), .A2(n_223), .B1(n_539), .B2(n_705), .Y(n_704) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_174), .Y(n_305) );
INVx1_ASAP7_75t_L g835 ( .A(n_175), .Y(n_835) );
INVx1_ASAP7_75t_L g496 ( .A(n_177), .Y(n_496) );
INVx1_ASAP7_75t_L g942 ( .A(n_178), .Y(n_942) );
INVx1_ASAP7_75t_L g451 ( .A(n_180), .Y(n_451) );
OAI211xp5_ASAP7_75t_L g458 ( .A1(n_180), .A2(n_459), .B(n_462), .C(n_463), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_181), .Y(n_258) );
INVx1_ASAP7_75t_L g900 ( .A(n_183), .Y(n_900) );
OAI211xp5_ASAP7_75t_SL g526 ( .A1(n_187), .A2(n_527), .B(n_530), .C(n_533), .Y(n_526) );
INVx1_ASAP7_75t_L g555 ( .A(n_187), .Y(n_555) );
INVx1_ASAP7_75t_L g772 ( .A(n_188), .Y(n_772) );
INVx1_ASAP7_75t_L g938 ( .A(n_190), .Y(n_938) );
INVx1_ASAP7_75t_L g671 ( .A(n_191), .Y(n_671) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_191), .A2(n_392), .B(n_680), .C(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g919 ( .A(n_192), .Y(n_919) );
INVx1_ASAP7_75t_L g945 ( .A(n_193), .Y(n_945) );
INVx1_ASAP7_75t_L g830 ( .A(n_194), .Y(n_830) );
INVx1_ASAP7_75t_L g612 ( .A(n_195), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g868 ( .A(n_196), .Y(n_868) );
INVx1_ASAP7_75t_L g770 ( .A(n_197), .Y(n_770) );
XOR2xp5_ASAP7_75t_L g851 ( .A(n_198), .B(n_852), .Y(n_851) );
BUFx3_ASAP7_75t_L g299 ( .A(n_201), .Y(n_299) );
INVx1_ASAP7_75t_L g361 ( .A(n_201), .Y(n_361) );
INVx1_ASAP7_75t_L g669 ( .A(n_202), .Y(n_669) );
XOR2x2_ASAP7_75t_L g688 ( .A(n_205), .B(n_689), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_206), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_207), .Y(n_860) );
INVx1_ASAP7_75t_L g607 ( .A(n_208), .Y(n_607) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_209), .A2(n_333), .B(n_446), .C(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g465 ( .A(n_209), .Y(n_465) );
INVx1_ASAP7_75t_L g602 ( .A(n_210), .Y(n_602) );
INVx1_ASAP7_75t_L g723 ( .A(n_211), .Y(n_723) );
INVx1_ASAP7_75t_L g765 ( .A(n_212), .Y(n_765) );
INVx1_ASAP7_75t_L g965 ( .A(n_214), .Y(n_965) );
OAI211xp5_ASAP7_75t_L g744 ( .A1(n_216), .A2(n_333), .B(n_745), .C(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g757 ( .A(n_216), .Y(n_757) );
INVx1_ASAP7_75t_L g247 ( .A(n_217), .Y(n_247) );
INVx2_ASAP7_75t_L g291 ( .A(n_217), .Y(n_291) );
INVx1_ASAP7_75t_L g521 ( .A(n_217), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_219), .Y(n_280) );
INVx1_ASAP7_75t_L g477 ( .A(n_220), .Y(n_477) );
INVx1_ASAP7_75t_L g651 ( .A(n_221), .Y(n_651) );
INVx1_ASAP7_75t_L g483 ( .A(n_222), .Y(n_483) );
INVx1_ASAP7_75t_L g725 ( .A(n_224), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g407 ( .A(n_226), .B(n_408), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g452 ( .A1(n_227), .A2(n_231), .B1(n_352), .B2(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g695 ( .A(n_228), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_228), .A2(n_530), .B(n_699), .C(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g1200 ( .A(n_229), .Y(n_1200) );
XNOR2xp5_ASAP7_75t_L g1259 ( .A(n_230), .B(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g647 ( .A(n_233), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_978), .B(n_987), .Y(n_234) );
XNOR2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_632), .Y(n_235) );
XOR2x1_ASAP7_75t_L g236 ( .A(n_237), .B(n_468), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_405), .B1(n_406), .B2(n_467), .Y(n_237) );
INVx1_ASAP7_75t_L g467 ( .A(n_238), .Y(n_467) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND3xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_330), .C(n_371), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g241 ( .A(n_242), .B(n_295), .Y(n_241) );
OAI33xp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_251), .A3(n_265), .B1(n_277), .B2(n_285), .B3(n_289), .Y(n_242) );
OAI33xp33_ASAP7_75t_L g432 ( .A1(n_243), .A2(n_289), .A3(n_433), .B1(n_436), .B2(n_440), .B3(n_443), .Y(n_432) );
OAI33xp33_ASAP7_75t_L g763 ( .A1(n_243), .A2(n_289), .A3(n_764), .B1(n_767), .B2(n_771), .B3(n_774), .Y(n_763) );
OAI33xp33_ASAP7_75t_L g854 ( .A1(n_243), .A2(n_289), .A3(n_855), .B1(n_859), .B2(n_862), .B3(n_866), .Y(n_854) );
OAI33xp33_ASAP7_75t_L g926 ( .A1(n_243), .A2(n_289), .A3(n_927), .B1(n_928), .B2(n_929), .B3(n_930), .Y(n_926) );
BUFx4f_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
BUFx2_ASAP7_75t_L g507 ( .A(n_244), .Y(n_507) );
BUFx4f_ASAP7_75t_L g653 ( .A(n_244), .Y(n_653) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_248), .Y(n_244) );
AND2x2_ASAP7_75t_SL g327 ( .A(n_245), .B(n_328), .Y(n_327) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_245), .Y(n_404) );
INVx1_ASAP7_75t_L g500 ( .A(n_245), .Y(n_500) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
BUFx2_ASAP7_75t_L g370 ( .A(n_246), .Y(n_370) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp33_ASAP7_75t_SL g248 ( .A(n_249), .B(n_250), .Y(n_248) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_249), .Y(n_402) );
AND3x4_ASAP7_75t_L g811 ( .A(n_249), .B(n_380), .C(n_812), .Y(n_811) );
INVx3_ASAP7_75t_L g294 ( .A(n_250), .Y(n_294) );
BUFx3_ASAP7_75t_L g380 ( .A(n_250), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B1(n_258), .B2(n_259), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_252), .A2(n_286), .B1(n_301), .B2(n_307), .Y(n_300) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_253), .A2(n_286), .B1(n_287), .B2(n_288), .Y(n_285) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_253), .A2(n_259), .B1(n_765), .B2(n_766), .Y(n_764) );
OAI22xp33_ASAP7_75t_L g774 ( .A1(n_253), .A2(n_287), .B1(n_775), .B2(n_776), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_253), .A2(n_856), .B1(n_857), .B2(n_858), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_253), .A2(n_287), .B1(n_867), .B2(n_868), .Y(n_866) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_253), .A2(n_916), .B1(n_922), .B2(n_931), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g951 ( .A1(n_253), .A2(n_857), .B1(n_941), .B2(n_948), .Y(n_951) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_253), .A2(n_287), .B1(n_942), .B2(n_949), .Y(n_957) );
BUFx4f_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x4_ASAP7_75t_L g373 ( .A(n_254), .B(n_374), .Y(n_373) );
OR2x4_ASAP7_75t_L g396 ( .A(n_254), .B(n_294), .Y(n_396) );
INVx2_ASAP7_75t_L g435 ( .A(n_254), .Y(n_435) );
BUFx3_ASAP7_75t_L g509 ( .A(n_254), .Y(n_509) );
BUFx3_ASAP7_75t_L g618 ( .A(n_254), .Y(n_618) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_255), .Y(n_264) );
INVx2_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_255), .B(n_263), .Y(n_275) );
AND2x4_ASAP7_75t_L g394 ( .A(n_255), .B(n_386), .Y(n_394) );
INVx1_ASAP7_75t_L g818 ( .A(n_256), .Y(n_818) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVxp67_ASAP7_75t_L g270 ( .A(n_257), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_258), .A2(n_288), .B1(n_313), .B2(n_317), .Y(n_321) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_259), .A2(n_413), .B1(n_423), .B2(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g573 ( .A(n_259), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_259), .A2(n_598), .B1(n_607), .B2(n_616), .Y(n_629) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_260), .Y(n_510) );
INVx4_ASAP7_75t_L g681 ( .A(n_260), .Y(n_681) );
INVx3_ASAP7_75t_L g714 ( .A(n_260), .Y(n_714) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx3_ASAP7_75t_L g287 ( .A(n_261), .Y(n_287) );
BUFx2_ASAP7_75t_L g461 ( .A(n_261), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
BUFx2_ASAP7_75t_L g390 ( .A(n_262), .Y(n_390) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g386 ( .A(n_263), .Y(n_386) );
BUFx2_ASAP7_75t_L g381 ( .A(n_264), .Y(n_381) );
INVx2_ASAP7_75t_L g388 ( .A(n_264), .Y(n_388) );
AND2x4_ASAP7_75t_L g810 ( .A(n_264), .B(n_385), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B1(n_272), .B2(n_276), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_266), .A2(n_280), .B1(n_313), .B2(n_317), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_267), .A2(n_281), .B1(n_772), .B2(n_773), .Y(n_771) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g769 ( .A(n_268), .Y(n_769) );
BUFx8_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_269), .Y(n_279) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_269), .Y(n_399) );
INVx2_ASAP7_75t_L g627 ( .A(n_269), .Y(n_627) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x4_ASAP7_75t_L g817 ( .A(n_271), .B(n_818), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_272), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_767) );
OAI22xp33_ASAP7_75t_SL g952 ( .A1(n_272), .A2(n_660), .B1(n_938), .B2(n_945), .Y(n_952) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x6_ASAP7_75t_L g375 ( .A(n_274), .B(n_294), .Y(n_375) );
BUFx3_ASAP7_75t_L g514 ( .A(n_274), .Y(n_514) );
BUFx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g283 ( .A(n_275), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_276), .A2(n_284), .B1(n_307), .B2(n_323), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B1(n_281), .B2(n_284), .Y(n_277) );
INVx2_ASAP7_75t_L g721 ( .A(n_278), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_278), .A2(n_438), .B1(n_918), .B2(n_924), .Y(n_928) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_SL g441 ( .A(n_279), .Y(n_441) );
INVx5_ASAP7_75t_L g660 ( .A(n_279), .Y(n_660) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_279), .Y(n_808) );
BUFx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g955 ( .A(n_282), .Y(n_955) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_283), .Y(n_439) );
OAI22xp33_ASAP7_75t_L g443 ( .A1(n_287), .A2(n_415), .B1(n_425), .B2(n_434), .Y(n_443) );
INVx2_ASAP7_75t_L g658 ( .A(n_287), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_287), .A2(n_434), .B1(n_915), .B2(n_921), .Y(n_927) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
AND2x4_ASAP7_75t_L g297 ( .A(n_290), .B(n_298), .Y(n_297) );
OR2x6_ASAP7_75t_L g956 ( .A(n_290), .B(n_292), .Y(n_956) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g812 ( .A(n_291), .Y(n_812) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND3x1_ASAP7_75t_L g519 ( .A(n_293), .B(n_294), .C(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g374 ( .A(n_294), .Y(n_374) );
AND2x4_ASAP7_75t_L g393 ( .A(n_294), .B(n_394), .Y(n_393) );
OAI33xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .A3(n_312), .B1(n_321), .B2(n_322), .B3(n_326), .Y(n_295) );
OAI33xp33_ASAP7_75t_L g777 ( .A1(n_296), .A2(n_326), .A3(n_778), .B1(n_780), .B2(n_781), .B3(n_782), .Y(n_777) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g411 ( .A(n_297), .Y(n_411) );
INVx2_ASAP7_75t_L g600 ( .A(n_297), .Y(n_600) );
INVx4_ASAP7_75t_L g801 ( .A(n_297), .Y(n_801) );
AND2x4_ASAP7_75t_L g328 ( .A(n_299), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g336 ( .A(n_299), .Y(n_336) );
BUFx2_ASAP7_75t_L g343 ( .A(n_299), .Y(n_343) );
AND2x4_ASAP7_75t_L g348 ( .A(n_299), .B(n_349), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_301), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_301), .A2(n_427), .B1(n_428), .B2(n_430), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_301), .A2(n_765), .B1(n_775), .B2(n_779), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_301), .A2(n_428), .B1(n_915), .B2(n_916), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_301), .A2(n_414), .B1(n_924), .B2(n_925), .Y(n_923) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_301), .A2(n_504), .B1(n_941), .B2(n_942), .Y(n_940) );
INVx4_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_302), .Y(n_597) );
INVx3_ASAP7_75t_L g641 ( .A(n_302), .Y(n_641) );
BUFx4f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g325 ( .A(n_303), .Y(n_325) );
INVx3_ASAP7_75t_L g354 ( .A(n_303), .Y(n_354) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx2_ASAP7_75t_L g311 ( .A(n_305), .Y(n_311) );
INVx2_ASAP7_75t_L g316 ( .A(n_305), .Y(n_316) );
NAND2x1_ASAP7_75t_L g320 ( .A(n_305), .B(n_306), .Y(n_320) );
AND2x2_ASAP7_75t_L g339 ( .A(n_305), .B(n_306), .Y(n_339) );
INVx1_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
AND2x2_ASAP7_75t_L g364 ( .A(n_305), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_306), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g315 ( .A(n_306), .B(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g344 ( .A(n_306), .Y(n_344) );
INVx2_ASAP7_75t_L g365 ( .A(n_306), .Y(n_365) );
INVx1_ASAP7_75t_L g797 ( .A(n_306), .Y(n_797) );
AND2x2_ASAP7_75t_L g799 ( .A(n_306), .B(n_311), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_307), .A2(n_323), .B1(n_770), .B2(n_773), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_307), .A2(n_861), .B1(n_864), .B2(n_871), .Y(n_877) );
INVx4_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_SL g414 ( .A(n_308), .Y(n_414) );
INVx2_ASAP7_75t_L g429 ( .A(n_308), .Y(n_429) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_308), .Y(n_481) );
INVx1_ASAP7_75t_L g504 ( .A(n_308), .Y(n_504) );
INVx1_ASAP7_75t_L g779 ( .A(n_308), .Y(n_779) );
INVx8_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g357 ( .A(n_309), .B(n_343), .Y(n_357) );
OR2x2_ASAP7_75t_L g750 ( .A(n_309), .B(n_335), .Y(n_750) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_313), .A2(n_317), .B1(n_768), .B2(n_772), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_313), .A2(n_421), .B1(n_766), .B2(n_776), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_313), .A2(n_860), .B1(n_863), .B2(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_313), .A2(n_424), .B1(n_938), .B2(n_939), .Y(n_937) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g603 ( .A(n_314), .Y(n_603) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g419 ( .A(n_315), .Y(n_419) );
BUFx2_ASAP7_75t_L g486 ( .A(n_315), .Y(n_486) );
BUFx3_ASAP7_75t_L g875 ( .A(n_315), .Y(n_875) );
AND2x2_ASAP7_75t_L g796 ( .A(n_316), .B(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g446 ( .A(n_318), .Y(n_446) );
INVx1_ASAP7_75t_L g582 ( .A(n_318), .Y(n_582) );
INVx2_ASAP7_75t_L g734 ( .A(n_318), .Y(n_734) );
INVx2_ASAP7_75t_L g876 ( .A(n_318), .Y(n_876) );
INVx4_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx4f_ASAP7_75t_L g332 ( .A(n_319), .Y(n_332) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_319), .Y(n_424) );
BUFx4f_ASAP7_75t_L g529 ( .A(n_319), .Y(n_529) );
BUFx4f_ASAP7_75t_L g873 ( .A(n_319), .Y(n_873) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g421 ( .A(n_320), .Y(n_421) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x6_ASAP7_75t_L g359 ( .A(n_325), .B(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g455 ( .A(n_325), .B(n_360), .Y(n_455) );
OR2x6_ASAP7_75t_L g543 ( .A(n_325), .B(n_353), .Y(n_543) );
OAI33xp33_ASAP7_75t_L g869 ( .A1(n_326), .A2(n_411), .A3(n_870), .B1(n_872), .B2(n_874), .B3(n_877), .Y(n_869) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g431 ( .A(n_327), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_327), .B(n_803), .C(n_805), .Y(n_802) );
AND2x4_ASAP7_75t_L g498 ( .A(n_328), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g368 ( .A(n_329), .Y(n_368) );
OAI31xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_351), .A3(n_358), .B(n_366), .Y(n_330) );
NAND3xp33_ASAP7_75t_L g828 ( .A(n_333), .B(n_829), .C(n_833), .Y(n_828) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_L g448 ( .A(n_335), .B(n_344), .Y(n_448) );
AND2x2_ASAP7_75t_L g531 ( .A(n_335), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVxp67_ASAP7_75t_L g353 ( .A(n_336), .Y(n_353) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g1241 ( .A(n_338), .Y(n_1241) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_339), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_345), .B2(n_346), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_342), .A2(n_575), .B1(n_585), .B2(n_586), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_342), .A2(n_670), .B1(n_694), .B2(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_342), .A2(n_450), .B1(n_962), .B2(n_963), .Y(n_961) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x4_ASAP7_75t_L g536 ( .A(n_343), .B(n_344), .Y(n_536) );
AND2x2_ASAP7_75t_L g831 ( .A(n_343), .B(n_795), .Y(n_831) );
AOI32xp33_ASAP7_75t_L g382 ( .A1(n_345), .A2(n_383), .A3(n_387), .B1(n_389), .B2(n_391), .Y(n_382) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g450 ( .A(n_348), .Y(n_450) );
INVx2_ASAP7_75t_L g587 ( .A(n_348), .Y(n_587) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x6_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
BUFx3_ASAP7_75t_L g478 ( .A(n_354), .Y(n_478) );
INVx2_ASAP7_75t_SL g611 ( .A(n_354), .Y(n_611) );
BUFx3_ASAP7_75t_L g871 ( .A(n_354), .Y(n_871) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g453 ( .A(n_357), .Y(n_453) );
INVx2_ASAP7_75t_L g541 ( .A(n_357), .Y(n_541) );
BUFx2_ASAP7_75t_L g539 ( .A(n_359), .Y(n_539) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_359), .Y(n_589) );
AND2x4_ASAP7_75t_L g363 ( .A(n_360), .B(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_363), .Y(n_362) );
INVx4_ASAP7_75t_L g666 ( .A(n_363), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_363), .A2(n_986), .B1(n_1199), .B2(n_1200), .Y(n_1248) );
BUFx3_ASAP7_75t_L g790 ( .A(n_364), .Y(n_790) );
INVx2_ASAP7_75t_L g1239 ( .A(n_364), .Y(n_1239) );
OAI31xp33_ASAP7_75t_L g444 ( .A1(n_366), .A2(n_445), .A3(n_452), .B(n_454), .Y(n_444) );
OAI31xp33_ASAP7_75t_L g958 ( .A1(n_366), .A2(n_959), .A3(n_960), .B(n_966), .Y(n_958) );
BUFx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g544 ( .A(n_367), .Y(n_544) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_367), .Y(n_591) );
OAI31xp33_ASAP7_75t_L g878 ( .A1(n_367), .A2(n_879), .A3(n_880), .B(n_884), .Y(n_878) );
OAI31xp33_ASAP7_75t_L g896 ( .A1(n_367), .A2(n_897), .A3(n_898), .B(n_902), .Y(n_896) );
INVx1_ASAP7_75t_L g1253 ( .A(n_367), .Y(n_1253) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g985 ( .A(n_368), .Y(n_985) );
NOR2xp33_ASAP7_75t_L g1256 ( .A(n_368), .B(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI31xp33_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_376), .A3(n_395), .B(n_400), .Y(n_371) );
BUFx2_ASAP7_75t_L g547 ( .A(n_373), .Y(n_547) );
BUFx3_ASAP7_75t_L g570 ( .A(n_373), .Y(n_570) );
INVx2_ASAP7_75t_SL g847 ( .A(n_373), .Y(n_847) );
BUFx2_ASAP7_75t_L g1203 ( .A(n_373), .Y(n_1203) );
AND2x2_ASAP7_75t_L g398 ( .A(n_374), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g562 ( .A(n_374), .B(n_399), .Y(n_562) );
BUFx3_ASAP7_75t_L g548 ( .A(n_375), .Y(n_548) );
INVx1_ASAP7_75t_L g686 ( .A(n_375), .Y(n_686) );
INVx2_ASAP7_75t_L g848 ( .A(n_375), .Y(n_848) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_378), .A2(n_557), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_378), .A2(n_389), .B1(n_747), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_378), .A2(n_557), .B1(n_962), .B2(n_965), .Y(n_971) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
AND2x2_ASAP7_75t_L g389 ( .A(n_379), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g464 ( .A(n_379), .B(n_381), .Y(n_464) );
AND2x2_ASAP7_75t_L g554 ( .A(n_379), .B(n_381), .Y(n_554) );
AND2x4_ASAP7_75t_L g557 ( .A(n_379), .B(n_390), .Y(n_557) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g383 ( .A(n_380), .B(n_384), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_383), .A2(n_464), .B1(n_882), .B2(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_389), .A2(n_449), .B1(n_464), .B2(n_465), .Y(n_463) );
INVxp67_ASAP7_75t_L g889 ( .A(n_389), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_389), .A2(n_464), .B1(n_900), .B2(n_909), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_392), .B(n_843), .C(n_846), .Y(n_842) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_392), .B(n_971), .C(n_972), .Y(n_970) );
CKINVDCx8_ASAP7_75t_R g392 ( .A(n_393), .Y(n_392) );
CKINVDCx8_ASAP7_75t_R g462 ( .A(n_393), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g1201 ( .A(n_393), .B(n_1202), .C(n_1205), .Y(n_1201) );
BUFx3_ASAP7_75t_L g760 ( .A(n_394), .Y(n_760) );
INVx2_ASAP7_75t_L g820 ( .A(n_394), .Y(n_820) );
BUFx2_ASAP7_75t_L g844 ( .A(n_394), .Y(n_844) );
BUFx2_ASAP7_75t_L g907 ( .A(n_394), .Y(n_907) );
BUFx2_ASAP7_75t_L g1224 ( .A(n_394), .Y(n_1224) );
INVx1_ASAP7_75t_L g560 ( .A(n_396), .Y(n_560) );
INVx2_ASAP7_75t_SL g677 ( .A(n_396), .Y(n_677) );
INVx2_ASAP7_75t_SL g841 ( .A(n_396), .Y(n_841) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g437 ( .A(n_399), .Y(n_437) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_399), .Y(n_513) );
INVx2_ASAP7_75t_L g516 ( .A(n_399), .Y(n_516) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_399), .Y(n_622) );
OAI31xp33_ASAP7_75t_SL g456 ( .A1(n_400), .A2(n_457), .A3(n_458), .B(n_466), .Y(n_456) );
OAI31xp33_ASAP7_75t_L g752 ( .A1(n_400), .A2(n_753), .A3(n_755), .B(n_761), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g838 ( .A1(n_400), .A2(n_839), .B(n_842), .Y(n_838) );
OAI31xp33_ASAP7_75t_SL g885 ( .A1(n_400), .A2(n_886), .A3(n_887), .B(n_888), .Y(n_885) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
AND2x2_ASAP7_75t_SL g564 ( .A(n_401), .B(n_403), .Y(n_564) );
AND2x4_ASAP7_75t_L g579 ( .A(n_401), .B(n_403), .Y(n_579) );
AND2x2_ASAP7_75t_L g911 ( .A(n_401), .B(n_403), .Y(n_911) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AND3x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_444), .C(n_456), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_432), .Y(n_409) );
OAI33xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .A3(n_416), .B1(n_422), .B2(n_426), .B3(n_431), .Y(n_410) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_411), .Y(n_475) );
OAI33xp33_ASAP7_75t_L g913 ( .A1(n_411), .A2(n_431), .A3(n_914), .B1(n_917), .B2(n_920), .B3(n_923), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_420), .B2(n_421), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_417), .A2(n_427), .B1(n_437), .B2(n_438), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_418), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_418), .A2(n_424), .B1(n_918), .B2(n_919), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_418), .A2(n_873), .B1(n_921), .B2(n_922), .Y(n_920) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g493 ( .A(n_419), .Y(n_493) );
BUFx2_ASAP7_75t_L g733 ( .A(n_419), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_420), .A2(n_430), .B1(n_441), .B2(n_442), .Y(n_440) );
INVx2_ASAP7_75t_SL g489 ( .A(n_421), .Y(n_489) );
BUFx2_ASAP7_75t_SL g495 ( .A(n_421), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_421), .A2(n_493), .B1(n_644), .B2(n_645), .Y(n_643) );
BUFx3_ASAP7_75t_L g701 ( .A(n_421), .Y(n_701) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_424), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_428), .A2(n_856), .B1(n_867), .B2(n_871), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_428), .A2(n_871), .B1(n_945), .B2(n_946), .Y(n_944) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI33xp33_ASAP7_75t_L g936 ( .A1(n_431), .A2(n_937), .A3(n_940), .B1(n_943), .B2(n_944), .B3(n_947), .Y(n_936) );
INVx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_437), .A2(n_438), .B1(n_860), .B2(n_861), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_437), .A2(n_865), .B1(n_919), .B2(n_925), .Y(n_929) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx3_ASAP7_75t_L g442 ( .A(n_439), .Y(n_442) );
CKINVDCx8_ASAP7_75t_R g623 ( .A(n_439), .Y(n_623) );
INVx3_ASAP7_75t_L g865 ( .A(n_439), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_441), .A2(n_514), .B1(n_645), .B2(n_651), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_441), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_446), .A2(n_712), .B1(n_726), .B2(n_732), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_450), .A2(n_534), .B1(n_535), .B2(n_537), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_450), .A2(n_536), .B1(n_747), .B2(n_748), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g833 ( .A1(n_450), .A2(n_536), .B1(n_791), .B2(n_834), .C1(n_835), .C2(n_836), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_450), .A2(n_536), .B1(n_882), .B2(n_883), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_450), .A2(n_536), .B1(n_900), .B2(n_901), .Y(n_899) );
INVx2_ASAP7_75t_SL g706 ( .A(n_453), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_459), .A2(n_642), .B1(n_648), .B2(n_655), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g724 ( .A1(n_459), .A2(n_509), .B1(n_725), .B2(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g524 ( .A(n_461), .Y(n_524) );
INVx1_ASAP7_75t_L g551 ( .A(n_461), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_462), .B(n_756), .C(n_758), .Y(n_755) );
NAND3xp33_ASAP7_75t_SL g905 ( .A(n_462), .B(n_906), .C(n_908), .Y(n_905) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
OA22x2_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_565), .B2(n_566), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_525), .C(n_545), .Y(n_472) );
NOR2xp33_ASAP7_75t_SL g473 ( .A(n_474), .B(n_506), .Y(n_473) );
OAI33xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .A3(n_482), .B1(n_490), .B2(n_497), .B3(n_501), .Y(n_474) );
INVx1_ASAP7_75t_L g1230 ( .A(n_475), .Y(n_1230) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_476) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_477), .A2(n_494), .B1(n_509), .B2(n_510), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_478), .A2(n_502), .B1(n_503), .B2(n_505), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_478), .A2(n_480), .B1(n_650), .B2(n_651), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_479), .A2(n_496), .B1(n_509), .B2(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g639 ( .A1(n_480), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_480), .A2(n_711), .B1(n_725), .B2(n_729), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_480), .A2(n_718), .B1(n_723), .B2(n_729), .Y(n_736) );
INVx6_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx5_ASAP7_75t_L g599 ( .A(n_481), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_487), .B2(n_488), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_483), .A2(n_502), .B1(n_512), .B2(n_514), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_484), .A2(n_495), .B1(n_647), .B2(n_648), .Y(n_646) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx4_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_487), .A2(n_505), .B1(n_514), .B2(n_516), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_488), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_601) );
INVx5_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI33xp33_ASAP7_75t_L g638 ( .A1(n_497), .A2(n_600), .A3(n_639), .B1(n_643), .B2(n_646), .B3(n_649), .Y(n_638) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_498), .Y(n_608) );
AOI33xp33_ASAP7_75t_L g1229 ( .A1(n_498), .A2(n_1230), .A3(n_1231), .B1(n_1235), .B2(n_1242), .B3(n_1243), .Y(n_1229) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OAI33xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .A3(n_511), .B1(n_515), .B2(n_517), .B3(n_522), .Y(n_506) );
OAI33xp33_ASAP7_75t_L g614 ( .A1(n_507), .A2(n_615), .A3(n_620), .B1(n_624), .B2(n_628), .B3(n_629), .Y(n_614) );
OAI33xp33_ASAP7_75t_L g709 ( .A1(n_507), .A2(n_517), .A3(n_710), .B1(n_715), .B2(n_719), .B3(n_724), .Y(n_709) );
OAI33xp33_ASAP7_75t_L g950 ( .A1(n_507), .A2(n_951), .A3(n_952), .B1(n_953), .B2(n_956), .B3(n_957), .Y(n_950) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_509), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_514), .A2(n_604), .B1(n_613), .B2(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_514), .A2(n_720), .B1(n_722), .B2(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g1228 ( .A(n_517), .Y(n_1228) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g628 ( .A(n_518), .Y(n_628) );
INVx2_ASAP7_75t_L g662 ( .A(n_518), .Y(n_662) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx3_ASAP7_75t_L g825 ( .A(n_519), .Y(n_825) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
OAI31xp33_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_538), .A3(n_542), .B(n_544), .Y(n_525) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_529), .A2(n_603), .B1(n_606), .B2(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g583 ( .A(n_531), .Y(n_583) );
INVx1_ASAP7_75t_L g672 ( .A(n_531), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g1249 ( .A(n_531), .B(n_1250), .C(n_1251), .Y(n_1249) );
BUFx3_ASAP7_75t_L g791 ( .A(n_532), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_534), .A2(n_553), .B1(n_555), .B2(n_556), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_535), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g1252 ( .A(n_536), .Y(n_1252) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_541), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
INVx1_ASAP7_75t_L g967 ( .A(n_541), .Y(n_967) );
INVx3_ASAP7_75t_L g986 ( .A(n_543), .Y(n_986) );
OAI31xp33_ASAP7_75t_L g664 ( .A1(n_544), .A2(n_665), .A3(n_667), .B(n_673), .Y(n_664) );
OAI31xp33_ASAP7_75t_L g697 ( .A1(n_544), .A2(n_698), .A3(n_704), .B(n_707), .Y(n_697) );
OAI31xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_549), .A3(n_558), .B(n_563), .Y(n_545) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g619 ( .A(n_551), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_553), .A2(n_556), .B1(n_669), .B2(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_553), .A2(n_556), .B1(n_694), .B2(n_695), .Y(n_693) );
BUFx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g845 ( .A(n_554), .Y(n_845) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI222xp33_ASAP7_75t_L g843 ( .A1(n_557), .A2(n_834), .B1(n_835), .B2(n_836), .C1(n_844), .C2(n_845), .Y(n_843) );
INVx1_ASAP7_75t_L g1207 ( .A(n_557), .Y(n_1207) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g578 ( .A(n_562), .Y(n_578) );
INVx1_ASAP7_75t_L g678 ( .A(n_562), .Y(n_678) );
INVx1_ASAP7_75t_L g754 ( .A(n_562), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_562), .A2(n_841), .B1(n_1199), .B2(n_1200), .Y(n_1198) );
OAI31xp33_ASAP7_75t_L g674 ( .A1(n_563), .A2(n_675), .A3(n_679), .B(n_684), .Y(n_674) );
OAI31xp33_ASAP7_75t_L g690 ( .A1(n_563), .A2(n_691), .A3(n_692), .B(n_696), .Y(n_690) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g630 ( .A(n_567), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_580), .C(n_592), .Y(n_567) );
OAI31xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_571), .A3(n_577), .B(n_579), .Y(n_568) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
CKINVDCx14_ASAP7_75t_R g1208 ( .A(n_579), .Y(n_1208) );
OAI31xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_588), .A3(n_590), .B(n_591), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g960 ( .A(n_583), .B(n_961), .C(n_964), .Y(n_960) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g670 ( .A(n_587), .Y(n_670) );
OAI31xp33_ASAP7_75t_SL g743 ( .A1(n_591), .A2(n_744), .A3(n_749), .B(n_751), .Y(n_743) );
OAI21xp5_ASAP7_75t_L g827 ( .A1(n_591), .A2(n_828), .B(n_837), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_614), .Y(n_592) );
OAI33xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_600), .A3(n_601), .B1(n_605), .B2(n_608), .B3(n_609), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_598), .B2(n_599), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_595), .A2(n_606), .B1(n_616), .B2(n_619), .Y(n_615) );
INVx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_599), .A2(n_610), .B1(n_612), .B2(n_613), .Y(n_609) );
OAI33xp33_ASAP7_75t_L g727 ( .A1(n_600), .A2(n_608), .A3(n_728), .B1(n_731), .B2(n_735), .B3(n_736), .Y(n_727) );
OAI22xp33_ASAP7_75t_L g620 ( .A1(n_602), .A2(n_612), .B1(n_621), .B2(n_623), .Y(n_620) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_618), .Y(n_656) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_623), .A2(n_644), .B1(n_650), .B2(n_660), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_623), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g1219 ( .A(n_627), .Y(n_1219) );
INVx1_ASAP7_75t_L g1226 ( .A(n_627), .Y(n_1226) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_738), .B1(n_976), .B2(n_977), .Y(n_632) );
OA21x2_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_687), .B(n_737), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g976 ( .A1(n_634), .A2(n_687), .B(n_737), .Y(n_976) );
INVx2_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g737 ( .A(n_635), .B(n_688), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_664), .C(n_674), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_652), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_640), .A2(n_647), .B1(n_655), .B2(n_657), .Y(n_654) );
INVx2_ASAP7_75t_SL g730 ( .A(n_641), .Y(n_730) );
OAI33xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .A3(n_659), .B1(n_661), .B2(n_662), .B3(n_663), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx3_ASAP7_75t_L g717 ( .A(n_660), .Y(n_717) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g931 ( .A(n_681), .Y(n_931) );
INVx1_ASAP7_75t_L g1206 ( .A(n_681), .Y(n_1206) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_697), .C(n_708), .Y(n_689) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_727), .Y(n_708) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_L g857 ( .A(n_714), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_716), .A2(n_722), .B1(n_732), .B2(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx4_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g977 ( .A(n_738), .Y(n_977) );
XNOR2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_849), .Y(n_738) );
INVx2_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
XNOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_783), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_752), .C(n_762), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_748), .B(n_759), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_777), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_769), .A2(n_939), .B1(n_946), .B2(n_954), .Y(n_953) );
NAND3xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_827), .C(n_838), .Y(n_784) );
AND4x1_ASAP7_75t_L g785 ( .A(n_786), .B(n_802), .C(n_806), .D(n_821), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_792), .C(n_800), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_791), .B(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_795), .Y(n_804) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx3_ASAP7_75t_L g1233 ( .A(n_796), .Y(n_1233) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_798), .Y(n_1234) );
BUFx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g1246 ( .A(n_799), .Y(n_1246) );
INVx1_ASAP7_75t_L g943 ( .A(n_800), .Y(n_943) );
INVx2_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
NAND3xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_811), .C(n_813), .Y(n_806) );
BUFx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx12f_ASAP7_75t_L g823 ( .A(n_810), .Y(n_823) );
INVx5_ASAP7_75t_L g1221 ( .A(n_810), .Y(n_1221) );
BUFx3_ASAP7_75t_L g1210 ( .A(n_811), .Y(n_1210) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
BUFx3_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
BUFx3_ASAP7_75t_L g1215 ( .A(n_817), .Y(n_1215) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g1216 ( .A(n_820), .Y(n_1216) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .C(n_826), .Y(n_821) );
BUFx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_830), .A2(n_832), .B1(n_847), .B2(n_848), .Y(n_846) );
INVx2_ASAP7_75t_SL g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g1204 ( .A(n_848), .Y(n_1204) );
XNOR2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_892), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_878), .C(n_885), .Y(n_852) );
NOR2xp33_ASAP7_75t_SL g853 ( .A(n_854), .B(n_869), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_858), .A2(n_868), .B1(n_875), .B2(n_876), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_873), .A2(n_875), .B1(n_948), .B2(n_949), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .B1(n_932), .B2(n_933), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
NAND3xp33_ASAP7_75t_SL g895 ( .A(n_896), .B(n_903), .C(n_912), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_901), .B(n_907), .Y(n_906) );
OAI31xp33_ASAP7_75t_SL g903 ( .A1(n_904), .A2(n_905), .A3(n_910), .B(n_911), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_907), .B(n_963), .Y(n_972) );
OAI31xp33_ASAP7_75t_L g968 ( .A1(n_911), .A2(n_969), .A3(n_970), .B(n_973), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_913), .B(n_926), .Y(n_912) );
INVx3_ASAP7_75t_SL g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g975 ( .A(n_934), .Y(n_975) );
NAND3xp33_ASAP7_75t_L g934 ( .A(n_935), .B(n_958), .C(n_968), .Y(n_934) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_936), .B(n_950), .Y(n_935) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
AND2x2_ASAP7_75t_L g978 ( .A(n_979), .B(n_984), .Y(n_978) );
INVx1_ASAP7_75t_L g1257 ( .A(n_979), .Y(n_1257) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_982), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g1263 ( .A(n_980), .B(n_983), .Y(n_1263) );
INVx1_ASAP7_75t_L g1265 ( .A(n_980), .Y(n_1265) );
HB1xp67_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_983), .B(n_1265), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_986), .Y(n_984) );
AND2x4_ASAP7_75t_SL g1255 ( .A(n_986), .B(n_1256), .Y(n_1255) );
OAI21xp33_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_994), .B(n_1193), .Y(n_987) );
BUFx2_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_990), .B(n_991), .Y(n_989) );
AND2x6_ASAP7_75t_L g1000 ( .A(n_990), .B(n_1001), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_990), .B(n_1003), .Y(n_1002) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_990), .B(n_991), .Y(n_1005) );
AND2x6_ASAP7_75t_L g1006 ( .A(n_990), .B(n_1007), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_990), .B(n_1003), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_990), .B(n_1003), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g1266 ( .A(n_991), .Y(n_1266) );
AND2x2_ASAP7_75t_L g991 ( .A(n_992), .B(n_993), .Y(n_991) );
NOR2xp67_ASAP7_75t_SL g994 ( .A(n_995), .B(n_1131), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_1092), .Y(n_995) );
A2O1A1Ixp33_ASAP7_75t_SL g996 ( .A1(n_997), .A2(n_1008), .B(n_1041), .C(n_1087), .Y(n_996) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_997), .B(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g1102 ( .A(n_997), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_997), .B(n_1130), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_997), .B(n_1079), .Y(n_1154) );
INVx1_ASAP7_75t_L g1185 ( .A(n_997), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_997), .B(n_1025), .Y(n_1190) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1044 ( .A(n_998), .Y(n_1044) );
INVx1_ASAP7_75t_L g1116 ( .A(n_998), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_998), .B(n_1039), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_998), .B(n_1086), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_998), .B(n_1025), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_999), .B(n_1004), .Y(n_998) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1024), .B1(n_1031), .B2(n_1040), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1021), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1011), .B(n_1028), .Y(n_1141) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_1012), .B(n_1050), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_1012), .B(n_1056), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1018), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1013), .B(n_1050), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1013), .B(n_1073), .Y(n_1072) );
A2O1A1Ixp33_ASAP7_75t_L g1134 ( .A1(n_1013), .A2(n_1116), .B(n_1135), .C(n_1137), .Y(n_1134) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_1014), .B(n_1023), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1014), .B(n_1018), .Y(n_1065) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1014), .B(n_1050), .Y(n_1160) );
NOR2xp33_ASAP7_75t_L g1165 ( .A(n_1014), .B(n_1166), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1018), .Y(n_1023) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1018), .Y(n_1040) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1018), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1018), .B(n_1056), .Y(n_1125) );
NAND2x1_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1020), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1021), .B(n_1056), .Y(n_1157) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_1022), .B(n_1056), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1028), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g1039 ( .A(n_1025), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_1025), .B(n_1036), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_1025), .B(n_1076), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_1025), .A2(n_1119), .B1(n_1138), .B2(n_1156), .Y(n_1155) );
AND2x4_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
INVx3_ASAP7_75t_L g1033 ( .A(n_1028), .Y(n_1033) );
CKINVDCx5p33_ASAP7_75t_R g1048 ( .A(n_1028), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1028), .B(n_1050), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1028), .B(n_1072), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1028), .B(n_1102), .Y(n_1126) );
AND2x4_ASAP7_75t_SL g1028 ( .A(n_1029), .B(n_1030), .Y(n_1028) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
NOR2xp33_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1034), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1033), .B(n_1056), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1033), .B(n_1035), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1144 ( .A(n_1033), .B(n_1145), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1033), .B(n_1065), .Y(n_1152) );
CKINVDCx14_ASAP7_75t_R g1171 ( .A(n_1033), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1033), .B(n_1054), .Y(n_1174) );
AOI211xp5_ASAP7_75t_L g1100 ( .A1(n_1034), .A2(n_1101), .B(n_1103), .C(n_1106), .Y(n_1100) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1039), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1035), .B(n_1096), .Y(n_1095) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1035), .Y(n_1145) );
NOR2xp33_ASAP7_75t_L g1168 ( .A(n_1035), .B(n_1097), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1035), .B(n_1170), .Y(n_1169) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_1036), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1036), .B(n_1039), .Y(n_1069) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1036), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1038), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_1039), .B(n_1044), .Y(n_1043) );
NAND3xp33_ASAP7_75t_L g1143 ( .A(n_1039), .B(n_1065), .C(n_1144), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1040), .B(n_1056), .Y(n_1148) );
NAND4xp25_ASAP7_75t_SL g1041 ( .A(n_1042), .B(n_1060), .C(n_1077), .D(n_1083), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g1042 ( .A1(n_1043), .A2(n_1045), .B1(n_1054), .B2(n_1057), .Y(n_1042) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1044), .Y(n_1099) );
OAI211xp5_ASAP7_75t_L g1163 ( .A1(n_1044), .A2(n_1164), .B(n_1167), .C(n_1169), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1053), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
OAI21xp5_ASAP7_75t_L g1111 ( .A1(n_1047), .A2(n_1058), .B(n_1112), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1049), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1048), .B(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1048), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_1048), .B(n_1118), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1048), .B(n_1075), .Y(n_1136) );
NOR2xp33_ASAP7_75t_L g1137 ( .A(n_1048), .B(n_1138), .Y(n_1137) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1050), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_1050), .B(n_1098), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1050), .B(n_1073), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_1050), .A2(n_1159), .B1(n_1161), .B2(n_1162), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1052), .Y(n_1050) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1053), .Y(n_1061) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_1055), .B(n_1085), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_1056), .B(n_1064), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1056), .B(n_1072), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1056), .B(n_1152), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1058), .B(n_1115), .Y(n_1114) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
O2A1O1Ixp33_ASAP7_75t_L g1060 ( .A1(n_1061), .A2(n_1062), .B(n_1066), .C(n_1070), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g1164 ( .A1(n_1061), .A2(n_1069), .B1(n_1145), .B2(n_1165), .Y(n_1164) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
AOI21xp5_ASAP7_75t_L g1070 ( .A1(n_1063), .A2(n_1071), .B(n_1075), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1081 ( .A(n_1064), .B(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1065), .B(n_1074), .Y(n_1096) );
OAI211xp5_ASAP7_75t_L g1123 ( .A1(n_1065), .A2(n_1068), .B(n_1124), .C(n_1126), .Y(n_1123) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1068), .Y(n_1138) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1069), .B(n_1185), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1074), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1072), .B(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1074), .Y(n_1166) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1075), .Y(n_1110) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1075), .Y(n_1130) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1076), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1080), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1101 ( .A(n_1079), .B(n_1102), .Y(n_1101) );
AOI21xp5_ASAP7_75t_L g1175 ( .A1(n_1079), .A2(n_1176), .B(n_1178), .Y(n_1175) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
A2O1A1Ixp33_ASAP7_75t_L g1107 ( .A1(n_1081), .A2(n_1108), .B(n_1109), .C(n_1111), .Y(n_1107) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1082), .Y(n_1177) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
CKINVDCx14_ASAP7_75t_R g1106 ( .A(n_1087), .Y(n_1106) );
A2O1A1Ixp33_ASAP7_75t_L g1172 ( .A1(n_1087), .A2(n_1173), .B(n_1175), .C(n_1180), .Y(n_1172) );
INVx3_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
OAI221xp5_ASAP7_75t_L g1146 ( .A1(n_1088), .A2(n_1117), .B1(n_1121), .B2(n_1147), .C(n_1149), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1091), .Y(n_1088) );
NOR5xp2_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1100), .C(n_1107), .D(n_1113), .E(n_1127), .Y(n_1092) );
AOI21xp33_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1097), .B(n_1099), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVxp67_ASAP7_75t_L g1108 ( .A(n_1096), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1105), .Y(n_1103) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1105), .Y(n_1112) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
AOI211xp5_ASAP7_75t_L g1139 ( .A1(n_1110), .A2(n_1140), .B(n_1142), .C(n_1146), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1112), .B(n_1171), .Y(n_1179) );
OAI221xp5_ASAP7_75t_SL g1113 ( .A1(n_1114), .A2(n_1117), .B1(n_1119), .B2(n_1121), .C(n_1123), .Y(n_1113) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1114), .Y(n_1162) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1129), .Y(n_1127) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1128), .Y(n_1153) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1129), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1182), .Y(n_1131) );
OAI21xp5_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1163), .B(n_1172), .Y(n_1132) );
NAND4xp25_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1139), .C(n_1150), .D(n_1158), .Y(n_1133) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
OAI21xp5_ASAP7_75t_SL g1183 ( .A1(n_1147), .A2(n_1184), .B(n_1186), .Y(n_1183) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
O2A1O1Ixp33_ASAP7_75t_L g1150 ( .A1(n_1151), .A2(n_1153), .B(n_1154), .C(n_1155), .Y(n_1150) );
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_1151), .A2(n_1171), .B1(n_1183), .B2(n_1191), .Y(n_1182) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1157), .B(n_1171), .Y(n_1170) );
OAI31xp33_ASAP7_75t_L g1186 ( .A1(n_1159), .A2(n_1187), .A3(n_1189), .B(n_1190), .Y(n_1186) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
A2O1A1Ixp33_ASAP7_75t_L g1191 ( .A1(n_1160), .A2(n_1184), .B(n_1188), .C(n_1192), .Y(n_1191) );
INVxp67_ASAP7_75t_SL g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1184), .Y(n_1189) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1190), .Y(n_1192) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g1261 ( .A(n_1196), .Y(n_1261) );
NAND4xp25_ASAP7_75t_SL g1196 ( .A(n_1197), .B(n_1209), .C(n_1229), .D(n_1247), .Y(n_1196) );
AO21x1_ASAP7_75t_L g1197 ( .A1(n_1198), .A2(n_1201), .B(n_1208), .Y(n_1197) );
AOI33xp33_ASAP7_75t_L g1209 ( .A1(n_1210), .A2(n_1211), .A3(n_1217), .B1(n_1222), .B2(n_1225), .B3(n_1228), .Y(n_1209) );
BUFx2_ASAP7_75t_SL g1212 ( .A(n_1213), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx2_ASAP7_75t_SL g1214 ( .A(n_1215), .Y(n_1214) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1221), .Y(n_1227) );
BUFx2_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx2_ASAP7_75t_SL g1244 ( .A(n_1233), .Y(n_1244) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
AO21x1_ASAP7_75t_L g1247 ( .A1(n_1248), .A2(n_1249), .B(n_1253), .Y(n_1247) );
BUFx3_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVxp67_ASAP7_75t_SL g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
HB1xp67_ASAP7_75t_SL g1262 ( .A(n_1263), .Y(n_1262) );
OAI21xp5_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1266), .B(n_1267), .Y(n_1264) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
endmodule