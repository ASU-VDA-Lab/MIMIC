module fake_netlist_1_12362_n_687 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_687);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_687;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_60), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_58), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_68), .Y(n_89) );
BUFx10_ASAP7_75t_L g90 ( .A(n_61), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_78), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_23), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_3), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_76), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_14), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_16), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_27), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_73), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_53), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_40), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_49), .Y(n_103) );
BUFx8_ASAP7_75t_SL g104 ( .A(n_39), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_21), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_32), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_62), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_65), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_81), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_10), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_16), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_4), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_85), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_5), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_63), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_0), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_83), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_84), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_34), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_56), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_30), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_36), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_44), .Y(n_123) );
BUFx6f_ASAP7_75t_SL g124 ( .A(n_80), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_46), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_120), .B(n_1), .Y(n_126) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_91), .A2(n_45), .B(n_79), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_120), .B(n_112), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_115), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_115), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_100), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_100), .B(n_1), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_101), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_92), .B(n_2), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_114), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_119), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_99), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_114), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_104), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_101), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_92), .B(n_5), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_119), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_132), .A2(n_94), .B1(n_95), .B2(n_98), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_133), .B(n_109), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_133), .B(n_109), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_131), .B(n_117), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_130), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_136), .Y(n_154) );
OAI22xp33_ASAP7_75t_L g155 ( .A1(n_141), .A2(n_98), .B1(n_95), .B2(n_93), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_132), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_130), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_127), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_130), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_128), .B(n_96), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_143), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_140), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_130), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_144), .Y(n_173) );
INVxp67_ASAP7_75t_SL g174 ( .A(n_126), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
AND2x6_ASAP7_75t_L g176 ( .A(n_135), .B(n_117), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_132), .B(n_118), .Y(n_177) );
XOR2x2_ASAP7_75t_SL g178 ( .A(n_141), .B(n_93), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_174), .B(n_126), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_177), .A2(n_138), .B(n_134), .C(n_129), .Y(n_181) );
NOR2x1p5_ASAP7_75t_L g182 ( .A(n_164), .B(n_146), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_174), .B(n_145), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_161), .B(n_134), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_156), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_148), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_161), .B(n_134), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_148), .B(n_137), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_176), .A2(n_145), .B1(n_137), .B2(n_138), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_149), .B(n_86), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g197 ( .A(n_158), .B(n_102), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_176), .A2(n_116), .B1(n_94), .B2(n_114), .Y(n_198) );
AOI222xp33_ASAP7_75t_L g199 ( .A1(n_155), .A2(n_97), .B1(n_116), .B2(n_110), .C1(n_105), .C2(n_142), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_149), .B(n_87), .Y(n_200) );
AND2x6_ASAP7_75t_SL g201 ( .A(n_178), .B(n_118), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_150), .B(n_90), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_155), .A2(n_108), .B1(n_129), .B2(n_111), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_176), .A2(n_124), .B1(n_129), .B2(n_130), .Y(n_205) );
BUFx5_ASAP7_75t_L g206 ( .A(n_176), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_158), .B(n_127), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_176), .B(n_89), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_176), .B(n_103), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_147), .B(n_90), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_176), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_176), .B(n_106), .Y(n_212) );
AND2x6_ASAP7_75t_SL g213 ( .A(n_178), .B(n_121), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_147), .B(n_90), .Y(n_214) );
O2A1O1Ixp5_ASAP7_75t_L g215 ( .A1(n_158), .A2(n_123), .B(n_121), .C(n_142), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_166), .B(n_90), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_176), .B(n_107), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_176), .B(n_113), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
NOR3xp33_ASAP7_75t_L g220 ( .A(n_178), .B(n_111), .C(n_123), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_183), .B(n_177), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_220), .A2(n_139), .B(n_173), .C(n_171), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_202), .A2(n_139), .B(n_130), .C(n_175), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_189), .A2(n_158), .B1(n_124), .B2(n_130), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_193), .Y(n_226) );
OR2x6_ASAP7_75t_SL g227 ( .A(n_204), .B(n_180), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_189), .B(n_6), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_191), .A2(n_127), .B(n_160), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_202), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_192), .A2(n_124), .B1(n_122), .B2(n_125), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_185), .A2(n_127), .B(n_163), .Y(n_232) );
INVx6_ASAP7_75t_L g233 ( .A(n_182), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_190), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_179), .A2(n_127), .B(n_163), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
AO32x2_ASAP7_75t_L g237 ( .A1(n_211), .A2(n_151), .A3(n_172), .B1(n_157), .B2(n_159), .Y(n_237) );
OAI22x1_ASAP7_75t_L g238 ( .A1(n_204), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_179), .A2(n_165), .B(n_152), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_186), .A2(n_165), .B(n_152), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_203), .B(n_7), .Y(n_241) );
OAI21xp33_ASAP7_75t_L g242 ( .A1(n_197), .A2(n_175), .B(n_173), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_216), .B(n_124), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_186), .A2(n_167), .B(n_154), .Y(n_244) );
NOR4xp25_ASAP7_75t_L g245 ( .A(n_181), .B(n_169), .C(n_171), .D(n_153), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_206), .B(n_168), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_182), .B(n_168), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_211), .B(n_8), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_199), .A2(n_169), .B(n_153), .C(n_160), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_193), .A2(n_167), .B(n_154), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_206), .B(n_168), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_199), .A2(n_170), .B(n_168), .C(n_172), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_193), .A2(n_172), .B(n_159), .Y(n_253) );
NAND2x1_ASAP7_75t_L g254 ( .A(n_184), .B(n_168), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_195), .B(n_9), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_235), .A2(n_207), .B(n_215), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_223), .A2(n_210), .B(n_214), .C(n_188), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_239), .A2(n_193), .B(n_187), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_225), .Y(n_259) );
AND2x6_ASAP7_75t_L g260 ( .A(n_228), .B(n_193), .Y(n_260) );
O2A1O1Ixp5_ASAP7_75t_SL g261 ( .A1(n_255), .A2(n_170), .B(n_207), .C(n_200), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_230), .A2(n_198), .B1(n_184), .B2(n_217), .Y(n_262) );
AOI221x1_ASAP7_75t_L g263 ( .A1(n_242), .A2(n_208), .B1(n_218), .B2(n_209), .C(n_212), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_228), .B(n_184), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_236), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_234), .A2(n_197), .B1(n_206), .B2(n_194), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_233), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_221), .A2(n_194), .B1(n_205), .B2(n_187), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_252), .A2(n_170), .B(n_201), .C(n_213), .Y(n_269) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_232), .A2(n_157), .A3(n_159), .B(n_196), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_229), .A2(n_207), .B(n_253), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_224), .A2(n_157), .B(n_196), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_224), .A2(n_219), .B(n_170), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_227), .B(n_201), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_240), .A2(n_219), .B(n_170), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_248), .B(n_206), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_222), .A2(n_213), .B(n_206), .C(n_11), .Y(n_278) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_238), .A2(n_206), .A3(n_10), .B(n_12), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_265), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_271), .A2(n_272), .B(n_273), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_265), .B(n_248), .Y(n_282) );
NAND3xp33_ASAP7_75t_L g283 ( .A(n_261), .B(n_245), .C(n_241), .Y(n_283) );
NAND2x1p5_ASAP7_75t_L g284 ( .A(n_277), .B(n_246), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_260), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_275), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_271), .A2(n_250), .B(n_244), .Y(n_287) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_273), .A2(n_251), .B(n_237), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_275), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_257), .A2(n_249), .B(n_254), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_274), .B(n_206), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_269), .B(n_206), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_270), .Y(n_293) );
AOI21xp33_ASAP7_75t_L g294 ( .A1(n_266), .A2(n_243), .B(n_231), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_259), .B(n_247), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_272), .A2(n_237), .B(n_247), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_258), .A2(n_237), .B(n_247), .Y(n_297) );
AOI22x1_ASAP7_75t_L g298 ( .A1(n_264), .A2(n_52), .B1(n_82), .B2(n_77), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_264), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_259), .B(n_233), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_278), .A2(n_9), .B(n_12), .C(n_13), .Y(n_301) );
AOI21x1_ASAP7_75t_L g302 ( .A1(n_263), .A2(n_51), .B(n_74), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_293), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_280), .B(n_260), .Y(n_304) );
INVx5_ASAP7_75t_L g305 ( .A(n_299), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_285), .Y(n_306) );
INVxp33_ASAP7_75t_L g307 ( .A(n_300), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_293), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_281), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_280), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_293), .B(n_264), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_286), .B(n_260), .Y(n_313) );
OR2x6_ASAP7_75t_L g314 ( .A(n_285), .B(n_256), .Y(n_314) );
OA21x2_ASAP7_75t_L g315 ( .A1(n_283), .A2(n_256), .B(n_261), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_295), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_289), .B(n_279), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_289), .B(n_279), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_282), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_295), .B(n_279), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_296), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_299), .B(n_279), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_288), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_282), .B(n_279), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_288), .Y(n_329) );
OAI321xp33_ASAP7_75t_L g330 ( .A1(n_301), .A2(n_262), .A3(n_268), .B1(n_260), .B2(n_276), .C(n_19), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_287), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_292), .B(n_270), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_288), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_288), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_303), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_328), .B(n_297), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_312), .B(n_308), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_328), .B(n_297), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_305), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_308), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_318), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_305), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_318), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_327), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_318), .B(n_292), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_317), .B(n_291), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_319), .B(n_283), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_327), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_310), .Y(n_355) );
NOR2x1_ASAP7_75t_SL g356 ( .A(n_314), .B(n_291), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_312), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_319), .B(n_270), .Y(n_358) );
NAND2x1_ASAP7_75t_L g359 ( .A(n_314), .B(n_260), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_311), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_314), .B(n_270), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_305), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_312), .B(n_270), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_323), .B(n_317), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_328), .B(n_290), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_329), .Y(n_367) );
OR2x6_ASAP7_75t_L g368 ( .A(n_314), .B(n_284), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_314), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_307), .B(n_267), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_316), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_325), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_314), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_314), .B(n_287), .Y(n_376) );
INVx4_ASAP7_75t_L g377 ( .A(n_305), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_325), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_323), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_323), .B(n_284), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_333), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_333), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_333), .B(n_260), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_304), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_335), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_321), .B(n_13), .Y(n_387) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_304), .B(n_298), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_316), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_381), .B(n_334), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_381), .B(n_334), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_382), .B(n_334), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_346), .B(n_332), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_346), .B(n_335), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_341), .B(n_322), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_348), .B(n_320), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_360), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_377), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_348), .B(n_320), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_376), .B(n_332), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_383), .A2(n_326), .B1(n_322), .B2(n_331), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_364), .B(n_320), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_355), .B(n_326), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_363), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_354), .B(n_320), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_354), .B(n_324), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_349), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_364), .B(n_324), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_358), .B(n_324), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_347), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_363), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_372), .B(n_331), .C(n_332), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_342), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_336), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_336), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_342), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_379), .B(n_332), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_352), .B(n_305), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_337), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_358), .B(n_316), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_349), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_350), .B(n_315), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_350), .B(n_315), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_357), .B(n_305), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_387), .B(n_15), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_347), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_387), .B(n_305), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_365), .B(n_315), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_337), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_370), .B(n_305), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_377), .A2(n_313), .B1(n_306), .B2(n_298), .Y(n_432) );
NAND2x1_ASAP7_75t_L g433 ( .A(n_377), .B(n_306), .Y(n_433) );
NOR2xp33_ASAP7_75t_SL g434 ( .A(n_344), .B(n_362), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_383), .A2(n_306), .B1(n_313), .B2(n_294), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_365), .B(n_315), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_347), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_370), .B(n_15), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_338), .B(n_343), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_374), .B(n_378), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_340), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_344), .B(n_17), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_353), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_374), .B(n_17), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_378), .B(n_309), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_338), .B(n_309), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_380), .B(n_309), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_338), .B(n_309), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_361), .B(n_309), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_362), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_380), .B(n_309), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_345), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_351), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_385), .B(n_309), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_345), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_343), .B(n_309), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_361), .B(n_302), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_343), .B(n_302), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_366), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_339), .B(n_18), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_366), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_384), .B(n_18), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_339), .B(n_19), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_385), .B(n_20), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_430), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_405), .B(n_386), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_394), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_412), .B(n_386), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_398), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_414), .B(n_369), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_417), .B(n_367), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_399), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_453), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_423), .B(n_361), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_408), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_421), .B(n_367), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_408), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_423), .B(n_361), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_424), .B(n_369), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_424), .B(n_371), .Y(n_480) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_433), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_390), .B(n_356), .Y(n_482) );
NAND2x1_ASAP7_75t_L g483 ( .A(n_399), .B(n_375), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_429), .B(n_375), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_429), .B(n_376), .Y(n_485) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_462), .B(n_330), .C(n_388), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_422), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_421), .B(n_368), .Y(n_488) );
AND2x4_ASAP7_75t_SL g489 ( .A(n_460), .B(n_368), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_439), .B(n_356), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_390), .B(n_389), .Y(n_492) );
INVx3_ASAP7_75t_SL g493 ( .A(n_450), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_440), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_415), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_415), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_416), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_391), .B(n_389), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_433), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_443), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_426), .A2(n_368), .B1(n_376), .B2(n_359), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_420), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_420), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_436), .B(n_368), .Y(n_505) );
INVxp67_ASAP7_75t_L g506 ( .A(n_413), .Y(n_506) );
AND2x4_ASAP7_75t_SL g507 ( .A(n_460), .B(n_373), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_391), .B(n_373), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_392), .B(n_359), .Y(n_509) );
NAND4xp25_ASAP7_75t_L g510 ( .A(n_402), .B(n_294), .C(n_21), .D(n_22), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_427), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_411), .B(n_330), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_441), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_436), .B(n_20), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_410), .B(n_22), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_410), .B(n_23), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_411), .B(n_24), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_439), .B(n_24), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_419), .B(n_25), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_392), .B(n_25), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_452), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_395), .B(n_26), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_395), .B(n_26), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_446), .B(n_27), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_446), .B(n_284), .Y(n_525) );
NOR2x1p5_ASAP7_75t_L g526 ( .A(n_425), .B(n_28), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_448), .B(n_29), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_448), .B(n_31), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_452), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_409), .B(n_33), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_455), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_455), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_456), .B(n_35), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_396), .Y(n_534) );
OR2x6_ASAP7_75t_L g535 ( .A(n_431), .B(n_37), .Y(n_535) );
BUFx2_ASAP7_75t_L g536 ( .A(n_437), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_404), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_434), .B(n_38), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_409), .B(n_41), .Y(n_539) );
NOR2xp33_ASAP7_75t_SL g540 ( .A(n_493), .B(n_432), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_465), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_465), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_474), .B(n_401), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_491), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_493), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_494), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_467), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_534), .B(n_407), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_472), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_510), .A2(n_442), .B(n_464), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_537), .B(n_407), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_473), .B(n_438), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_476), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_500), .B(n_401), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_495), .B(n_406), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_474), .B(n_401), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_469), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_475), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_478), .B(n_401), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_511), .B(n_444), .Y(n_560) );
XNOR2xp5_ASAP7_75t_L g561 ( .A(n_518), .B(n_464), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_502), .A2(n_428), .B1(n_435), .B2(n_463), .Y(n_562) );
AOI21xp5_ASAP7_75t_SL g563 ( .A1(n_526), .A2(n_463), .B(n_457), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_536), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_496), .B(n_397), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_515), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_497), .B(n_400), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_478), .B(n_393), .Y(n_568) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_477), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_514), .B(n_406), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_475), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_503), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_504), .B(n_461), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_507), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_480), .B(n_418), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_485), .B(n_393), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_471), .B(n_418), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_485), .B(n_449), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_468), .B(n_403), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_489), .A2(n_449), .B1(n_458), .B2(n_457), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_479), .B(n_403), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_519), .B(n_518), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_486), .A2(n_449), .B1(n_447), .B2(n_451), .Y(n_583) );
NOR3x1_ASAP7_75t_L g584 ( .A(n_483), .B(n_451), .C(n_447), .Y(n_584) );
OR2x6_ASAP7_75t_L g585 ( .A(n_500), .B(n_445), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_513), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_521), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_505), .B(n_458), .Y(n_588) );
OAI21xp33_ASAP7_75t_SL g589 ( .A1(n_490), .A2(n_461), .B(n_454), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_529), .B(n_459), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_505), .B(n_454), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_492), .B(n_457), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_531), .B(n_42), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_484), .B(n_43), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_532), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_484), .B(n_47), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_506), .B(n_48), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_481), .B(n_50), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_470), .B(n_54), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_541), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_542), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_548), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_545), .B(n_522), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_561), .A2(n_516), .B1(n_517), .B2(n_535), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_581), .B(n_508), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_589), .A2(n_564), .B(n_517), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_548), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_579), .B(n_499), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_550), .A2(n_486), .B1(n_523), .B2(n_525), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_551), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_564), .B(n_520), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_574), .A2(n_535), .B1(n_482), .B2(n_515), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_566), .B(n_466), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_578), .B(n_525), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_585), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_543), .B(n_524), .Y(n_617) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_585), .A2(n_538), .B(n_512), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_563), .A2(n_538), .B(n_540), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_577), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_556), .B(n_524), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_555), .Y(n_622) );
NAND4xp25_ASAP7_75t_SL g623 ( .A(n_574), .B(n_523), .C(n_509), .D(n_488), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_540), .A2(n_481), .B(n_535), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_569), .B(n_481), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_549), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_565), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_558), .Y(n_628) );
OAI22xp33_ASAP7_75t_SL g629 ( .A1(n_584), .A2(n_512), .B1(n_539), .B2(n_530), .Y(n_629) );
INVxp33_ASAP7_75t_L g630 ( .A(n_582), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_565), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_598), .A2(n_481), .B(n_477), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_562), .A2(n_533), .B1(n_527), .B2(n_528), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_567), .Y(n_634) );
INVxp67_ASAP7_75t_L g635 ( .A(n_560), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_567), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_580), .A2(n_501), .B1(n_498), .B2(n_487), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_552), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_609), .A2(n_583), .B1(n_554), .B2(n_570), .Y(n_639) );
NAND4xp25_ASAP7_75t_L g640 ( .A(n_609), .B(n_597), .C(n_596), .D(n_594), .Y(n_640) );
AOI32xp33_ASAP7_75t_L g641 ( .A1(n_604), .A2(n_554), .A3(n_559), .B1(n_568), .B2(n_576), .Y(n_641) );
AOI32xp33_ASAP7_75t_L g642 ( .A1(n_637), .A2(n_599), .A3(n_588), .B1(n_591), .B2(n_553), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_623), .A2(n_612), .B1(n_635), .B2(n_638), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_606), .A2(n_544), .B1(n_546), .B2(n_597), .C(n_592), .Y(n_644) );
INVxp67_ASAP7_75t_SL g645 ( .A(n_625), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g646 ( .A1(n_638), .A2(n_595), .B1(n_547), .B2(n_557), .C1(n_587), .C2(n_586), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_619), .A2(n_572), .B(n_593), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g648 ( .A1(n_611), .A2(n_575), .A3(n_571), .B1(n_573), .B2(n_590), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_616), .B(n_590), .Y(n_649) );
NOR3xp33_ASAP7_75t_L g650 ( .A(n_618), .B(n_593), .C(n_573), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_633), .A2(n_55), .B1(n_57), .B2(n_59), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_622), .Y(n_652) );
AOI211xp5_ASAP7_75t_SL g653 ( .A1(n_624), .A2(n_64), .B(n_66), .C(n_67), .Y(n_653) );
AO21x1_ASAP7_75t_L g654 ( .A1(n_625), .A2(n_69), .B(n_70), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_632), .A2(n_71), .B(n_72), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g656 ( .A1(n_630), .A2(n_75), .B(n_603), .C(n_626), .Y(n_656) );
OAI31xp33_ASAP7_75t_L g657 ( .A1(n_633), .A2(n_614), .A3(n_610), .B(n_602), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_628), .B(n_613), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_627), .A2(n_636), .B(n_634), .Y(n_659) );
AOI21xp33_ASAP7_75t_SL g660 ( .A1(n_614), .A2(n_600), .B(n_601), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_631), .A2(n_607), .B1(n_620), .B2(n_608), .C(n_605), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_617), .A2(n_621), .B(n_615), .Y(n_662) );
NAND5xp2_ASAP7_75t_L g663 ( .A(n_619), .B(n_609), .C(n_624), .D(n_606), .E(n_540), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_638), .B(n_635), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_618), .A2(n_606), .B(n_619), .C(n_629), .Y(n_665) );
NAND3xp33_ASAP7_75t_SL g666 ( .A(n_665), .B(n_656), .C(n_654), .Y(n_666) );
NOR2x1_ASAP7_75t_L g667 ( .A(n_663), .B(n_647), .Y(n_667) );
AOI221x1_ASAP7_75t_L g668 ( .A1(n_664), .A2(n_650), .B1(n_651), .B2(n_660), .C(n_639), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_664), .B(n_643), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_646), .B(n_657), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_649), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_667), .A2(n_641), .B1(n_642), .B2(n_661), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_669), .B(n_648), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_671), .B(n_662), .Y(n_674) );
AOI211x1_ASAP7_75t_SL g675 ( .A1(n_670), .A2(n_640), .B(n_658), .C(n_655), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_674), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_675), .B(n_668), .Y(n_677) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_672), .B(n_666), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_676), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_678), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_679), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g682 ( .A(n_680), .B(n_677), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_681), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_682), .B(n_673), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_684), .A2(n_645), .B(n_653), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_685), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_644), .B1(n_659), .B2(n_652), .Y(n_687) );
endmodule