module fake_jpeg_9737_n_224 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_23),
.Y(n_46)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_21),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

OR2x4_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_1),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_37),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_19),
.B1(n_34),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_56),
.B1(n_25),
.B2(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_60),
.Y(n_79)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_17),
.B1(n_24),
.B2(n_30),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_31),
.A3(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_27),
.B(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_33),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_30),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_67),
.B(n_88),
.Y(n_109)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_70),
.Y(n_111)
);

XNOR2x1_ASAP7_75t_SL g110 ( 
.A(n_69),
.B(n_92),
.Y(n_110)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_36),
.B1(n_41),
.B2(n_38),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_78),
.B1(n_54),
.B2(n_59),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_41),
.B1(n_36),
.B2(n_45),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_75),
.B1(n_94),
.B2(n_4),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_45),
.B1(n_37),
.B2(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_22),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_31),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_25),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_86),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_28),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_57),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_5),
.Y(n_114)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_2),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_37),
.C(n_33),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_59),
.C(n_54),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_37),
.B1(n_33),
.B2(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_5),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_93),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_114),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_120),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_95),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_67),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_R g121 ( 
.A(n_110),
.B(n_69),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_130),
.B(n_135),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_105),
.C(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_129),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_109),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_136),
.C(n_114),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_71),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_106),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_142),
.Y(n_162)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_134),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_71),
.B(n_69),
.Y(n_135)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_96),
.A3(n_92),
.B1(n_73),
.B2(n_77),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_94),
.B1(n_91),
.B2(n_88),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_140),
.B1(n_108),
.B2(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_76),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_115),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_92),
.B1(n_89),
.B2(n_76),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_89),
.B1(n_14),
.B2(n_11),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_108),
.B1(n_114),
.B2(n_11),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_102),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_127),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_152),
.B1(n_158),
.B2(n_161),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_97),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_130),
.C(n_121),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_156),
.B(n_122),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_116),
.B(n_99),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_163),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_99),
.B1(n_101),
.B2(n_12),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_169),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_176),
.C(n_145),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_177),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_128),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_178),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_125),
.C(n_133),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_142),
.C(n_134),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g178 ( 
.A(n_161),
.B(n_132),
.C(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_171),
.C(n_167),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_165),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_190),
.B(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_152),
.B1(n_151),
.B2(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_154),
.B(n_163),
.C(n_160),
.D(n_150),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_144),
.B(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_193),
.C(n_194),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_176),
.C(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_144),
.C(n_164),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_166),
.C(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_199),
.C(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_147),
.C(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_147),
.C(n_124),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_208),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

AOI321xp33_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_190),
.A3(n_191),
.B1(n_183),
.B2(n_184),
.C(n_187),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_184),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_187),
.C(n_183),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_212),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_180),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_207),
.Y(n_216)
);

OA21x2_ASAP7_75t_SL g215 ( 
.A1(n_213),
.A2(n_202),
.B(n_211),
.Y(n_215)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_16),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_217),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_124),
.B(n_12),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_14),
.B(n_15),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_9),
.B(n_10),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_218),
.B(n_10),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_222),
.Y(n_224)
);


endmodule