module fake_jpeg_23355_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_20),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_38),
.B(n_0),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_7),
.B(n_14),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_49),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_18),
.B1(n_31),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_35),
.B1(n_18),
.B2(n_23),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_53),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_30),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_34),
.C(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_17),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_17),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_73),
.B(n_37),
.Y(n_103)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NAND2x1_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_29),
.Y(n_73)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_82),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_35),
.B1(n_42),
.B2(n_20),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_19),
.B1(n_24),
.B2(n_51),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_78),
.B1(n_54),
.B2(n_69),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_65),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_90),
.B(n_22),
.Y(n_130)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_94),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_49),
.B1(n_50),
.B2(n_42),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_54),
.B1(n_51),
.B2(n_42),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_37),
.A3(n_27),
.B1(n_32),
.B2(n_41),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_79),
.A3(n_73),
.B1(n_32),
.B2(n_40),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_62),
.B(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_37),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_56),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_110),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_41),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_48),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_69),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_31),
.B1(n_45),
.B2(n_32),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_34),
.B1(n_19),
.B2(n_24),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_34),
.B1(n_48),
.B2(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_30),
.Y(n_116)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_123),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_127),
.B(n_110),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g124 ( 
.A(n_99),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_60),
.B1(n_75),
.B2(n_67),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_100),
.B1(n_112),
.B2(n_91),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_102),
.B(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_40),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_130),
.Y(n_154)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_131),
.Y(n_159)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_80),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_40),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_97),
.B1(n_101),
.B2(n_98),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_137),
.A2(n_142),
.B1(n_148),
.B2(n_151),
.Y(n_178)
);

OAI22x1_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_126),
.B1(n_117),
.B2(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_149),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_141),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_127),
.B(n_95),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_107),
.B1(n_93),
.B2(n_108),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_135),
.A2(n_21),
.B1(n_22),
.B2(n_75),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_41),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_145),
.C(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_29),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_158),
.B(n_125),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_77),
.B1(n_43),
.B2(n_40),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_41),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_132),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_121),
.B(n_29),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_141),
.C(n_145),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_21),
.B(n_29),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_10),
.Y(n_160)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_117),
.B(n_118),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_172),
.B(n_176),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_173),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_183),
.B1(n_158),
.B2(n_143),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_177),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_156),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_128),
.A3(n_136),
.B1(n_130),
.B2(n_115),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_155),
.Y(n_197)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_124),
.B1(n_129),
.B2(n_131),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_131),
.B1(n_129),
.B2(n_119),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_151),
.B1(n_124),
.B2(n_119),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_193),
.B1(n_199),
.B2(n_200),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_157),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_192),
.C(n_194),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_176),
.B1(n_163),
.B2(n_169),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_201),
.B1(n_26),
.B2(n_1),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_152),
.C(n_140),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_142),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_148),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_197),
.C(n_8),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_124),
.B1(n_89),
.B2(n_72),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_89),
.B1(n_72),
.B2(n_26),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_169),
.A2(n_26),
.B1(n_29),
.B2(n_2),
.Y(n_201)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_165),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_212),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_167),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_216),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_177),
.B1(n_172),
.B2(n_168),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_190),
.B(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_172),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_184),
.B1(n_182),
.B2(n_181),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_188),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_187),
.Y(n_219)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_195),
.C(n_194),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_230),
.C(n_232),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_197),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_208),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_220),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_202),
.C(n_200),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_196),
.C(n_6),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_206),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_221),
.B1(n_215),
.B2(n_214),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_211),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_223),
.C(n_232),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_242),
.A2(n_226),
.B(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_208),
.B(n_205),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_8),
.B(n_10),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_253),
.C(n_239),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_222),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_236),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_256),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_253),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_242),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_259),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_239),
.C(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_250),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_11),
.B(n_12),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_238),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_11),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_10),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_266),
.B(n_267),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_262),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_264),
.B(n_12),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_270),
.A2(n_11),
.B(n_14),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_14),
.Y(n_272)
);


endmodule