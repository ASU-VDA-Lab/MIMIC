module fake_jpeg_8220_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_1),
.C(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx2_ASAP7_75t_SL g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_19),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_36),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_20),
.B1(n_22),
.B2(n_26),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_54),
.B1(n_59),
.B2(n_63),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_20),
.B1(n_22),
.B2(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_33),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_18),
.B1(n_26),
.B2(n_42),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_27),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_63)
);

NAND2x1_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_43),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_43),
.Y(n_98)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_69),
.Y(n_90)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_75),
.Y(n_99)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_80),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_35),
.B1(n_37),
.B2(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_34),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_83),
.B1(n_61),
.B2(n_47),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_39),
.B1(n_17),
.B2(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_105),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_106),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_64),
.C(n_65),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_100),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_30),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_68),
.C(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_32),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_39),
.B1(n_57),
.B2(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_3),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_84),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_4),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_81),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_47),
.B1(n_57),
.B2(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_126),
.B1(n_96),
.B2(n_94),
.Y(n_144)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_129),
.B(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_43),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_127),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_25),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_28),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_28),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_106),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_85),
.B1(n_69),
.B2(n_31),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_79),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_93),
.B1(n_115),
.B2(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_95),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_131),
.B(n_136),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_109),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_100),
.B(n_95),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_120),
.B1(n_88),
.B2(n_31),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_140),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_107),
.C(n_105),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_109),
.B1(n_113),
.B2(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_145),
.B(n_147),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_159),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_125),
.C(n_118),
.Y(n_150)
);

AOI321xp33_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_140),
.A3(n_145),
.B1(n_134),
.B2(n_144),
.C(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_88),
.B(n_29),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_160),
.B(n_161),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_158),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_13),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_5),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_28),
.B(n_79),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_29),
.B(n_28),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_143),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_142),
.C(n_136),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_163),
.A2(n_171),
.B(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_141),
.C(n_132),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_169),
.C(n_173),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_172),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_154),
.C(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_133),
.C(n_30),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_153),
.B(n_162),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_177),
.B(n_179),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_154),
.B1(n_148),
.B2(n_160),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_181),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_160),
.C(n_30),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_6),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_167),
.B(n_172),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_184),
.A2(n_187),
.B(n_8),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_186),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_6),
.B(n_7),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_190),
.B(n_176),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_175),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_176),
.B(n_11),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_194),
.B(n_10),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_196),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_12),
.C(n_13),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_198),
.C(n_200),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_201),
.Y(n_202)
);


endmodule