module fake_jpeg_21514_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_48),
.B1(n_15),
.B2(n_17),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_25),
.B1(n_22),
.B2(n_18),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_21),
.B1(n_17),
.B2(n_31),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_30),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_49),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_34),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_28),
.B1(n_15),
.B2(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_76),
.B(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_42),
.Y(n_70)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_39),
.CI(n_30),
.CON(n_93),
.SN(n_93)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_27),
.B1(n_31),
.B2(n_17),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_53),
.B1(n_54),
.B2(n_44),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_23),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_84),
.Y(n_103)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_30),
.B(n_19),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_80),
.B1(n_82),
.B2(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_55),
.Y(n_79)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_81),
.Y(n_110)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_32),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_55),
.B(n_35),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_55),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_54),
.B1(n_53),
.B2(n_44),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_101),
.B1(n_106),
.B2(n_107),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_64),
.B(n_59),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_105),
.B1(n_112),
.B2(n_79),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_109),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_54),
.B1(n_53),
.B2(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_62),
.A2(n_53),
.B1(n_44),
.B2(n_20),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_55),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_30),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_49),
.B(n_15),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_118),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_126),
.B(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_65),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_128),
.B1(n_129),
.B2(n_132),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_56),
.C(n_57),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_131),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_135),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_95),
.B1(n_86),
.B2(n_102),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_56),
.B1(n_78),
.B2(n_79),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_134),
.B1(n_95),
.B2(n_108),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_63),
.B1(n_75),
.B2(n_81),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_96),
.A2(n_75),
.B1(n_58),
.B2(n_61),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_90),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_61),
.B1(n_58),
.B2(n_68),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_82),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_49),
.B(n_21),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_113),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_101),
.A2(n_80),
.B1(n_29),
.B2(n_72),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_110),
.B1(n_90),
.B2(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_145),
.B1(n_167),
.B2(n_119),
.Y(n_173)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_94),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_166),
.C(n_169),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_113),
.A3(n_108),
.B1(n_112),
.B2(n_97),
.C1(n_29),
.C2(n_27),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_149),
.C(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_158),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_172),
.B1(n_126),
.B2(n_114),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_23),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_164),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_111),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_97),
.B1(n_99),
.B2(n_21),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_97),
.B(n_27),
.Y(n_168)
);

AOI22x1_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_10),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_170),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_29),
.B1(n_26),
.B2(n_28),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_124),
.B1(n_149),
.B2(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_92),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_190),
.B1(n_195),
.B2(n_196),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_178),
.B1(n_193),
.B2(n_147),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_176),
.B(n_159),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_130),
.B(n_131),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_179),
.A2(n_182),
.B(n_189),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_117),
.C(n_115),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_188),
.C(n_169),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_127),
.B(n_122),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_127),
.C(n_122),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_136),
.B(n_129),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_138),
.B1(n_92),
.B2(n_26),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_197),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_142),
.B(n_158),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_0),
.B(n_1),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_0),
.B(n_2),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_0),
.B(n_3),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_168),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_215),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_205),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_143),
.C(n_152),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_168),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_147),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_209),
.B(n_216),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_192),
.B1(n_200),
.B2(n_195),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_162),
.B1(n_160),
.B2(n_159),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_211),
.A2(n_200),
.B1(n_182),
.B2(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_148),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_193),
.Y(n_235)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_230),
.B1(n_239),
.B2(n_216),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_214),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_238),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_175),
.B1(n_201),
.B2(n_179),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_203),
.B1(n_212),
.B2(n_175),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_188),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_221),
.B(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_236),
.A2(n_208),
.B1(n_217),
.B2(n_205),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_241),
.A2(n_235),
.B1(n_228),
.B2(n_226),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_252),
.B(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_210),
.B1(n_212),
.B2(n_225),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_246),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_204),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_191),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_206),
.C(n_177),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_250),
.C(n_251),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_216),
.C(n_183),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_203),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_222),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_198),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_237),
.C(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_263),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_232),
.B(n_229),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_267),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_185),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_197),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_266),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_213),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_241),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_207),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_261),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_276),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_256),
.A2(n_252),
.B(n_242),
.Y(n_273)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_273),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_251),
.B1(n_207),
.B2(n_255),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_269),
.B1(n_268),
.B2(n_275),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_246),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_191),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_257),
.B(n_263),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_8),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_257),
.B(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_283),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_14),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_10),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_289),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_290),
.A2(n_8),
.B(n_12),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_286),
.A2(n_282),
.B(n_281),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_293),
.C(n_292),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.C(n_11),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_291),
.A2(n_288),
.B(n_11),
.C(n_13),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_13),
.B(n_5),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_4),
.B(n_5),
.Y(n_298)
);

O2A1O1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_298),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_300)
);


endmodule