module fake_netlist_6_4703_n_739 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_739);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_739;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_671;
wire n_726;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_594;
wire n_719;
wire n_565;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g151 ( 
.A(n_52),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_36),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_28),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_1),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_23),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_22),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_15),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_14),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_43),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_61),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_65),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_26),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

CKINVDCx11_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_141),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_64),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_119),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_113),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_29),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_76),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_48),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_95),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_39),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_51),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_10),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_68),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_79),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_19),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_73),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_27),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_30),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_144),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_47),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_40),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_53),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_12),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_101),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_122),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_126),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_83),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_173),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_0),
.B(n_2),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_152),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_173),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_158),
.B(n_3),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_4),
.B(n_5),
.Y(n_225)
);

BUFx8_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_165),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_6),
.Y(n_233)
);

BUFx8_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_151),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_160),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_162),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_200),
.B(n_8),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_207),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_165),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_207),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_229),
.B1(n_233),
.B2(n_217),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_161),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_182),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_219),
.B(n_182),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_250),
.B1(n_219),
.B2(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_248),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_169),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_220),
.B(n_201),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_171),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_220),
.B(n_201),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_172),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_246),
.B(n_155),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_212),
.B(n_230),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_212),
.B(n_157),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_212),
.B(n_178),
.Y(n_282)
);

BUFx6f_ASAP7_75t_SL g283 ( 
.A(n_237),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_208),
.B(n_174),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_243),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_L g289 ( 
.A(n_228),
.B(n_175),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_226),
.B(n_183),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_228),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_214),
.A2(n_206),
.B1(n_179),
.B2(n_199),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_226),
.B(n_185),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_221),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_237),
.A2(n_177),
.B1(n_180),
.B2(n_196),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_215),
.B1(n_225),
.B2(n_210),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_226),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_266),
.B(n_187),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_256),
.Y(n_304)
);

NAND2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_184),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_234),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_294),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_242),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_256),
.A2(n_186),
.B1(n_194),
.B2(n_227),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_251),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_269),
.A2(n_215),
.B1(n_225),
.B2(n_210),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_221),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_253),
.B(n_189),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_296),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_287),
.Y(n_318)
);

INVx8_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_231),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_209),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_231),
.Y(n_322)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_251),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_231),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_252),
.Y(n_328)
);

OR2x6_ASAP7_75t_L g329 ( 
.A(n_258),
.B(n_211),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_211),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_271),
.B(n_231),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_272),
.B(n_213),
.C(n_216),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_254),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_231),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_270),
.B(n_241),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_270),
.B(n_241),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_293),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_241),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_295),
.B(n_190),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_292),
.B(n_241),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_284),
.A2(n_191),
.B1(n_193),
.B2(n_197),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_209),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_274),
.B(n_241),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_289),
.A2(n_235),
.B(n_228),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_252),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_257),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_276),
.B(n_235),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_276),
.B(n_204),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_277),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_277),
.B(n_279),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_279),
.B(n_288),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_257),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_288),
.B(n_216),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_284),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_298),
.B(n_213),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_282),
.B(n_210),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_261),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_260),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_261),
.B(n_18),
.Y(n_359)
);

NOR2x1p5_ASAP7_75t_L g360 ( 
.A(n_262),
.B(n_8),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_321),
.B(n_259),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_262),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_314),
.A2(n_264),
.B(n_268),
.C(n_254),
.Y(n_363)
);

CKINVDCx6p67_ASAP7_75t_R g364 ( 
.A(n_319),
.Y(n_364)
);

A2O1A1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_314),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_356),
.A2(n_84),
.B(n_148),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_356),
.A2(n_81),
.B(n_147),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_312),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_20),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_21),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_9),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_304),
.A2(n_80),
.B1(n_143),
.B2(n_142),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_303),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_350),
.A2(n_78),
.B(n_140),
.Y(n_375)
);

O2A1O1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_315),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_304),
.A2(n_85),
.B1(n_138),
.B2(n_137),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_301),
.B(n_13),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_24),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_351),
.A2(n_75),
.B(n_133),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_334),
.A2(n_74),
.B(n_131),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_72),
.B(n_130),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_309),
.Y(n_384)
);

O2A1O1Ixp33_ASAP7_75t_SL g385 ( 
.A1(n_302),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_385)
);

O2A1O1Ixp33_ASAP7_75t_L g386 ( 
.A1(n_315),
.A2(n_16),
.B(n_17),
.C(n_25),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_313),
.B(n_31),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_306),
.B(n_32),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_310),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_299),
.B(n_37),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_317),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_299),
.B(n_44),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_307),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_302),
.B(n_45),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_307),
.B(n_46),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_339),
.B(n_326),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_353),
.A2(n_49),
.B(n_50),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_54),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_308),
.B(n_56),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_327),
.B(n_57),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_329),
.B(n_58),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_333),
.B(n_59),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_333),
.B(n_60),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_348),
.A2(n_341),
.B(n_359),
.Y(n_407)
);

OAI21xp33_ASAP7_75t_L g408 ( 
.A1(n_311),
.A2(n_62),
.B(n_63),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_325),
.A2(n_331),
.B(n_336),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_335),
.A2(n_66),
.B(n_67),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_358),
.B(n_69),
.Y(n_411)
);

A2O1A1Ixp33_ASAP7_75t_L g412 ( 
.A1(n_332),
.A2(n_70),
.B(n_71),
.C(n_86),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_305),
.A2(n_87),
.B(n_88),
.Y(n_413)
);

NOR3xp33_ASAP7_75t_L g414 ( 
.A(n_316),
.B(n_90),
.C(n_91),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_338),
.A2(n_340),
.B(n_322),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_320),
.A2(n_92),
.B(n_93),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_347),
.A2(n_94),
.B(n_96),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_349),
.B(n_97),
.Y(n_419)
);

O2A1O1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_329),
.A2(n_98),
.B(n_99),
.C(n_100),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_329),
.B(n_102),
.Y(n_421)
);

O2A1O1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_324),
.A2(n_346),
.B(n_345),
.C(n_328),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_360),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_357),
.B(n_107),
.Y(n_424)
);

AOI21x1_ASAP7_75t_L g425 ( 
.A1(n_324),
.A2(n_108),
.B(n_109),
.Y(n_425)
);

NOR2x1_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_346),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_372),
.B(n_323),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_384),
.A2(n_344),
.B(n_111),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_383),
.Y(n_430)
);

BUFx2_ASAP7_75t_SL g431 ( 
.A(n_396),
.Y(n_431)
);

CKINVDCx11_ASAP7_75t_R g432 ( 
.A(n_364),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_361),
.B(n_323),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_110),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_323),
.B(n_319),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_392),
.A2(n_319),
.B(n_115),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_409),
.A2(n_149),
.B(n_117),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_415),
.A2(n_128),
.B(n_120),
.Y(n_439)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_127),
.B(n_121),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_394),
.A2(n_112),
.B(n_123),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_418),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_362),
.B(n_124),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_374),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_404),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_379),
.A2(n_371),
.B1(n_378),
.B2(n_365),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_369),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_407),
.A2(n_399),
.B(n_397),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_421),
.B(n_411),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_423),
.B(n_398),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_422),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_390),
.A2(n_370),
.B(n_401),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_366),
.A2(n_367),
.B(n_413),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_408),
.B(n_424),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_376),
.A2(n_393),
.B1(n_373),
.B2(n_377),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_376),
.B(n_405),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_406),
.A2(n_425),
.B(n_419),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_403),
.Y(n_460)
);

OAI21xp33_ASAP7_75t_SL g461 ( 
.A1(n_391),
.A2(n_382),
.B(n_380),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_386),
.B(n_385),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_375),
.A2(n_400),
.B(n_417),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_386),
.B(n_414),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_412),
.A2(n_420),
.B(n_381),
.Y(n_465)
);

AND3x4_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_410),
.C(n_416),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_362),
.B(n_300),
.Y(n_467)
);

OA22x2_ASAP7_75t_L g468 ( 
.A1(n_361),
.A2(n_311),
.B1(n_304),
.B2(n_315),
.Y(n_468)
);

CKINVDCx9p33_ASAP7_75t_R g469 ( 
.A(n_402),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_372),
.B(n_354),
.Y(n_470)
);

O2A1O1Ixp5_ASAP7_75t_L g471 ( 
.A1(n_379),
.A2(n_302),
.B(n_407),
.C(n_369),
.Y(n_471)
);

OA21x2_ASAP7_75t_L g472 ( 
.A1(n_392),
.A2(n_394),
.B(n_299),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_384),
.B(n_362),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_372),
.B(n_304),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_372),
.B(n_304),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_372),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_432),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_475),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_433),
.Y(n_479)
);

NAND2x1p5_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_428),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_458),
.A2(n_471),
.B(n_450),
.Y(n_481)
);

AO21x1_ASAP7_75t_L g482 ( 
.A1(n_447),
.A2(n_452),
.B(n_457),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_468),
.A2(n_447),
.B1(n_457),
.B2(n_464),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_448),
.A2(n_455),
.B1(n_449),
.B2(n_446),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_440),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_445),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_456),
.A2(n_473),
.B(n_444),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_476),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_468),
.A2(n_473),
.B1(n_451),
.B2(n_462),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_429),
.A2(n_455),
.B(n_465),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_451),
.A2(n_470),
.B1(n_434),
.B2(n_435),
.Y(n_491)
);

OAI21xp33_ASAP7_75t_L g492 ( 
.A1(n_427),
.A2(n_435),
.B(n_430),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_453),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_456),
.A2(n_429),
.B(n_465),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_466),
.A2(n_443),
.B1(n_428),
.B2(n_472),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_461),
.A2(n_472),
.B(n_437),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_443),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_440),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_431),
.B(n_426),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_440),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_469),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_442),
.A2(n_460),
.B1(n_439),
.B2(n_441),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_436),
.A2(n_468),
.B1(n_408),
.B2(n_452),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_463),
.A2(n_458),
.B(n_394),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_474),
.B(n_361),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_476),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_458),
.A2(n_394),
.B(n_392),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_455),
.B(n_452),
.Y(n_510)
);

AOI221xp5_ASAP7_75t_L g511 ( 
.A1(n_457),
.A2(n_253),
.B1(n_256),
.B2(n_315),
.C(n_304),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_361),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g514 ( 
.A(n_474),
.B(n_256),
.C(n_378),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_467),
.B(n_474),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_440),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_361),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_455),
.A2(n_450),
.B(n_454),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_508),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_493),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_493),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_497),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_483),
.A2(n_478),
.B1(n_515),
.B2(n_511),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_497),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_500),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_490),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_490),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_485),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_507),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_496),
.A2(n_518),
.B(n_505),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_502),
.A2(n_481),
.B(n_503),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_485),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_482),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_483),
.B(n_489),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_486),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_490),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_487),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_485),
.Y(n_539)
);

AO21x2_ASAP7_75t_L g540 ( 
.A1(n_494),
.A2(n_510),
.B(n_509),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_479),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_498),
.Y(n_543)
);

AO21x2_ASAP7_75t_L g544 ( 
.A1(n_510),
.A2(n_506),
.B(n_484),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_513),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_512),
.B(n_517),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_489),
.B(n_491),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_495),
.B(n_504),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_480),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_495),
.B(n_504),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_500),
.B(n_516),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_498),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_498),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_514),
.B(n_501),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_492),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_519),
.Y(n_556)
);

AO21x2_ASAP7_75t_L g557 ( 
.A1(n_531),
.A2(n_499),
.B(n_502),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_542),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_542),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_542),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_547),
.B(n_501),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_524),
.B(n_498),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_520),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_524),
.B(n_516),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_516),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_523),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_523),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_516),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_546),
.B(n_477),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_520),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_535),
.B(n_477),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_552),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_534),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_535),
.B(n_522),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_534),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_538),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_530),
.B(n_554),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_538),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_527),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_525),
.B(n_548),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_551),
.B(n_552),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_540),
.B(n_537),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_552),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_530),
.B(n_536),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_548),
.B(n_550),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_533),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_536),
.B(n_541),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_528),
.Y(n_589)
);

NOR2x1_ASAP7_75t_L g590 ( 
.A(n_540),
.B(n_544),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_550),
.B(n_545),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_541),
.B(n_545),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_529),
.B(n_543),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_586),
.B(n_528),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_572),
.B(n_549),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_583),
.B(n_558),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_556),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_586),
.B(n_537),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_583),
.B(n_540),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_585),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_574),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_591),
.B(n_540),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_559),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_544),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_574),
.Y(n_606)
);

NAND2x1p5_ASAP7_75t_L g607 ( 
.A(n_590),
.B(n_532),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_581),
.B(n_544),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_572),
.B(n_582),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_559),
.B(n_544),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_560),
.B(n_531),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_560),
.B(n_531),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_571),
.B(n_526),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_575),
.B(n_532),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_566),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_567),
.B(n_556),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_588),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_561),
.B(n_553),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_576),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_576),
.Y(n_620)
);

NOR2x1p5_ASAP7_75t_L g621 ( 
.A(n_571),
.B(n_543),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_563),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_569),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_575),
.B(n_532),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_563),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_570),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_582),
.B(n_549),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_570),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_609),
.B(n_579),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_602),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_617),
.B(n_566),
.Y(n_631)
);

AND2x4_ASAP7_75t_SL g632 ( 
.A(n_615),
.B(n_587),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_623),
.A2(n_561),
.B1(n_569),
.B2(n_555),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_602),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_604),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_603),
.B(n_590),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_609),
.B(n_577),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_606),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_603),
.B(n_555),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_601),
.B(n_616),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_605),
.B(n_564),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_618),
.B(n_564),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_594),
.B(n_562),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_606),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_605),
.B(n_562),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_609),
.B(n_611),
.Y(n_646)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_598),
.B(n_568),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_594),
.B(n_568),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_619),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_608),
.B(n_580),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_608),
.B(n_580),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_619),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_620),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_620),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_622),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_599),
.B(n_573),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_604),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_614),
.B(n_589),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_625),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_626),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_633),
.A2(n_613),
.B1(n_621),
.B2(n_595),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_660),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_650),
.B(n_610),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_639),
.B(n_600),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_659),
.Y(n_665)
);

NAND2x1p5_ASAP7_75t_L g666 ( 
.A(n_647),
.B(n_610),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_659),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_646),
.B(n_611),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_660),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_655),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_630),
.Y(n_671)
);

NAND2x1_ASAP7_75t_L g672 ( 
.A(n_630),
.B(n_612),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_646),
.B(n_624),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_646),
.B(n_624),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_650),
.B(n_612),
.Y(n_675)
);

NAND2x1p5_ASAP7_75t_L g676 ( 
.A(n_629),
.B(n_596),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_634),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_670),
.B(n_640),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_661),
.A2(n_631),
.B(n_642),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_665),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_661),
.A2(n_637),
.B1(n_629),
.B2(n_627),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_666),
.B(n_629),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_662),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_667),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_673),
.B(n_674),
.Y(n_685)
);

NAND2x1p5_ASAP7_75t_L g686 ( 
.A(n_672),
.B(n_637),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_668),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_671),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_666),
.A2(n_637),
.B1(n_595),
.B2(n_627),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_SL g690 ( 
.A(n_682),
.B(n_587),
.Y(n_690)
);

OAI31xp33_ASAP7_75t_L g691 ( 
.A1(n_686),
.A2(n_676),
.A3(n_632),
.B(n_639),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_678),
.B(n_664),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_681),
.A2(n_689),
.B1(n_679),
.B2(n_687),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_680),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_684),
.B(n_641),
.Y(n_695)
);

OAI32xp33_ASAP7_75t_L g696 ( 
.A1(n_688),
.A2(n_676),
.A3(n_663),
.B1(n_675),
.B2(n_677),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_685),
.B(n_668),
.Y(n_697)
);

OAI21xp33_ASAP7_75t_SL g698 ( 
.A1(n_691),
.A2(n_681),
.B(n_689),
.Y(n_698)
);

AOI211xp5_ASAP7_75t_L g699 ( 
.A1(n_693),
.A2(n_683),
.B(n_669),
.C(n_648),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_696),
.A2(n_656),
.B(n_643),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_694),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_690),
.A2(n_636),
.B1(n_641),
.B2(n_645),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_697),
.A2(n_645),
.B(n_663),
.C(n_675),
.Y(n_703)
);

AOI221xp5_ASAP7_75t_L g704 ( 
.A1(n_699),
.A2(n_695),
.B1(n_692),
.B2(n_636),
.C(n_638),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_701),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_698),
.B(n_632),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_703),
.B(n_651),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_700),
.A2(n_702),
.B(n_649),
.Y(n_708)
);

AND2x2_ASAP7_75t_SL g709 ( 
.A(n_706),
.B(n_584),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_705),
.B(n_652),
.Y(n_710)
);

NOR2x1_ASAP7_75t_L g711 ( 
.A(n_708),
.B(n_592),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_710),
.B(n_707),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_711),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_709),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_SL g715 ( 
.A1(n_711),
.A2(n_704),
.B(n_635),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_714),
.B(n_651),
.Y(n_716)
);

XNOR2xp5_ASAP7_75t_L g717 ( 
.A(n_713),
.B(n_712),
.Y(n_717)
);

XNOR2xp5_ASAP7_75t_L g718 ( 
.A(n_715),
.B(n_584),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_713),
.B(n_654),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_713),
.B(n_653),
.Y(n_720)
);

AOI21xp33_ASAP7_75t_L g721 ( 
.A1(n_717),
.A2(n_526),
.B(n_557),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_719),
.Y(n_722)
);

OAI21x1_ASAP7_75t_SL g723 ( 
.A1(n_720),
.A2(n_533),
.B(n_644),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_716),
.B(n_657),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_718),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_722),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_725),
.A2(n_724),
.B1(n_721),
.B2(n_723),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_724),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_SL g729 ( 
.A(n_722),
.B(n_553),
.C(n_573),
.Y(n_729)
);

OA22x2_ASAP7_75t_L g730 ( 
.A1(n_728),
.A2(n_565),
.B1(n_593),
.B2(n_584),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_726),
.B(n_658),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_729),
.Y(n_732)
);

XNOR2x1_ASAP7_75t_L g733 ( 
.A(n_732),
.B(n_727),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_731),
.A2(n_628),
.B1(n_597),
.B2(n_607),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_730),
.B(n_587),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_734),
.A2(n_733),
.B(n_735),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_736),
.B(n_565),
.Y(n_737)
);

XNOR2xp5_ASAP7_75t_L g738 ( 
.A(n_737),
.B(n_565),
.Y(n_738)
);

AOI21xp33_ASAP7_75t_L g739 ( 
.A1(n_738),
.A2(n_539),
.B(n_543),
.Y(n_739)
);


endmodule