module fake_ibex_1791_n_1134 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1134);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1134;

wire n_1084;
wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_972;
wire n_947;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_959;
wire n_336;
wire n_930;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_1106;
wire n_1129;
wire n_449;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_375;
wire n_317;
wire n_340;
wire n_698;
wire n_901;
wire n_1096;
wire n_187;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_1109;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_1112;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_736;
wire n_550;
wire n_1055;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_641;
wire n_557;
wire n_1103;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1068;
wire n_1057;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_719;
wire n_370;
wire n_431;
wire n_614;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_1082;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_968;
wire n_625;
wire n_953;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_705;
wire n_488;
wire n_1038;
wire n_1092;
wire n_999;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_1126;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1100;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_564;
wire n_506;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_223;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_247;
wire n_379;
wire n_285;
wire n_1128;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_729;
wire n_430;
wire n_414;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1119;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_1095;
wire n_361;
wire n_1085;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_890;
wire n_874;
wire n_912;
wire n_921;
wire n_1058;
wire n_1105;
wire n_677;
wire n_489;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_1000;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_SL g180 ( 
.A(n_74),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_34),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_147),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_41),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_18),
.B(n_178),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_161),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_13),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_63),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_12),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_43),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_140),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_11),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_51),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_49),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_82),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_45),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_29),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_56),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_29),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_94),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_100),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_133),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_12),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_38),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_79),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_23),
.Y(n_216)
);

INVxp33_ASAP7_75t_SL g217 ( 
.A(n_170),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_20),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_65),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_25),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_114),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_25),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_26),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_95),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_16),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_31),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_57),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_85),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_15),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_123),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_72),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_39),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_23),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_13),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_76),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_92),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_15),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_106),
.Y(n_248)
);

BUFx2_ASAP7_75t_SL g249 ( 
.A(n_172),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_168),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_30),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_101),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_99),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_177),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_44),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_86),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_84),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_126),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_26),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_132),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_116),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_137),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_71),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_50),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_98),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_6),
.Y(n_266)
);

INVxp33_ASAP7_75t_SL g267 ( 
.A(n_58),
.Y(n_267)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_36),
.Y(n_268)
);

INVxp33_ASAP7_75t_SL g269 ( 
.A(n_6),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_160),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_27),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_152),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_124),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_144),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_21),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_111),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_96),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_146),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_141),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_143),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_70),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_11),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_139),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_129),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_150),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_119),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_33),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_83),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_35),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_24),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_37),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_31),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_75),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_30),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_120),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_20),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_42),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_145),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_1),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_181),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_283),
.A2(n_197),
.B1(n_291),
.B2(n_269),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_194),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_203),
.B(n_0),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_221),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_207),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_221),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_283),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_203),
.B(n_2),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_231),
.B(n_259),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_191),
.B(n_3),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_210),
.A2(n_215),
.B(n_194),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_212),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_316)
);

NOR2x1_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_185),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_215),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_182),
.Y(n_323)
);

OAI21x1_ASAP7_75t_L g324 ( 
.A1(n_255),
.A2(n_78),
.B(n_176),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_183),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_212),
.B(n_4),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_221),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_261),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_184),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_187),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_261),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_221),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_221),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_268),
.B(n_7),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_188),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_262),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_195),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_8),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_196),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_198),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_8),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_262),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_258),
.B(n_9),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_242),
.Y(n_347)
);

BUFx8_ASAP7_75t_L g348 ( 
.A(n_193),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_213),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_242),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_242),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_216),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_219),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_182),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_222),
.B(n_9),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_258),
.B(n_10),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_199),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_201),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_279),
.B(n_10),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_242),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_226),
.B(n_14),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_222),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g364 ( 
.A(n_230),
.B(n_40),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_233),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_279),
.B(n_14),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_256),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_234),
.B(n_16),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_202),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_204),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_208),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_240),
.B(n_17),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_193),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_286),
.B(n_17),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_237),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_209),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_214),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_218),
.B(n_18),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_256),
.B(n_19),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_220),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_263),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_263),
.B(n_19),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_223),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_241),
.B(n_21),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_224),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_243),
.B(n_22),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_256),
.B(n_22),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_256),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_260),
.B(n_24),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_244),
.B(n_27),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_227),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_228),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_247),
.Y(n_394)
);

BUFx12f_ASAP7_75t_L g395 ( 
.A(n_186),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_323),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_301),
.B(n_186),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_318),
.B(n_229),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_324),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_344),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_314),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_306),
.B(n_320),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_318),
.B(n_235),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_344),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_192),
.Y(n_407)
);

AND2x6_ASAP7_75t_L g408 ( 
.A(n_356),
.B(n_239),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_323),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_395),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_395),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_360),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_345),
.B(n_192),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_307),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_311),
.B(n_211),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_348),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_360),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_376),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_307),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_375),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

OAI22xp33_ASAP7_75t_L g422 ( 
.A1(n_362),
.A2(n_240),
.B1(n_269),
.B2(n_225),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_302),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_325),
.B(n_217),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_325),
.B(n_246),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_304),
.B(n_251),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_304),
.A2(n_238),
.B1(n_190),
.B2(n_236),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_310),
.B(n_349),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_329),
.B(n_217),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_304),
.B(n_275),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_330),
.B(n_267),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_383),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_307),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_307),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_356),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_334),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_356),
.B(n_211),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_335),
.B(n_267),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_335),
.B(n_250),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_337),
.B(n_252),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_337),
.B(n_232),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_355),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_317),
.B(n_282),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_309),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_334),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_339),
.A2(n_316),
.B1(n_375),
.B2(n_373),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_309),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_339),
.B(n_292),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_303),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_340),
.B(n_253),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_340),
.B(n_293),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_303),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_L g459 ( 
.A(n_341),
.B(n_232),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_305),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_357),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_363),
.Y(n_462)
);

NAND2x1p5_ASAP7_75t_L g463 ( 
.A(n_362),
.B(n_353),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_319),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_341),
.Y(n_465)
);

INVx5_ASAP7_75t_L g466 ( 
.A(n_305),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_354),
.B(n_295),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_358),
.B(n_254),
.Y(n_468)
);

AO22x2_ASAP7_75t_L g469 ( 
.A1(n_313),
.A2(n_205),
.B1(n_266),
.B2(n_297),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_365),
.B(n_193),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_358),
.B(n_359),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_359),
.B(n_257),
.Y(n_472)
);

NOR3xp33_ASAP7_75t_L g473 ( 
.A(n_308),
.B(n_342),
.C(n_368),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_373),
.A2(n_190),
.B1(n_206),
.B2(n_236),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_315),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_319),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_370),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_382),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_370),
.B(n_193),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_315),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_394),
.B(n_245),
.Y(n_482)
);

OR2x2_ASAP7_75t_SL g483 ( 
.A(n_385),
.B(n_387),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_309),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_321),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_305),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_315),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_307),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_321),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_371),
.B(n_265),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_364),
.B(n_272),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_379),
.B(n_206),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_371),
.B(n_193),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_328),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_328),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_372),
.B(n_276),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_372),
.B(n_277),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_315),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_377),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_377),
.B(n_378),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_331),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_331),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_336),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_327),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_327),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_336),
.Y(n_506)
);

INVx8_ASAP7_75t_L g507 ( 
.A(n_312),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_378),
.B(n_281),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_381),
.B(n_245),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_381),
.A2(n_249),
.B1(n_294),
.B2(n_284),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_384),
.B(n_285),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_384),
.B(n_287),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_386),
.B(n_296),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_305),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_343),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_322),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_327),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_386),
.B(n_238),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_392),
.B(n_298),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_393),
.B(n_270),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_393),
.B(n_264),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_343),
.B(n_260),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_312),
.B(n_278),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_312),
.B(n_322),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_346),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_346),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_351),
.B(n_274),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_351),
.Y(n_528)
);

NAND3x1_ASAP7_75t_L g529 ( 
.A(n_391),
.B(n_189),
.C(n_32),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_305),
.B(n_278),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_374),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_380),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_463),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_463),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_401),
.B(n_405),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_465),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_481),
.Y(n_537)
);

NOR2x1p5_ASAP7_75t_L g538 ( 
.A(n_425),
.B(n_289),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_402),
.B(n_28),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_411),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_481),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_499),
.B(n_289),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_480),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_498),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_480),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_499),
.B(n_299),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_420),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_400),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_412),
.B(n_388),
.Y(n_551)
);

BUFx12f_ASAP7_75t_L g552 ( 
.A(n_410),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_400),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_399),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_400),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_493),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_523),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_426),
.B(n_299),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_471),
.Y(n_560)
);

BUFx4f_ASAP7_75t_SL g561 ( 
.A(n_427),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_406),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_510),
.A2(n_390),
.B1(n_249),
.B2(n_374),
.Y(n_564)
);

AOI22x1_ASAP7_75t_L g565 ( 
.A1(n_406),
.A2(n_273),
.B1(n_260),
.B2(n_367),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_471),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_516),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_432),
.B(n_434),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_441),
.B(n_180),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

OR2x6_ASAP7_75t_L g571 ( 
.A(n_469),
.B(n_260),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_514),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_477),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_420),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_507),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_521),
.B(n_200),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_406),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_447),
.Y(n_578)
);

AOI211xp5_ASAP7_75t_L g579 ( 
.A1(n_422),
.A2(n_260),
.B(n_273),
.C(n_374),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_518),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_407),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_510),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_423),
.Y(n_583)
);

NOR2x1p5_ASAP7_75t_L g584 ( 
.A(n_431),
.B(n_415),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_520),
.B(n_273),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_469),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_449),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_507),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_467),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_493),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_511),
.B(n_273),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_524),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_511),
.B(n_327),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_439),
.B(n_28),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_474),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_478),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_446),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_475),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_524),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_450),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_451),
.B(n_32),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_507),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_462),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_438),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

AND2x6_ASAP7_75t_SL g607 ( 
.A(n_403),
.B(n_33),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_450),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_475),
.B(n_487),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_408),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_513),
.B(n_327),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_453),
.Y(n_612)
);

CKINVDCx16_ASAP7_75t_R g613 ( 
.A(n_518),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_453),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_501),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_522),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_417),
.B(n_332),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_408),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_408),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_484),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_490),
.B(n_332),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_484),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_455),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_458),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_520),
.B(n_332),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_487),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_435),
.A2(n_350),
.B1(n_367),
.B2(n_361),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_482),
.B(n_333),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_461),
.B(n_333),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_526),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_457),
.B(n_429),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_464),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_408),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_476),
.Y(n_634)
);

NOR2x1p5_ASAP7_75t_L g635 ( 
.A(n_454),
.B(n_34),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_490),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_L g637 ( 
.A(n_430),
.B(n_35),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_527),
.B(n_333),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_457),
.B(n_37),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_492),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_430),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_485),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_489),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_454),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_429),
.B(n_38),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_494),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_527),
.B(n_333),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_495),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_474),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_483),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_452),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_433),
.B(n_333),
.Y(n_652)
);

OR2x2_ASAP7_75t_SL g653 ( 
.A(n_473),
.B(n_39),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_502),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_532),
.B(n_338),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_522),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_433),
.B(n_338),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_503),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_537),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_568),
.B(n_452),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_560),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_566),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_575),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_583),
.B(n_492),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_533),
.B(n_534),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_563),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_598),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_535),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_542),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_597),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_613),
.B(n_541),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_568),
.A2(n_497),
.B(n_443),
.C(n_496),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_536),
.B(n_448),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_549),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_542),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_535),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_549),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_575),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_631),
.B(n_442),
.Y(n_680)
);

AOI222xp33_ASAP7_75t_L g681 ( 
.A1(n_651),
.A2(n_448),
.B1(n_397),
.B2(n_512),
.C1(n_444),
.C2(n_472),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_540),
.B(n_459),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_582),
.A2(n_571),
.B1(n_558),
.B2(n_535),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_570),
.A2(n_440),
.B1(n_398),
.B2(n_404),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_631),
.B(n_413),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_626),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_588),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_571),
.A2(n_500),
.B1(n_491),
.B2(n_528),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_631),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_551),
.B(n_445),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_551),
.B(n_509),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_597),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_545),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_545),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_551),
.B(n_428),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_588),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_626),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_618),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_597),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_618),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_584),
.B(n_442),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_571),
.A2(n_491),
.B1(n_528),
.B2(n_398),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_541),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_618),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_589),
.B(n_428),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_618),
.B(n_396),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_639),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_645),
.A2(n_639),
.B1(n_650),
.B2(n_637),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_602),
.A2(n_491),
.B1(n_404),
.B2(n_468),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_633),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_581),
.B(n_444),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_597),
.Y(n_712)
);

AND3x1_ASAP7_75t_SL g713 ( 
.A(n_635),
.B(n_529),
.C(n_525),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_559),
.B(n_456),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_644),
.B(n_636),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_632),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_559),
.B(n_456),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_586),
.A2(n_639),
.B1(n_641),
.B2(n_649),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_602),
.A2(n_645),
.B1(n_547),
.B2(n_564),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_602),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_645),
.B(n_468),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_552),
.B(n_472),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_629),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_552),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_619),
.A2(n_519),
.B1(n_508),
.B2(n_512),
.Y(n_725)
);

CKINVDCx16_ASAP7_75t_R g726 ( 
.A(n_573),
.Y(n_726)
);

BUFx12f_ASAP7_75t_L g727 ( 
.A(n_607),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_561),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_543),
.B(n_491),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_633),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_R g731 ( 
.A(n_574),
.B(n_506),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_548),
.A2(n_409),
.B1(n_530),
.B2(n_515),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_576),
.B(n_569),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_603),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_561),
.Y(n_735)
);

NOR2x1p5_ASAP7_75t_SL g736 ( 
.A(n_550),
.B(n_553),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_633),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_592),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_599),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_554),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_633),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_603),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_610),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_605),
.B(n_421),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_544),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_632),
.B(n_424),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_634),
.B(n_522),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_544),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_634),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_572),
.Y(n_750)
);

OAI21x1_ASAP7_75t_SL g751 ( 
.A1(n_564),
.A2(n_46),
.B(n_47),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_572),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_652),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_594),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_652),
.Y(n_755)
);

BUFx8_ASAP7_75t_SL g756 ( 
.A(n_595),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_619),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_554),
.B(n_460),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_556),
.B(n_460),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_653),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_539),
.B(n_338),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_623),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_546),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_572),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_572),
.Y(n_765)
);

OR2x6_ASAP7_75t_L g766 ( 
.A(n_610),
.B(n_347),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_621),
.A2(n_436),
.B(n_517),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_619),
.A2(n_531),
.B1(n_460),
.B2(n_466),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_595),
.Y(n_769)
);

OR2x6_ASAP7_75t_L g770 ( 
.A(n_652),
.B(n_347),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_538),
.Y(n_771)
);

INVx5_ASAP7_75t_SL g772 ( 
.A(n_617),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_722),
.B(n_556),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_711),
.B(n_580),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_660),
.A2(n_640),
.B1(n_557),
.B2(n_546),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_703),
.B(n_642),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_683),
.A2(n_658),
.B1(n_642),
.B2(n_646),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_733),
.A2(n_546),
.B1(n_557),
.B2(n_590),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_683),
.A2(n_719),
.B1(n_709),
.B2(n_721),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_719),
.A2(n_658),
.B1(n_646),
.B2(n_654),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_722),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_722),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_733),
.A2(n_557),
.B1(n_585),
.B2(n_643),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_709),
.A2(n_654),
.B1(n_624),
.B2(n_648),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_659),
.Y(n_785)
);

AO31x2_ASAP7_75t_L g786 ( 
.A1(n_673),
.A2(n_585),
.A3(n_555),
.B(n_562),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_762),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_666),
.A2(n_579),
.B1(n_567),
.B2(n_625),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_659),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_770),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_661),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_731),
.Y(n_792)
);

AOI222xp33_ASAP7_75t_L g793 ( 
.A1(n_760),
.A2(n_601),
.B1(n_622),
.B2(n_608),
.C1(n_612),
.C2(n_614),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_681),
.B(n_604),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_SL g795 ( 
.A1(n_672),
.A2(n_609),
.B1(n_591),
.B2(n_606),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_662),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_SL g797 ( 
.A1(n_731),
.A2(n_604),
.B1(n_606),
.B2(n_625),
.Y(n_797)
);

CKINVDCx16_ASAP7_75t_R g798 ( 
.A(n_726),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_705),
.B(n_628),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_724),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_716),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_770),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_721),
.A2(n_702),
.B1(n_717),
.B2(n_714),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_715),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_702),
.A2(n_617),
.B1(n_615),
.B2(n_630),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_669),
.Y(n_806)
);

AOI221xp5_ASAP7_75t_L g807 ( 
.A1(n_718),
.A2(n_620),
.B1(n_638),
.B2(n_647),
.C(n_657),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_688),
.B(n_627),
.C(n_617),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_716),
.Y(n_809)
);

AOI222xp33_ASAP7_75t_SL g810 ( 
.A1(n_675),
.A2(n_630),
.B1(n_615),
.B2(n_596),
.C1(n_587),
.C2(n_578),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_677),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_708),
.A2(n_615),
.B1(n_630),
.B2(n_596),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_728),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_688),
.A2(n_578),
.B1(n_587),
.B2(n_611),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_728),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_718),
.A2(n_657),
.B1(n_593),
.B2(n_655),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_749),
.Y(n_817)
);

AOI211x1_ASAP7_75t_L g818 ( 
.A1(n_684),
.A2(n_627),
.B(n_600),
.C(n_53),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_678),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_720),
.A2(n_577),
.B1(n_562),
.B2(n_600),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_664),
.B(n_600),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_686),
.A2(n_577),
.B(n_565),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_678),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_735),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_707),
.A2(n_600),
.B1(n_656),
.B2(n_616),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_696),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_749),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_696),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_695),
.A2(n_656),
.B1(n_616),
.B2(n_347),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_725),
.A2(n_656),
.B1(n_616),
.B2(n_347),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_686),
.A2(n_347),
.B1(n_350),
.B2(n_352),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_758),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_680),
.B(n_701),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_698),
.B(n_616),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_L g835 ( 
.A1(n_734),
.A2(n_350),
.B1(n_352),
.B2(n_361),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_665),
.B(n_531),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_765),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_SL g838 ( 
.A1(n_706),
.A2(n_48),
.B(n_52),
.C(n_54),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_738),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_668),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_739),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_723),
.A2(n_350),
.B1(n_352),
.B2(n_361),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_670),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_680),
.A2(n_531),
.B1(n_466),
.B2(n_486),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_676),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_769),
.B(n_350),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_665),
.B(n_352),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_693),
.A2(n_517),
.B(n_505),
.Y(n_848)
);

BUFx12f_ASAP7_75t_L g849 ( 
.A(n_727),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_689),
.A2(n_352),
.B1(n_361),
.B2(n_367),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_754),
.Y(n_851)
);

AOI222xp33_ASAP7_75t_L g852 ( 
.A1(n_674),
.A2(n_361),
.B1(n_367),
.B2(n_369),
.C1(n_486),
.C2(n_466),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_765),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_693),
.A2(n_486),
.B(n_369),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_770),
.Y(n_855)
);

NAND2x1_ASAP7_75t_L g856 ( 
.A(n_766),
.B(n_367),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_SL g857 ( 
.A1(n_771),
.A2(n_369),
.B1(n_59),
.B2(n_60),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_758),
.Y(n_858)
);

INVx8_ASAP7_75t_L g859 ( 
.A(n_700),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_690),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_691),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_729),
.A2(n_369),
.B(n_504),
.C(n_488),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_698),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_685),
.A2(n_756),
.B1(n_755),
.B2(n_753),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_772),
.A2(n_734),
.B1(n_742),
.B2(n_753),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_679),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_744),
.A2(n_505),
.B1(n_504),
.B2(n_488),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_761),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_772),
.A2(n_505),
.B1(n_504),
.B2(n_488),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_745),
.Y(n_870)
);

OAI221xp5_ASAP7_75t_SL g871 ( 
.A1(n_682),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.C(n_64),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_742),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_748),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_679),
.Y(n_874)
);

OAI22x1_ASAP7_75t_L g875 ( 
.A1(n_713),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_875)
);

AOI222xp33_ASAP7_75t_L g876 ( 
.A1(n_740),
.A2(n_437),
.B1(n_436),
.B2(n_419),
.C1(n_414),
.C2(n_81),
.Y(n_876)
);

BUFx12f_ASAP7_75t_L g877 ( 
.A(n_759),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_SL g878 ( 
.A1(n_772),
.A2(n_437),
.B1(n_419),
.B2(n_414),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_763),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_SL g880 ( 
.A1(n_751),
.A2(n_437),
.B1(n_419),
.B2(n_77),
.Y(n_880)
);

CKINVDCx11_ASAP7_75t_R g881 ( 
.A(n_663),
.Y(n_881)
);

BUFx4f_ASAP7_75t_L g882 ( 
.A(n_750),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_755),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_744),
.A2(n_69),
.B1(n_73),
.B2(n_80),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_756),
.A2(n_663),
.B1(n_687),
.B2(n_750),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_687),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_746),
.A2(n_764),
.B1(n_752),
.B2(n_694),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_752),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_698),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_764),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_759),
.B(n_87),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_712),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_757),
.B(n_88),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_700),
.Y(n_894)
);

BUFx2_ASAP7_75t_L g895 ( 
.A(n_712),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_732),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_700),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_671),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_671),
.B(n_89),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_833),
.B(n_692),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_787),
.Y(n_901)
);

OAI22xp33_ASAP7_75t_L g902 ( 
.A1(n_792),
.A2(n_713),
.B1(n_757),
.B2(n_700),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_896),
.A2(n_736),
.B(n_692),
.C(n_699),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_859),
.Y(n_904)
);

AOI221xp5_ASAP7_75t_L g905 ( 
.A1(n_803),
.A2(n_699),
.B1(n_747),
.B2(n_730),
.C(n_768),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_851),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_791),
.Y(n_907)
);

OAI221xp5_ASAP7_75t_L g908 ( 
.A1(n_794),
.A2(n_730),
.B1(n_766),
.B2(n_743),
.C(n_667),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_781),
.B(n_704),
.Y(n_909)
);

HB1xp67_ASAP7_75t_L g910 ( 
.A(n_804),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_796),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_773),
.B(n_704),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_774),
.B(n_704),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_779),
.A2(n_697),
.B1(n_743),
.B2(n_766),
.Y(n_914)
);

AOI221xp5_ASAP7_75t_L g915 ( 
.A1(n_860),
.A2(n_861),
.B1(n_839),
.B2(n_841),
.C(n_807),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_776),
.B(n_743),
.Y(n_916)
);

OAI211xp5_ASAP7_75t_L g917 ( 
.A1(n_864),
.A2(n_767),
.B(n_741),
.C(n_737),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_807),
.B(n_741),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_819),
.A2(n_816),
.B1(n_782),
.B2(n_797),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_798),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_806),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_811),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_816),
.A2(n_741),
.B1(n_737),
.B2(n_710),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_SL g924 ( 
.A1(n_782),
.A2(n_710),
.B1(n_698),
.B2(n_97),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_859),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_785),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_780),
.A2(n_710),
.B1(n_93),
.B2(n_102),
.Y(n_927)
);

AOI221xp5_ASAP7_75t_L g928 ( 
.A1(n_783),
.A2(n_91),
.B1(n_103),
.B2(n_104),
.C(n_105),
.Y(n_928)
);

OAI221xp5_ASAP7_75t_L g929 ( 
.A1(n_775),
.A2(n_108),
.B1(n_110),
.B2(n_113),
.C(n_117),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_883),
.Y(n_930)
);

OAI211xp5_ASAP7_75t_L g931 ( 
.A1(n_793),
.A2(n_118),
.B(n_125),
.C(n_127),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_872),
.B(n_128),
.Y(n_932)
);

AOI221xp5_ASAP7_75t_SL g933 ( 
.A1(n_783),
.A2(n_142),
.B1(n_149),
.B2(n_151),
.C(n_153),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_810),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_934)
);

OAI221xp5_ASAP7_75t_L g935 ( 
.A1(n_775),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.C(n_164),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_826),
.Y(n_936)
);

AOI221xp5_ASAP7_75t_L g937 ( 
.A1(n_784),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.C(n_174),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_828),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_822),
.A2(n_175),
.B(n_179),
.Y(n_939)
);

AOI221xp5_ASAP7_75t_L g940 ( 
.A1(n_778),
.A2(n_777),
.B1(n_823),
.B2(n_868),
.C(n_885),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_872),
.A2(n_799),
.B1(n_887),
.B2(n_865),
.Y(n_941)
);

OAI221xp5_ASAP7_75t_L g942 ( 
.A1(n_778),
.A2(n_788),
.B1(n_773),
.B2(n_824),
.C(n_846),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_870),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_773),
.B(n_813),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_800),
.B(n_832),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_887),
.A2(n_871),
.B1(n_855),
.B2(n_790),
.Y(n_946)
);

AOI222xp33_ASAP7_75t_L g947 ( 
.A1(n_875),
.A2(n_849),
.B1(n_881),
.B2(n_877),
.C1(n_858),
.C2(n_857),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_873),
.Y(n_948)
);

OAI222xp33_ASAP7_75t_L g949 ( 
.A1(n_871),
.A2(n_795),
.B1(n_884),
.B2(n_866),
.C1(n_880),
.C2(n_805),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_790),
.A2(n_855),
.B1(n_802),
.B2(n_878),
.Y(n_950)
);

OAI211xp5_ASAP7_75t_SL g951 ( 
.A1(n_852),
.A2(n_815),
.B(n_890),
.C(n_888),
.Y(n_951)
);

OAI221xp5_ASAP7_75t_L g952 ( 
.A1(n_880),
.A2(n_795),
.B1(n_812),
.B2(n_884),
.C(n_847),
.Y(n_952)
);

OAI22xp33_ASAP7_75t_L g953 ( 
.A1(n_882),
.A2(n_874),
.B1(n_859),
.B2(n_802),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_821),
.A2(n_891),
.B1(n_836),
.B2(n_874),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_837),
.A2(n_853),
.B1(n_886),
.B2(n_808),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_837),
.A2(n_853),
.B1(n_886),
.B2(n_879),
.Y(n_956)
);

AOI222xp33_ASAP7_75t_L g957 ( 
.A1(n_882),
.A2(n_827),
.B1(n_817),
.B2(n_801),
.C1(n_809),
.C2(n_814),
.Y(n_957)
);

AO31x2_ASAP7_75t_L g958 ( 
.A1(n_862),
.A2(n_830),
.A3(n_820),
.B(n_848),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_789),
.B(n_843),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_SL g960 ( 
.A1(n_893),
.A2(n_835),
.B(n_831),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_840),
.B(n_845),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_SL g962 ( 
.A1(n_897),
.A2(n_894),
.B1(n_892),
.B2(n_895),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_898),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_876),
.A2(n_897),
.B1(n_844),
.B2(n_899),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_863),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_786),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_848),
.A2(n_831),
.B(n_854),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_786),
.B(n_818),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_878),
.A2(n_842),
.B1(n_867),
.B2(n_829),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_863),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_829),
.A2(n_842),
.B1(n_825),
.B2(n_889),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_786),
.B(n_825),
.Y(n_972)
);

AOI221xp5_ASAP7_75t_L g973 ( 
.A1(n_838),
.A2(n_869),
.B1(n_867),
.B2(n_850),
.C(n_856),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_786),
.Y(n_974)
);

AOI21xp33_ASAP7_75t_L g975 ( 
.A1(n_834),
.A2(n_863),
.B(n_889),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_889),
.A2(n_733),
.B(n_673),
.C(n_717),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_779),
.A2(n_760),
.B1(n_651),
.B2(n_641),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_785),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_896),
.A2(n_733),
.B(n_673),
.C(n_717),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_919),
.A2(n_979),
.B1(n_941),
.B2(n_977),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_926),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_941),
.A2(n_964),
.B1(n_942),
.B2(n_934),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_SL g983 ( 
.A1(n_950),
.A2(n_946),
.B1(n_931),
.B2(n_944),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_912),
.B(n_916),
.Y(n_984)
);

AO21x2_ASAP7_75t_L g985 ( 
.A1(n_968),
.A2(n_972),
.B(n_967),
.Y(n_985)
);

OAI221xp5_ASAP7_75t_L g986 ( 
.A1(n_940),
.A2(n_976),
.B1(n_915),
.B2(n_954),
.C(n_947),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_910),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_920),
.B(n_945),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_944),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_959),
.B(n_978),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_961),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_947),
.A2(n_951),
.B1(n_946),
.B2(n_900),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_936),
.B(n_938),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_950),
.A2(n_952),
.B1(n_960),
.B2(n_962),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_901),
.B(n_911),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_907),
.B(n_906),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_943),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_957),
.A2(n_913),
.B1(n_912),
.B2(n_904),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_904),
.B(n_965),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_925),
.Y(n_1000)
);

OAI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_914),
.A2(n_933),
.B1(n_955),
.B2(n_930),
.C(n_922),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_921),
.B(n_948),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_966),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_974),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_963),
.Y(n_1005)
);

OAI31xp33_ASAP7_75t_L g1006 ( 
.A1(n_949),
.A2(n_902),
.A3(n_953),
.B(n_969),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_918),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_965),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_903),
.A2(n_927),
.B(n_969),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_L g1010 ( 
.A(n_957),
.B(n_928),
.C(n_937),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_970),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_925),
.A2(n_909),
.B1(n_927),
.B2(n_956),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_909),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_929),
.A2(n_935),
.B1(n_905),
.B2(n_908),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_958),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_932),
.A2(n_924),
.B1(n_971),
.B2(n_923),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_917),
.B(n_939),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_958),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_L g1019 ( 
.A(n_973),
.B(n_975),
.C(n_958),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_979),
.B(n_651),
.Y(n_1020)
);

NOR4xp25_ASAP7_75t_L g1021 ( 
.A(n_979),
.B(n_718),
.C(n_529),
.D(n_977),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_SL g1022 ( 
.A1(n_950),
.A2(n_518),
.B1(n_613),
.B2(n_672),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_965),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_979),
.B(n_651),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_959),
.B(n_926),
.Y(n_1025)
);

AO21x2_ASAP7_75t_L g1026 ( 
.A1(n_968),
.A2(n_972),
.B(n_967),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_926),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1003),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1003),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_SL g1030 ( 
.A1(n_1022),
.A2(n_983),
.B(n_992),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1004),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1004),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_980),
.A2(n_982),
.B1(n_986),
.B2(n_1020),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1007),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_990),
.B(n_1025),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_1023),
.B(n_1013),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_993),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_990),
.B(n_1025),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_1023),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_1023),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_997),
.B(n_1005),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1024),
.B(n_1007),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_988),
.B(n_989),
.Y(n_1043)
);

AO21x2_ASAP7_75t_L g1044 ( 
.A1(n_1009),
.A2(n_1019),
.B(n_1018),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_L g1045 ( 
.A(n_1013),
.B(n_994),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_991),
.B(n_981),
.Y(n_1046)
);

NOR2x1p5_ASAP7_75t_L g1047 ( 
.A(n_1023),
.B(n_1015),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_1023),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_SL g1049 ( 
.A(n_998),
.B(n_1000),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1027),
.B(n_1026),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1027),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_985),
.B(n_1026),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_985),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_995),
.B(n_985),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_1014),
.A2(n_1010),
.B1(n_1012),
.B2(n_1001),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_1035),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_1048),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1050),
.B(n_1031),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1035),
.B(n_995),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1032),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_1040),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1032),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1028),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1050),
.B(n_1038),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1028),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_1054),
.B(n_1026),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1038),
.B(n_984),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_R g1068 ( 
.A(n_1049),
.B(n_1000),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_L g1069 ( 
.A(n_1030),
.B(n_987),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1029),
.Y(n_1070)
);

INVxp33_ASAP7_75t_L g1071 ( 
.A(n_1068),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_1064),
.B(n_1054),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_1064),
.B(n_1052),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1058),
.B(n_1052),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1056),
.B(n_1053),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1063),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1062),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1059),
.B(n_1041),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1058),
.B(n_1041),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_1061),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1063),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1067),
.B(n_1070),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_1061),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1065),
.Y(n_1084)
);

OAI321xp33_ASAP7_75t_L g1085 ( 
.A1(n_1083),
.A2(n_1055),
.A3(n_1033),
.B1(n_1066),
.B2(n_1037),
.C(n_1036),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1077),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_1075),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1076),
.Y(n_1088)
);

XNOR2xp5_ASAP7_75t_L g1089 ( 
.A(n_1071),
.B(n_1069),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1083),
.A2(n_1030),
.B1(n_1055),
.B2(n_1033),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1076),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1074),
.B(n_1067),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1080),
.A2(n_1045),
.B(n_1006),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_1072),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1074),
.B(n_1070),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1082),
.B(n_1065),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1072),
.B(n_1066),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_1089),
.B(n_1085),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1088),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1090),
.A2(n_1089),
.B1(n_1093),
.B2(n_1045),
.Y(n_1101)
);

OAI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_1087),
.A2(n_1021),
.B1(n_1043),
.B2(n_1073),
.C(n_1075),
.Y(n_1102)
);

AOI31xp33_ASAP7_75t_L g1103 ( 
.A1(n_1092),
.A2(n_999),
.A3(n_1073),
.B(n_1036),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1087),
.B(n_1079),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1091),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1087),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1097),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1086),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_L g1109 ( 
.A(n_1086),
.B(n_1047),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1100),
.Y(n_1110)
);

OAI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1103),
.A2(n_1078),
.B1(n_1096),
.B2(n_1057),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1104),
.B(n_1057),
.Y(n_1112)
);

XNOR2xp5_ASAP7_75t_L g1113 ( 
.A(n_1101),
.B(n_1047),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1099),
.A2(n_1081),
.B1(n_1084),
.B2(n_1044),
.Y(n_1114)
);

NAND4xp75_ASAP7_75t_L g1115 ( 
.A(n_1109),
.B(n_1053),
.C(n_1084),
.D(n_1042),
.Y(n_1115)
);

NAND4xp25_ASAP7_75t_L g1116 ( 
.A(n_1114),
.B(n_1102),
.C(n_1098),
.D(n_1107),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1110),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1113),
.A2(n_1106),
.B1(n_1104),
.B2(n_1105),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1111),
.A2(n_1106),
.B1(n_1057),
.B2(n_1108),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1111),
.A2(n_1112),
.B(n_1108),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_SL g1121 ( 
.A(n_1119),
.B(n_999),
.C(n_1036),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_L g1122 ( 
.A(n_1116),
.B(n_1115),
.Y(n_1122)
);

AOI211xp5_ASAP7_75t_L g1123 ( 
.A1(n_1120),
.A2(n_1042),
.B(n_1051),
.C(n_1057),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1118),
.A2(n_1044),
.B1(n_1029),
.B2(n_984),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1122),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1123),
.A2(n_1117),
.B1(n_1016),
.B2(n_1077),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1124),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1125),
.A2(n_1121),
.B1(n_999),
.B2(n_1034),
.Y(n_1128)
);

OAI222xp33_ASAP7_75t_L g1129 ( 
.A1(n_1127),
.A2(n_1017),
.B1(n_996),
.B2(n_1040),
.C1(n_1002),
.C2(n_1051),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1126),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1130),
.A2(n_1034),
.B1(n_1046),
.B2(n_1060),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1131),
.A2(n_1128),
.B1(n_1129),
.B2(n_1046),
.Y(n_1132)
);

OAI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1132),
.A2(n_1017),
.B1(n_1039),
.B2(n_1048),
.Y(n_1133)
);

AOI221xp5_ASAP7_75t_L g1134 ( 
.A1(n_1133),
.A2(n_1008),
.B1(n_984),
.B2(n_1039),
.C(n_1011),
.Y(n_1134)
);


endmodule