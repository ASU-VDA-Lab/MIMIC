module fake_jpeg_6700_n_178 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_1),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_27),
.B1(n_28),
.B2(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_27),
.B1(n_28),
.B2(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_51),
.Y(n_54)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_50),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_22),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_32),
.C(n_35),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_72),
.B(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_66),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_51),
.B1(n_49),
.B2(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_70),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_30),
.B1(n_35),
.B2(n_34),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_49),
.B1(n_34),
.B2(n_26),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_30),
.B1(n_34),
.B2(n_19),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_14),
.B1(n_20),
.B2(n_26),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_30),
.C(n_33),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_21),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_83),
.B1(n_14),
.B2(n_20),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_17),
.B(n_33),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_82),
.A3(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_85),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_86),
.B1(n_73),
.B2(n_69),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_33),
.A3(n_48),
.B1(n_50),
.B2(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_48),
.B1(n_25),
.B2(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_92),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_25),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_85),
.B1(n_88),
.B2(n_87),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_75),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_111),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_58),
.B1(n_72),
.B2(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_77),
.B(n_80),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_81),
.A2(n_65),
.B1(n_56),
.B2(n_57),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_16),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_82),
.B1(n_93),
.B2(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_114),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_20),
.B1(n_14),
.B2(n_22),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_84),
.B(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_126),
.B(n_111),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_118),
.B(n_119),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_92),
.B(n_90),
.Y(n_118)
);

NOR2xp67_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_78),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_99),
.B1(n_97),
.B2(n_103),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_17),
.CI(n_22),
.CON(n_121),
.SN(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_125),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_19),
.B1(n_63),
.B2(n_5),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_16),
.B(n_24),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_3),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_13),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_16),
.B(n_63),
.Y(n_126)
);

AOI221xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_101),
.B1(n_104),
.B2(n_102),
.C(n_105),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_16),
.C(n_4),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_97),
.C(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_135),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_125),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_139),
.C(n_141),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_108),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_143),
.C(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_3),
.C(n_4),
.Y(n_143)
);

OAI322xp33_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_115),
.A3(n_116),
.B1(n_128),
.B2(n_117),
.C1(n_121),
.C2(n_118),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_151),
.B1(n_7),
.B2(n_8),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_144),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_126),
.C(n_129),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_143),
.C(n_140),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_124),
.C(n_121),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_150),
.A2(n_9),
.B(n_10),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_127),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_3),
.B(n_4),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_9),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_156),
.C(n_150),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_146),
.A2(n_136),
.B1(n_6),
.B2(n_7),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_160),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_136),
.C(n_6),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_5),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_12),
.B(n_9),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_161),
.B(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_165),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_166),
.B(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_162),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_11),
.B(n_12),
.Y(n_171)
);

NAND2x1_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_11),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_166),
.C(n_170),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_172),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.Y(n_178)
);


endmodule