module fake_aes_8398_n_24 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_24);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
NOR2xp67_ASAP7_75t_L g12 ( .A(n_7), .B(n_1), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_10), .B(n_5), .Y(n_15) );
INVx4_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_14), .B(n_0), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
NAND3xp33_ASAP7_75t_SL g19 ( .A(n_18), .B(n_11), .C(n_13), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_17), .B(n_12), .Y(n_20) );
NAND3xp33_ASAP7_75t_L g21 ( .A(n_20), .B(n_15), .C(n_0), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_22), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_4), .B1(n_6), .B2(n_8), .Y(n_24) );
endmodule