module fake_jpeg_26795_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

MAJIxp5_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_2),
.C(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx4_ASAP7_75t_SL g11 ( 
.A(n_2),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_16),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_10),
.B(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_3),
.B1(n_4),
.B2(n_13),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_21),
.B1(n_8),
.B2(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_4),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_8),
.B(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_12),
.B1(n_11),
.B2(n_7),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_24),
.B(n_17),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_21),
.B1(n_20),
.B2(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_30),
.B(n_32),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_16),
.B1(n_22),
.B2(n_19),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_40),
.C(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_14),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_45),
.Y(n_47)
);


endmodule