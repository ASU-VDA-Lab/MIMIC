module fake_jpeg_13834_n_576 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_576);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_576;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_10),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_56),
.B(n_61),
.Y(n_149)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_62),
.B(n_63),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_18),
.B(n_8),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_18),
.B(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_66),
.B(n_70),
.Y(n_163)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g167 ( 
.A(n_72),
.Y(n_167)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_76),
.B(n_78),
.Y(n_171)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_77),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_28),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_21),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_82),
.B(n_95),
.Y(n_178)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_90),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_44),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_98),
.B(n_106),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_101),
.Y(n_170)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_17),
.Y(n_103)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_29),
.B(n_8),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_107),
.B(n_113),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_47),
.Y(n_113)
);

OR2x2_ASAP7_75t_SL g114 ( 
.A(n_56),
.B(n_30),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_114),
.B(n_49),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_33),
.B1(n_52),
.B2(n_54),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_115),
.A2(n_138),
.B1(n_90),
.B2(n_112),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_52),
.B1(n_42),
.B2(n_54),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_126),
.A2(n_23),
.B1(n_94),
.B2(n_93),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_29),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_127),
.B(n_23),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_130),
.B(n_158),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_59),
.A2(n_54),
.B1(n_42),
.B2(n_28),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_131),
.A2(n_168),
.B1(n_40),
.B2(n_50),
.Y(n_238)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_84),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_132),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_73),
.B(n_20),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_140),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_75),
.A2(n_33),
.B1(n_42),
.B2(n_35),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_20),
.Y(n_140)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_75),
.Y(n_142)
);

CKINVDCx6p67_ASAP7_75t_R g192 ( 
.A(n_142),
.Y(n_192)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_96),
.A2(n_110),
.B1(n_102),
.B2(n_100),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_154),
.A2(n_68),
.B1(n_104),
.B2(n_69),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_20),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_72),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_86),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_80),
.A2(n_43),
.B1(n_50),
.B2(n_31),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_103),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_60),
.Y(n_181)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_64),
.Y(n_184)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_65),
.Y(n_185)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_188),
.Y(n_281)
);

CKINVDCx12_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_189),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_191),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_193),
.A2(n_219),
.B1(n_74),
.B2(n_177),
.Y(n_269)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g289 ( 
.A(n_194),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_195),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_197),
.B(n_204),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_198),
.B(n_200),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_199),
.B(n_201),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_140),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_92),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_99),
.B1(n_97),
.B2(n_58),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_138),
.C(n_115),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_178),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g308 ( 
.A(n_205),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_43),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_206),
.B(n_210),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_207),
.A2(n_225),
.B1(n_177),
.B2(n_123),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_208),
.B(n_209),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_159),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_34),
.Y(n_210)
);

CKINVDCx12_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_211),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_120),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_212),
.B(n_216),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_214),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_34),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_215),
.B(n_218),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_153),
.B(n_47),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_135),
.Y(n_217)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_31),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_30),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_222),
.B(n_226),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_131),
.A2(n_91),
.B1(n_87),
.B2(n_79),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_224),
.A2(n_118),
.B1(n_133),
.B2(n_124),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_125),
.A2(n_35),
.B1(n_37),
.B2(n_55),
.Y(n_225)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_134),
.B(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_231),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_136),
.B(n_40),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_232),
.B(n_242),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_235),
.Y(n_273)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_147),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_237),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_48),
.B1(n_123),
.B2(n_118),
.Y(n_263)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_148),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_162),
.Y(n_241)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_151),
.B(n_55),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_116),
.Y(n_243)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_116),
.Y(n_244)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_132),
.Y(n_247)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

INVx11_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_164),
.B(n_49),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_251),
.B(n_20),
.Y(n_270)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_173),
.B(n_48),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_150),
.Y(n_252)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_252),
.Y(n_306)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_117),
.Y(n_253)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_129),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_255),
.B(n_257),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_190),
.B(n_213),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_258),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_154),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_259),
.B(n_266),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_260),
.B(n_105),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_263),
.A2(n_192),
.B1(n_240),
.B2(n_245),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_234),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_269),
.A2(n_271),
.B1(n_305),
.B2(n_240),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_270),
.B(n_223),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_226),
.A2(n_154),
.B(n_167),
.C(n_174),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_274),
.B(n_294),
.Y(n_344)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_228),
.B(n_141),
.CI(n_144),
.CON(n_277),
.SN(n_277)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_285),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_228),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_230),
.B(n_196),
.C(n_227),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_286),
.B(n_298),
.C(n_195),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_207),
.A2(n_139),
.B1(n_170),
.B2(n_121),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_236),
.B(n_124),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_192),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_223),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_203),
.B(n_170),
.C(n_139),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_221),
.B(n_133),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_300),
.B(n_235),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_219),
.A2(n_137),
.B1(n_143),
.B2(n_119),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_187),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_314),
.B(n_256),
.C(n_278),
.Y(n_394)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_280),
.Y(n_315)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_317),
.A2(n_357),
.B(n_358),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_192),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_321),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_275),
.B(n_303),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_324),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_294),
.Y(n_321)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_323),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_309),
.B(n_287),
.Y(n_324)
);

BUFx12_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_325),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_301),
.B(n_217),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_326),
.B(n_335),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_259),
.A2(n_193),
.B1(n_224),
.B2(n_225),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_327),
.A2(n_340),
.B1(n_308),
.B2(n_289),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_329),
.A2(n_349),
.B1(n_353),
.B2(n_355),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_330),
.A2(n_345),
.B1(n_347),
.B2(n_350),
.Y(n_391)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_332),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_309),
.B(n_250),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_336),
.Y(n_366)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_223),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_255),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_276),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_247),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_342),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_260),
.A2(n_137),
.B1(n_244),
.B2(n_243),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_302),
.B(n_241),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_343),
.B(n_351),
.Y(n_396)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_348),
.Y(n_368)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_267),
.Y(n_347)
);

INVx13_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_191),
.Y(n_349)
);

BUFx8_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_352),
.A2(n_268),
.B1(n_261),
.B2(n_265),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_288),
.B(n_237),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_292),
.A2(n_205),
.B1(n_220),
.B2(n_253),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_292),
.A2(n_248),
.B(n_152),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_356),
.A2(n_268),
.B(n_288),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_256),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_277),
.B(n_194),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_361),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_274),
.A2(n_147),
.B(n_169),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_360),
.A2(n_293),
.B(n_296),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_277),
.B(n_0),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_344),
.A2(n_298),
.B1(n_271),
.B2(n_282),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_364),
.A2(n_375),
.B1(n_385),
.B2(n_386),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_370),
.A2(n_374),
.B1(n_379),
.B2(n_383),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_327),
.A2(n_282),
.B1(n_273),
.B2(n_289),
.Y(n_374)
);

OAI22x1_ASAP7_75t_SL g375 ( 
.A1(n_329),
.A2(n_268),
.B1(n_280),
.B2(n_310),
.Y(n_375)
);

OA22x2_ASAP7_75t_L g378 ( 
.A1(n_344),
.A2(n_295),
.B1(n_306),
.B2(n_284),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_378),
.B(n_380),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_323),
.B1(n_321),
.B2(n_336),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_341),
.A2(n_273),
.B1(n_299),
.B2(n_265),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_341),
.A2(n_316),
.B1(n_359),
.B2(n_357),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_331),
.A2(n_299),
.B1(n_202),
.B2(n_188),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_357),
.A2(n_295),
.B1(n_261),
.B2(n_306),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_328),
.A2(n_284),
.B1(n_281),
.B2(n_291),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_387),
.A2(n_399),
.B1(n_402),
.B2(n_354),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_314),
.B(n_311),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_389),
.B(n_400),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_311),
.C(n_293),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_356),
.C(n_345),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_392),
.A2(n_395),
.B(n_354),
.Y(n_433)
);

XNOR2x1_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_350),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_360),
.A2(n_296),
.B(n_304),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_328),
.A2(n_291),
.B1(n_281),
.B2(n_233),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_331),
.B(n_333),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g401 ( 
.A1(n_361),
.A2(n_278),
.A3(n_214),
.B1(n_310),
.B2(n_304),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_330),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_346),
.A2(n_176),
.B1(n_117),
.B2(n_37),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_397),
.Y(n_403)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_404),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_405),
.A2(n_421),
.B1(n_434),
.B2(n_374),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_365),
.B(n_319),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_406),
.B(n_408),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_372),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_407),
.B(n_414),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_368),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_324),
.Y(n_410)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_398),
.Y(n_411)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_411),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_396),
.B(n_343),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_415),
.C(n_417),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_372),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_342),
.C(n_334),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_397),
.Y(n_418)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_418),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_320),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_425),
.C(n_429),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_347),
.Y(n_420)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_420),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_368),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_428),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_365),
.B(n_332),
.Y(n_423)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_369),
.B(n_332),
.Y(n_424)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_424),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_389),
.B(n_339),
.C(n_358),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_363),
.B(n_352),
.Y(n_426)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_426),
.Y(n_465)
);

CKINVDCx12_ASAP7_75t_R g427 ( 
.A(n_362),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_427),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_368),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_318),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_383),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_378),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_425),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_433),
.A2(n_392),
.B(n_391),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_315),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_394),
.B(n_325),
.C(n_348),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_386),
.C(n_388),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_409),
.A2(n_364),
.B1(n_393),
.B2(n_375),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_442),
.A2(n_449),
.B1(n_450),
.B2(n_454),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_443),
.A2(n_464),
.B1(n_468),
.B2(n_37),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_407),
.A2(n_370),
.B1(n_379),
.B2(n_384),
.Y(n_444)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_444),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_414),
.A2(n_421),
.B1(n_412),
.B2(n_409),
.Y(n_446)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_446),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_435),
.A2(n_367),
.B1(n_377),
.B2(n_368),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_416),
.A2(n_366),
.B1(n_371),
.B2(n_385),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_416),
.A2(n_366),
.B1(n_378),
.B2(n_401),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_388),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_440),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_432),
.C(n_417),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_431),
.A2(n_378),
.B1(n_395),
.B2(n_402),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_458),
.A2(n_350),
.B1(n_325),
.B2(n_176),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_430),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_462),
.A2(n_12),
.B(n_2),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_403),
.B(n_418),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_463),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_412),
.A2(n_387),
.B1(n_399),
.B2(n_382),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_466),
.B(n_436),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_430),
.A2(n_382),
.B1(n_380),
.B2(n_398),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_433),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_469),
.B(n_470),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_404),
.Y(n_470)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_471),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_411),
.Y(n_472)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_472),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_441),
.B(n_429),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_473),
.A2(n_478),
.B1(n_483),
.B2(n_487),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_474),
.B(n_479),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_477),
.C(n_482),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_415),
.C(n_436),
.Y(n_477)
);

OAI22x1_ASAP7_75t_L g478 ( 
.A1(n_454),
.A2(n_422),
.B1(n_428),
.B2(n_419),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_440),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_481),
.B(n_3),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_451),
.B(n_437),
.C(n_325),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_348),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_484),
.A2(n_490),
.B1(n_438),
.B2(n_491),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_350),
.C(n_108),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_494),
.C(n_0),
.Y(n_513)
);

NOR3xp33_ASAP7_75t_L g487 ( 
.A(n_448),
.B(n_12),
.C(n_2),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_488),
.A2(n_463),
.B(n_459),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_445),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_445),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_491),
.A2(n_438),
.B1(n_467),
.B2(n_447),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_492),
.A2(n_458),
.B1(n_439),
.B2(n_467),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_455),
.B(n_37),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_449),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_35),
.C(n_0),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_492),
.A2(n_453),
.B1(n_442),
.B2(n_448),
.Y(n_498)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_498),
.Y(n_521)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_499),
.Y(n_526)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_501),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_482),
.A2(n_460),
.B(n_452),
.Y(n_502)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_502),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_479),
.B(n_450),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_503),
.B(n_504),
.Y(n_520)
);

INVxp33_ASAP7_75t_SL g505 ( 
.A(n_469),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_469),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_506),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_508),
.A2(n_510),
.B(n_488),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_480),
.A2(n_485),
.B1(n_476),
.B2(n_464),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_509),
.A2(n_513),
.B1(n_495),
.B2(n_508),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_489),
.A2(n_468),
.B1(n_2),
.B2(n_3),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_513),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_11),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_514),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_474),
.B(n_475),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_516),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_3),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_518),
.A2(n_503),
.B(n_504),
.Y(n_534)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_519),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_491),
.Y(n_522)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_522),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_494),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_527),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_499),
.B(n_485),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_530),
.A2(n_521),
.B1(n_518),
.B2(n_529),
.Y(n_540)
);

AO21x1_ASAP7_75t_L g531 ( 
.A1(n_505),
.A2(n_478),
.B(n_486),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_531),
.A2(n_496),
.B1(n_493),
.B2(n_7),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_512),
.B(n_490),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_515),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_536),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_519),
.A2(n_500),
.B(n_514),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_516),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_537),
.B(n_539),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_524),
.B(n_500),
.C(n_496),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_541),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_542),
.B(n_517),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_529),
.A2(n_4),
.B1(n_5),
.B2(n_11),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_543),
.B(n_544),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_4),
.C(n_12),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_520),
.B(n_4),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_546),
.B(n_547),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_520),
.B(n_13),
.C(n_14),
.Y(n_547)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_549),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_531),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_551),
.B(n_552),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_533),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_SL g556 ( 
.A(n_535),
.B(n_522),
.C(n_527),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_556),
.A2(n_557),
.B(n_526),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_523),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_545),
.Y(n_558)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_558),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_549),
.B(n_526),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_560),
.A2(n_562),
.B(n_564),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_534),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_563),
.A2(n_542),
.B1(n_556),
.B2(n_547),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_555),
.B(n_539),
.C(n_546),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_565),
.Y(n_570)
);

AOI322xp5_ASAP7_75t_L g566 ( 
.A1(n_561),
.A2(n_554),
.A3(n_543),
.B1(n_548),
.B2(n_544),
.C1(n_525),
.C2(n_16),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_566),
.B(n_559),
.C(n_563),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_569),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_570),
.C(n_567),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_568),
.B(n_564),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_573),
.A2(n_525),
.B(n_14),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_13),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_15),
.Y(n_576)
);


endmodule