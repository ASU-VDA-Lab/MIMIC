module fake_netlist_1_9054_n_1253 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1253);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1253;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_271;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_272;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_710;
wire n_270;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_269;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g269 ( .A(n_77), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_58), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_187), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_19), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_223), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_161), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_2), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_120), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_70), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_1), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_182), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_227), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_69), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_79), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_231), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_168), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_90), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_57), .Y(n_286) );
BUFx2_ASAP7_75t_SL g287 ( .A(n_0), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_85), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_86), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_195), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_189), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_170), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_16), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_222), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_122), .Y(n_295) );
BUFx10_ASAP7_75t_L g296 ( .A(n_113), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_112), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_11), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_106), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_262), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_82), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_98), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_266), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_80), .Y(n_304) );
INVxp33_ASAP7_75t_SL g305 ( .A(n_263), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_265), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_185), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_125), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_124), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_108), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_76), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_0), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_9), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_12), .Y(n_315) );
CKINVDCx14_ASAP7_75t_R g316 ( .A(n_251), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_121), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_257), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_142), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_8), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_179), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_72), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_232), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_171), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_138), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_111), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_186), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_136), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_169), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_39), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_87), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_104), .Y(n_332) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_117), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_123), .Y(n_334) );
NOR2xp67_ASAP7_75t_L g335 ( .A(n_198), .B(n_261), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_253), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_224), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_178), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_95), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_256), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_219), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_35), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_75), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_103), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_4), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_67), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_159), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_28), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_131), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_73), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_199), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_150), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_7), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_226), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_148), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_248), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_45), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_97), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_119), .Y(n_359) );
INVxp33_ASAP7_75t_SL g360 ( .A(n_207), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_110), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_132), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_240), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_183), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_204), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_52), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_58), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_235), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_156), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_152), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_44), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_65), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_51), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_255), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_245), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_118), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_53), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_14), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_243), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_37), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_101), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_30), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_94), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_20), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_211), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_21), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_109), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_93), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_89), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_246), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_62), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_6), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_44), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_114), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_71), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_218), .B(n_244), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_206), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_83), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_162), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_7), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_74), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_146), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_65), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_27), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g405 ( .A(n_84), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_2), .Y(n_406) );
INVxp67_ASAP7_75t_SL g407 ( .A(n_134), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_22), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_209), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_91), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_297), .B(n_1), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_275), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_291), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_378), .B(n_3), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_284), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_379), .B(n_3), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_275), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_284), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_322), .B(n_4), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_405), .Y(n_420) );
INVx5_ASAP7_75t_L g421 ( .A(n_284), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_316), .B(n_5), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_315), .Y(n_423) );
AND2x6_ASAP7_75t_L g424 ( .A(n_291), .B(n_78), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_386), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_383), .B(n_5), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_372), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_387), .B(n_6), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_284), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_353), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_323), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_384), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_409), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_323), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_384), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_393), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_316), .B(n_8), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_274), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_323), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_315), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_441) );
NOR2xp33_ASAP7_75t_R g442 ( .A(n_324), .B(n_81), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_323), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_340), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_421), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_422), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_425), .B(n_394), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_431), .B(n_305), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_415), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_425), .B(n_296), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_415), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_413), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_432), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_413), .B(n_314), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_414), .B(n_296), .Y(n_455) );
AND2x6_ASAP7_75t_L g456 ( .A(n_422), .B(n_269), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_415), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_418), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_441), .B(n_287), .Y(n_460) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_432), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_414), .B(n_296), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_420), .B(n_305), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_418), .Y(n_465) );
BUFx3_ASAP7_75t_L g466 ( .A(n_424), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_438), .A2(n_272), .B1(n_278), .B2(n_270), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_434), .B(n_360), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_419), .A2(n_400), .B1(n_314), .B2(n_392), .Y(n_469) );
AND2x6_ASAP7_75t_L g470 ( .A(n_438), .B(n_271), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_419), .B(n_273), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_412), .B(n_400), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_417), .B(n_273), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_417), .B(n_276), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_439), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_423), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_427), .B(n_360), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_427), .B(n_276), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_426), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_426), .A2(n_312), .B1(n_321), .B2(n_274), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_428), .B(n_283), .Y(n_484) );
AND2x6_ASAP7_75t_L g485 ( .A(n_428), .B(n_277), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_430), .Y(n_486) );
AND2x6_ASAP7_75t_L g487 ( .A(n_424), .B(n_410), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_442), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g489 ( .A(n_411), .B(n_386), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_466), .B(n_279), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_466), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_487), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_482), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_463), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_482), .B(n_280), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_455), .B(n_283), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_487), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_455), .B(n_290), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_463), .Y(n_499) );
AND2x6_ASAP7_75t_SL g500 ( .A(n_460), .B(n_441), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_463), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_462), .B(n_290), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_446), .Y(n_503) );
NOR2x2_ASAP7_75t_L g504 ( .A(n_460), .B(n_366), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_452), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_473), .B(n_416), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_462), .B(n_295), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_480), .B(n_295), .Y(n_508) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_487), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_485), .A2(n_424), .B1(n_433), .B2(n_429), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_447), .B(n_308), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_479), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_478), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_452), .B(n_281), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_446), .Y(n_516) );
BUFx2_ASAP7_75t_L g517 ( .A(n_456), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_487), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_485), .A2(n_424), .B1(n_433), .B2(n_429), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_476), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_457), .Y(n_521) );
AND2x4_ASAP7_75t_SL g522 ( .A(n_483), .B(n_312), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_454), .B(n_308), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_484), .B(n_436), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_448), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_457), .B(n_282), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_489), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_485), .A2(n_424), .B1(n_437), .B2(n_436), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_477), .B(n_310), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_450), .B(n_286), .Y(n_530) );
AND2x6_ASAP7_75t_L g531 ( .A(n_457), .B(n_285), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_481), .B(n_310), .Y(n_532) );
BUFx12f_ASAP7_75t_L g533 ( .A(n_460), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_489), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_475), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_489), .B(n_437), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_456), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_460), .A2(n_392), .B1(n_403), .B2(n_366), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_485), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_485), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_485), .B(n_362), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_456), .B(n_362), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_456), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_449), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_488), .B(n_370), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_456), .B(n_370), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_488), .B(n_381), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_449), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_470), .B(n_381), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_470), .A2(n_424), .B1(n_293), .B2(n_313), .Y(n_550) );
BUFx2_ASAP7_75t_L g551 ( .A(n_470), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_470), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_470), .B(n_388), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_470), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_467), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_464), .B(n_388), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_445), .B(n_288), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_451), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_451), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_458), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_445), .B(n_294), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_468), .B(n_321), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g563 ( .A(n_458), .B(n_10), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_459), .Y(n_564) );
BUFx8_ASAP7_75t_SL g565 ( .A(n_469), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_459), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_487), .B(n_326), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_487), .B(n_327), .Y(n_568) );
O2A1O1Ixp5_ASAP7_75t_L g569 ( .A1(n_472), .A2(n_374), .B(n_407), .C(n_333), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_472), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_474), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_474), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_465), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_465), .Y(n_574) );
INVx4_ASAP7_75t_L g575 ( .A(n_453), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_471), .B(n_299), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_471), .B(n_339), .Y(n_577) );
OAI22xp5_ASAP7_75t_SL g578 ( .A1(n_486), .A2(n_404), .B1(n_403), .B2(n_363), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_494), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_493), .B(n_339), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_555), .A2(n_320), .B(n_330), .C(n_298), .Y(n_581) );
BUFx2_ASAP7_75t_L g582 ( .A(n_493), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_L g583 ( .A1(n_495), .A2(n_345), .B(n_346), .C(n_342), .Y(n_583) );
BUFx3_ASAP7_75t_L g584 ( .A(n_513), .Y(n_584) );
O2A1O1Ixp33_ASAP7_75t_L g585 ( .A1(n_495), .A2(n_357), .B(n_367), .C(n_348), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_535), .B(n_363), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_520), .B(n_371), .Y(n_587) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_491), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_503), .Y(n_589) );
BUFx3_ASAP7_75t_L g590 ( .A(n_533), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_525), .B(n_369), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_496), .B(n_369), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_498), .A2(n_377), .B(n_380), .C(n_373), .Y(n_593) );
AND2x2_ASAP7_75t_SL g594 ( .A(n_522), .B(n_401), .Y(n_594) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_491), .Y(n_595) );
INVx3_ASAP7_75t_SL g596 ( .A(n_504), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_512), .B(n_382), .Y(n_597) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_491), .Y(n_598) );
BUFx2_ASAP7_75t_R g599 ( .A(n_565), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_578), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_494), .Y(n_601) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_577), .Y(n_602) );
AND2x6_ASAP7_75t_L g603 ( .A(n_537), .B(n_300), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_515), .B(n_401), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_577), .A2(n_404), .B1(n_406), .B2(n_391), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_505), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_502), .B(n_408), .Y(n_607) );
AOI221x1_ASAP7_75t_L g608 ( .A1(n_543), .A2(n_352), .B1(n_302), .B2(n_303), .C(n_304), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_517), .B(n_395), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_499), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_538), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_507), .A2(n_393), .B(n_307), .C(n_309), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_501), .A2(n_486), .B(n_311), .Y(n_613) );
NOR2x1_ASAP7_75t_SL g614 ( .A(n_492), .B(n_306), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_529), .A2(n_318), .B(n_317), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_544), .Y(n_616) );
OR2x6_ASAP7_75t_L g617 ( .A(n_562), .B(n_335), .Y(n_617) );
BUFx12f_ASAP7_75t_L g618 ( .A(n_500), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_532), .A2(n_523), .B(n_490), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_516), .B(n_319), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g621 ( .A1(n_511), .A2(n_329), .B(n_331), .C(n_325), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_506), .B(n_398), .Y(n_622) );
OAI22xp5_ASAP7_75t_SL g623 ( .A1(n_562), .A2(n_336), .B1(n_337), .B2(n_332), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_505), .Y(n_624) );
BUFx2_ASAP7_75t_L g625 ( .A(n_531), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_522), .B(n_12), .Y(n_626) );
INVx2_ASAP7_75t_SL g627 ( .A(n_527), .Y(n_627) );
OR2x6_ASAP7_75t_L g628 ( .A(n_534), .B(n_338), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g629 ( .A1(n_536), .A2(n_343), .B(n_344), .C(n_341), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_544), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_531), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_506), .A2(n_351), .B1(n_375), .B2(n_399), .C1(n_397), .C2(n_390), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_545), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_524), .B(n_402), .Y(n_634) );
INVx4_ASAP7_75t_L g635 ( .A(n_537), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_536), .A2(n_424), .B1(n_349), .B2(n_350), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_490), .A2(n_355), .B(n_347), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_524), .B(n_358), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_556), .B(n_359), .Y(n_639) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_491), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_548), .Y(n_641) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_492), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_574), .A2(n_364), .B(n_361), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_559), .A2(n_376), .B(n_368), .C(n_385), .Y(n_644) );
NOR2x1_ASAP7_75t_SL g645 ( .A(n_492), .B(n_389), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_530), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_566), .A2(n_365), .B(n_292), .C(n_301), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_558), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_551), .A2(n_289), .B1(n_292), .B2(n_301), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_558), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_514), .A2(n_328), .B(n_289), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_508), .B(n_328), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_531), .B(n_334), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_531), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_560), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_554), .B(n_334), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_514), .A2(n_365), .B(n_356), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_526), .A2(n_356), .B(n_435), .C(n_440), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_526), .A2(n_396), .B(n_421), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g660 ( .A1(n_576), .A2(n_435), .B(n_440), .C(n_443), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_564), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_554), .A2(n_435), .B1(n_443), .B2(n_440), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_573), .A2(n_444), .B(n_443), .C(n_340), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_541), .A2(n_421), .B(n_444), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_531), .B(n_13), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_530), .B(n_14), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_576), .A2(n_444), .B(n_16), .C(n_17), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_545), .B(n_15), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_542), .Y(n_669) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_492), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_521), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_571), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_552), .A2(n_354), .B1(n_340), .B2(n_432), .Y(n_673) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_497), .Y(n_674) );
AO22x1_ASAP7_75t_L g675 ( .A1(n_547), .A2(n_340), .B1(n_354), .B2(n_18), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_539), .B(n_15), .Y(n_676) );
BUFx12f_ASAP7_75t_L g677 ( .A(n_540), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_571), .B(n_17), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_546), .B(n_20), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_550), .A2(n_432), .B1(n_22), .B2(n_23), .Y(n_680) );
INVxp67_ASAP7_75t_SL g681 ( .A(n_497), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_549), .B(n_21), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_553), .A2(n_453), .B1(n_461), .B2(n_25), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_497), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_572), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_572), .Y(n_686) );
INVxp67_ASAP7_75t_L g687 ( .A(n_557), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_567), .B(n_23), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_570), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_510), .A2(n_461), .B(n_453), .C(n_26), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_510), .A2(n_461), .B(n_453), .C(n_26), .Y(n_691) );
INVx5_ASAP7_75t_L g692 ( .A(n_509), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_568), .A2(n_461), .B(n_453), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_557), .Y(n_694) );
INVx3_ASAP7_75t_L g695 ( .A(n_509), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_575), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_561), .B(n_24), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_575), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_561), .A2(n_461), .B1(n_25), .B2(n_27), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_563), .A2(n_24), .B(n_28), .C(n_29), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_509), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_701) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_509), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_586), .A2(n_528), .B1(n_519), .B2(n_518), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_616), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_616), .B(n_519), .Y(n_705) );
OAI21x1_ASAP7_75t_L g706 ( .A1(n_693), .A2(n_528), .B(n_518), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_630), .A2(n_518), .B1(n_32), .B2(n_33), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_582), .Y(n_708) );
OAI21xp5_ASAP7_75t_L g709 ( .A1(n_619), .A2(n_518), .B(n_31), .Y(n_709) );
BUFx3_ASAP7_75t_L g710 ( .A(n_584), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_589), .Y(n_711) );
OAI21xp33_ASAP7_75t_SL g712 ( .A1(n_630), .A2(n_32), .B(n_33), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_648), .B(n_34), .Y(n_713) );
INVx3_ASAP7_75t_L g714 ( .A(n_635), .Y(n_714) );
OAI21x1_ASAP7_75t_L g715 ( .A1(n_664), .A2(n_92), .B(n_88), .Y(n_715) );
INVx3_ASAP7_75t_L g716 ( .A(n_635), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_648), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_612), .A2(n_34), .B(n_35), .C(n_36), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_650), .B(n_36), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_661), .B(n_37), .Y(n_720) );
NAND2x1_ASAP7_75t_L g721 ( .A(n_661), .B(n_96), .Y(n_721) );
OAI21x1_ASAP7_75t_L g722 ( .A1(n_610), .A2(n_100), .B(n_99), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_672), .B(n_38), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_641), .Y(n_724) );
O2A1O1Ixp33_ASAP7_75t_SL g725 ( .A1(n_690), .A2(n_691), .B(n_647), .C(n_629), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_678), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_628), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_610), .A2(n_40), .B(n_42), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_581), .A2(n_42), .B1(n_43), .B2(n_45), .C(n_46), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_596), .Y(n_730) );
NAND2x1p5_ASAP7_75t_L g731 ( .A(n_692), .B(n_43), .Y(n_731) );
AO31x2_ASAP7_75t_L g732 ( .A1(n_608), .A2(n_46), .A3(n_47), .B(n_48), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_655), .A2(n_47), .B(n_48), .Y(n_733) );
OAI21x1_ASAP7_75t_L g734 ( .A1(n_659), .A2(n_176), .B(n_267), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_587), .Y(n_735) );
OAI21x1_ASAP7_75t_L g736 ( .A1(n_613), .A2(n_175), .B(n_264), .Y(n_736) );
BUFx4f_ASAP7_75t_L g737 ( .A(n_594), .Y(n_737) );
NOR2xp67_ASAP7_75t_L g738 ( .A(n_586), .B(n_49), .Y(n_738) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_628), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_602), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_740) );
INVx2_ASAP7_75t_SL g741 ( .A(n_590), .Y(n_741) );
AO21x2_ASAP7_75t_L g742 ( .A1(n_683), .A2(n_177), .B(n_260), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_621), .A2(n_50), .B(n_52), .C(n_53), .Y(n_743) );
CKINVDCx14_ASAP7_75t_R g744 ( .A(n_580), .Y(n_744) );
AOI21x1_ASAP7_75t_L g745 ( .A1(n_675), .A2(n_181), .B(n_259), .Y(n_745) );
AO31x2_ASAP7_75t_L g746 ( .A1(n_644), .A2(n_54), .A3(n_55), .B(n_56), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_580), .B(n_54), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_591), .B(n_605), .Y(n_748) );
OA21x2_ASAP7_75t_L g749 ( .A1(n_663), .A2(n_180), .B(n_258), .Y(n_749) );
OR2x6_ASAP7_75t_L g750 ( .A(n_625), .B(n_55), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_592), .B(n_56), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_646), .B(n_57), .Y(n_752) );
OR2x6_ASAP7_75t_L g753 ( .A(n_626), .B(n_59), .Y(n_753) );
NOR2xp67_ASAP7_75t_L g754 ( .A(n_618), .B(n_59), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_620), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_643), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_756) );
AO21x2_ASAP7_75t_L g757 ( .A1(n_653), .A2(n_184), .B(n_254), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_607), .B(n_60), .Y(n_758) );
AO31x2_ASAP7_75t_L g759 ( .A1(n_614), .A2(n_61), .A3(n_63), .B(n_64), .Y(n_759) );
NAND2x1p5_ASAP7_75t_L g760 ( .A(n_692), .B(n_63), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_676), .Y(n_761) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_615), .A2(n_64), .B(n_66), .Y(n_762) );
INVx3_ASAP7_75t_L g763 ( .A(n_677), .Y(n_763) );
OA21x2_ASAP7_75t_L g764 ( .A1(n_651), .A2(n_190), .B(n_250), .Y(n_764) );
AO21x2_ASAP7_75t_L g765 ( .A1(n_679), .A2(n_188), .B(n_249), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_652), .A2(n_174), .B(n_247), .Y(n_766) );
OR2x6_ASAP7_75t_L g767 ( .A(n_604), .B(n_66), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_597), .B(n_67), .Y(n_768) );
BUFx12f_ASAP7_75t_L g769 ( .A(n_617), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_620), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_666), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_632), .A2(n_68), .B1(n_102), .B2(n_105), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_657), .A2(n_192), .B(n_107), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_697), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_676), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_583), .Y(n_776) );
OA21x2_ASAP7_75t_L g777 ( .A1(n_636), .A2(n_193), .B(n_115), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_638), .B(n_68), .Y(n_778) );
INVx1_ASAP7_75t_SL g779 ( .A(n_631), .Y(n_779) );
BUFx3_ASAP7_75t_L g780 ( .A(n_600), .Y(n_780) );
OA21x2_ASAP7_75t_L g781 ( .A1(n_665), .A2(n_116), .B(n_126), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_686), .A2(n_127), .B(n_128), .Y(n_782) );
OA21x2_ASAP7_75t_L g783 ( .A1(n_673), .A2(n_129), .B(n_130), .Y(n_783) );
OAI21x1_ASAP7_75t_SL g784 ( .A1(n_645), .A2(n_133), .B(n_135), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_639), .A2(n_137), .B(n_139), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_623), .A2(n_140), .B1(n_141), .B2(n_143), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_611), .B(n_144), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_585), .Y(n_788) );
OA21x2_ASAP7_75t_L g789 ( .A1(n_688), .A2(n_145), .B(n_147), .Y(n_789) );
AND2x4_ASAP7_75t_L g790 ( .A(n_627), .B(n_268), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_692), .Y(n_791) );
OAI21x1_ASAP7_75t_L g792 ( .A1(n_658), .A2(n_149), .B(n_151), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_593), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_633), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_794) );
BUFx2_ASAP7_75t_L g795 ( .A(n_603), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_637), .A2(n_157), .B(n_158), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_694), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_654), .B(n_242), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_700), .Y(n_799) );
AO21x2_ASAP7_75t_L g800 ( .A1(n_668), .A2(n_160), .B(n_163), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_682), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_622), .B(n_164), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_669), .B(n_165), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_634), .A2(n_166), .B(n_167), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_671), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_696), .Y(n_806) );
OAI21x1_ASAP7_75t_L g807 ( .A1(n_660), .A2(n_172), .B(n_173), .Y(n_807) );
OAI211xp5_ASAP7_75t_L g808 ( .A1(n_649), .A2(n_191), .B(n_194), .C(n_196), .Y(n_808) );
A2O1A1Ixp33_ASAP7_75t_L g809 ( .A1(n_667), .A2(n_197), .B(n_200), .C(n_201), .Y(n_809) );
OAI21x1_ASAP7_75t_L g810 ( .A1(n_656), .A2(n_662), .B(n_606), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_603), .A2(n_202), .B1(n_203), .B2(n_205), .Y(n_811) );
O2A1O1Ixp33_ASAP7_75t_SL g812 ( .A1(n_701), .A2(n_208), .B(n_210), .C(n_212), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_687), .B(n_213), .Y(n_813) );
AND2x4_ASAP7_75t_L g814 ( .A(n_689), .B(n_624), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_603), .A2(n_214), .B1(n_215), .B2(n_216), .Y(n_815) );
AND2x4_ASAP7_75t_L g816 ( .A(n_606), .B(n_217), .Y(n_816) );
OAI21x1_ASAP7_75t_L g817 ( .A1(n_624), .A2(n_220), .B(n_221), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_699), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_579), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_601), .B(n_225), .Y(n_820) );
OAI21x1_ASAP7_75t_L g821 ( .A1(n_695), .A2(n_228), .B(n_229), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_599), .Y(n_822) );
AO21x2_ASAP7_75t_L g823 ( .A1(n_680), .A2(n_230), .B(n_233), .Y(n_823) );
AO31x2_ASAP7_75t_L g824 ( .A1(n_685), .A2(n_234), .A3(n_236), .B(n_237), .Y(n_824) );
BUFx2_ASAP7_75t_L g825 ( .A(n_603), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_588), .A2(n_238), .B1(n_239), .B2(n_241), .Y(n_826) );
AND2x4_ASAP7_75t_L g827 ( .A(n_609), .B(n_698), .Y(n_827) );
INVx3_ASAP7_75t_L g828 ( .A(n_642), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_681), .B(n_588), .Y(n_829) );
INVx1_ASAP7_75t_SL g830 ( .A(n_588), .Y(n_830) );
AND2x4_ASAP7_75t_L g831 ( .A(n_642), .B(n_674), .Y(n_831) );
OA21x2_ASAP7_75t_L g832 ( .A1(n_595), .A2(n_598), .B(n_640), .Y(n_832) );
INVx3_ASAP7_75t_L g833 ( .A(n_670), .Y(n_833) );
OA21x2_ASAP7_75t_L g834 ( .A1(n_706), .A2(n_595), .B(n_598), .Y(n_834) );
OAI221xp5_ASAP7_75t_L g835 ( .A1(n_748), .A2(n_640), .B1(n_670), .B2(n_674), .C(n_684), .Y(n_835) );
OAI221xp5_ASAP7_75t_L g836 ( .A1(n_737), .A2(n_640), .B1(n_670), .B2(n_684), .C(n_702), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_704), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_739), .A2(n_702), .B1(n_797), .B2(n_744), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_750), .A2(n_775), .B1(n_761), .B2(n_739), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_767), .A2(n_793), .B1(n_799), .B2(n_747), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_767), .A2(n_753), .B1(n_750), .B2(n_769), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_725), .A2(n_778), .B(n_709), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_795), .B(n_825), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_727), .A2(n_756), .B1(n_729), .B2(n_726), .C(n_801), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g845 ( .A1(n_750), .A2(n_767), .B1(n_753), .B2(n_768), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_753), .A2(n_751), .B1(n_776), .B2(n_788), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_708), .B(n_752), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_771), .A2(n_738), .B1(n_761), .B2(n_770), .Y(n_848) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_717), .Y(n_849) );
AOI21xp33_ASAP7_75t_L g850 ( .A1(n_802), .A2(n_818), .B(n_778), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_724), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_711), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_723), .Y(n_853) );
O2A1O1Ixp33_ASAP7_75t_L g854 ( .A1(n_743), .A2(n_718), .B(n_756), .C(n_727), .Y(n_854) );
INVxp67_ASAP7_75t_L g855 ( .A(n_752), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g856 ( .A1(n_755), .A2(n_772), .B1(n_758), .B2(n_729), .C(n_762), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_775), .A2(n_707), .B1(n_728), .B2(n_760), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_774), .A2(n_772), .B1(n_780), .B2(n_758), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_805), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_703), .A2(n_719), .B1(n_720), .B2(n_713), .Y(n_860) );
INVx1_ASAP7_75t_SL g861 ( .A(n_710), .Y(n_861) );
OAI222xp33_ASAP7_75t_L g862 ( .A1(n_707), .A2(n_731), .B1(n_760), .B2(n_713), .C1(n_720), .C2(n_719), .Y(n_862) );
AND2x4_ASAP7_75t_L g863 ( .A(n_790), .B(n_814), .Y(n_863) );
NAND2x1p5_ASAP7_75t_L g864 ( .A(n_714), .B(n_716), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_723), .A2(n_790), .B1(n_827), .B2(n_762), .Y(n_865) );
A2O1A1Ixp33_ASAP7_75t_L g866 ( .A1(n_712), .A2(n_728), .B(n_733), .C(n_785), .Y(n_866) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_822), .Y(n_867) );
O2A1O1Ixp33_ASAP7_75t_L g868 ( .A1(n_733), .A2(n_809), .B(n_705), .C(n_740), .Y(n_868) );
AOI221xp5_ASAP7_75t_L g869 ( .A1(n_730), .A2(n_786), .B1(n_787), .B2(n_741), .C(n_705), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_746), .Y(n_870) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_786), .A2(n_763), .B1(n_812), .B2(n_785), .C(n_819), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_746), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_806), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_814), .B(n_754), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_763), .B(n_791), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_731), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_732), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_827), .B(n_791), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_820), .A2(n_813), .B(n_766), .Y(n_879) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_830), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_803), .A2(n_816), .B1(n_779), .B2(n_815), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_816), .A2(n_779), .B1(n_815), .B2(n_811), .Y(n_882) );
INVx6_ASAP7_75t_SL g883 ( .A(n_798), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_732), .Y(n_884) );
BUFx12f_ASAP7_75t_L g885 ( .A(n_798), .Y(n_885) );
NOR2x1p5_ASAP7_75t_L g886 ( .A(n_714), .B(n_716), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_813), .A2(n_823), .B1(n_800), .B2(n_742), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_820), .A2(n_804), .B(n_832), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_732), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_823), .A2(n_829), .B1(n_796), .B2(n_777), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_830), .B(n_833), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_759), .Y(n_892) );
AOI21x1_ASAP7_75t_L g893 ( .A1(n_832), .A2(n_745), .B(n_789), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_828), .B(n_833), .Y(n_894) );
OR2x2_ASAP7_75t_L g895 ( .A(n_759), .B(n_828), .Y(n_895) );
OAI211xp5_ASAP7_75t_L g896 ( .A1(n_811), .A2(n_826), .B(n_794), .C(n_808), .Y(n_896) );
INVx3_ASAP7_75t_L g897 ( .A(n_831), .Y(n_897) );
CKINVDCx6p67_ASAP7_75t_R g898 ( .A(n_831), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_759), .B(n_826), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_824), .B(n_796), .Y(n_900) );
AOI222xp33_ASAP7_75t_L g901 ( .A1(n_808), .A2(n_784), .B1(n_722), .B2(n_736), .C1(n_810), .C2(n_817), .Y(n_901) );
AND2x4_ASAP7_75t_L g902 ( .A(n_734), .B(n_821), .Y(n_902) );
AO221x2_ASAP7_75t_L g903 ( .A1(n_824), .A2(n_789), .B1(n_777), .B2(n_781), .C(n_765), .Y(n_903) );
AOI221xp5_ASAP7_75t_L g904 ( .A1(n_721), .A2(n_757), .B1(n_765), .B2(n_824), .C(n_749), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_757), .A2(n_783), .B1(n_781), .B2(n_764), .Y(n_905) );
OAI22xp33_ASAP7_75t_L g906 ( .A1(n_783), .A2(n_764), .B1(n_749), .B2(n_782), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_715), .A2(n_792), .B1(n_773), .B2(n_807), .Y(n_907) );
OAI221xp5_ASAP7_75t_SL g908 ( .A1(n_748), .A2(n_460), .B1(n_605), .B2(n_483), .C(n_744), .Y(n_908) );
OAI22xp5_ASAP7_75t_SL g909 ( .A1(n_744), .A2(n_594), .B1(n_423), .B2(n_538), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_737), .A2(n_594), .B1(n_748), .B2(n_522), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_704), .Y(n_911) );
A2O1A1Ixp33_ASAP7_75t_L g912 ( .A1(n_799), .A2(n_793), .B(n_735), .C(n_712), .Y(n_912) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_704), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_735), .B(n_493), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_711), .Y(n_915) );
OAI221xp5_ASAP7_75t_L g916 ( .A1(n_748), .A2(n_737), .B1(n_617), .B2(n_623), .C(n_483), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_735), .B(n_493), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_750), .A2(n_775), .B1(n_577), .B2(n_594), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g919 ( .A1(n_735), .A2(n_605), .B1(n_555), .B2(n_581), .C(n_469), .Y(n_919) );
AOI221xp5_ASAP7_75t_SL g920 ( .A1(n_799), .A2(n_605), .B1(n_623), .B2(n_581), .C(n_593), .Y(n_920) );
OAI21xp5_ASAP7_75t_L g921 ( .A1(n_735), .A2(n_569), .B(n_629), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_725), .A2(n_693), .B(n_778), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_711), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_737), .A2(n_594), .B1(n_748), .B2(n_522), .Y(n_924) );
CKINVDCx11_ASAP7_75t_R g925 ( .A(n_710), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_737), .A2(n_594), .B1(n_748), .B2(n_522), .Y(n_926) );
BUFx2_ASAP7_75t_L g927 ( .A(n_739), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_711), .Y(n_928) );
OAI221xp5_ASAP7_75t_L g929 ( .A1(n_748), .A2(n_737), .B1(n_617), .B2(n_623), .C(n_483), .Y(n_929) );
AOI221xp5_ASAP7_75t_L g930 ( .A1(n_735), .A2(n_605), .B1(n_555), .B2(n_581), .C(n_469), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_737), .A2(n_594), .B1(n_748), .B2(n_522), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_711), .Y(n_932) );
OAI221xp5_ASAP7_75t_SL g933 ( .A1(n_748), .A2(n_460), .B1(n_605), .B2(n_483), .C(n_744), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_711), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_735), .B(n_493), .Y(n_935) );
INVx3_ASAP7_75t_L g936 ( .A(n_714), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g937 ( .A1(n_737), .A2(n_594), .B1(n_578), .B2(n_586), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_711), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_750), .A2(n_775), .B1(n_577), .B2(n_594), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_750), .A2(n_775), .B1(n_577), .B2(n_594), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_711), .Y(n_941) );
AOI21xp33_ASAP7_75t_L g942 ( .A1(n_799), .A2(n_748), .B(n_612), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_739), .B(n_493), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_711), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g945 ( .A(n_748), .B(n_479), .Y(n_945) );
AND2x4_ASAP7_75t_L g946 ( .A(n_735), .B(n_739), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_704), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_737), .A2(n_594), .B1(n_748), .B2(n_522), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_737), .A2(n_594), .B1(n_748), .B2(n_522), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_735), .B(n_493), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_711), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_870), .Y(n_952) );
BUFx2_ASAP7_75t_L g953 ( .A(n_883), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_834), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_849), .B(n_913), .Y(n_955) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_943), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_849), .B(n_913), .Y(n_957) );
A2O1A1Ixp33_ASAP7_75t_L g958 ( .A1(n_854), .A2(n_844), .B(n_869), .C(n_850), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_872), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_877), .Y(n_960) );
BUFx3_ASAP7_75t_L g961 ( .A(n_898), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_884), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_834), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_837), .B(n_911), .Y(n_964) );
BUFx2_ASAP7_75t_L g965 ( .A(n_883), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_947), .B(n_851), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_889), .Y(n_967) );
INVx2_ASAP7_75t_L g968 ( .A(n_893), .Y(n_968) );
BUFx2_ASAP7_75t_L g969 ( .A(n_880), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_916), .A2(n_929), .B1(n_845), .B2(n_844), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_892), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_852), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_859), .B(n_853), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_915), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_923), .B(n_928), .Y(n_975) );
AOI221xp5_ASAP7_75t_L g976 ( .A1(n_908), .A2(n_933), .B1(n_945), .B2(n_942), .C(n_930), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_932), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_934), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_938), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_908), .B(n_933), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_941), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_919), .B(n_930), .Y(n_982) );
AND2x4_ASAP7_75t_L g983 ( .A(n_876), .B(n_897), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_944), .B(n_951), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_873), .B(n_912), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_895), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_946), .B(n_863), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_918), .A2(n_939), .B1(n_940), .B2(n_926), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_880), .Y(n_989) );
INVxp67_ASAP7_75t_SL g990 ( .A(n_855), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_946), .B(n_863), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_865), .B(n_855), .Y(n_992) );
INVx5_ASAP7_75t_L g993 ( .A(n_885), .Y(n_993) );
INVx1_ASAP7_75t_SL g994 ( .A(n_927), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_858), .B(n_846), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_891), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_866), .B(n_842), .Y(n_997) );
OAI211xp5_ASAP7_75t_L g998 ( .A1(n_841), .A2(n_931), .B(n_949), .C(n_924), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_840), .B(n_897), .Y(n_999) );
INVxp67_ASAP7_75t_SL g1000 ( .A(n_857), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_894), .Y(n_1001) );
INVx8_ASAP7_75t_L g1002 ( .A(n_843), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_860), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_914), .B(n_950), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_899), .Y(n_1005) );
BUFx3_ASAP7_75t_L g1006 ( .A(n_864), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_917), .B(n_935), .Y(n_1007) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_864), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_842), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_902), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_919), .B(n_920), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_902), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_886), .B(n_847), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_936), .B(n_921), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_875), .Y(n_1015) );
OR2x2_ASAP7_75t_L g1016 ( .A(n_878), .B(n_839), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_922), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_848), .B(n_869), .Y(n_1018) );
AND2x4_ASAP7_75t_SL g1019 ( .A(n_838), .B(n_874), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_910), .B(n_948), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_854), .B(n_900), .Y(n_1021) );
INVx2_ASAP7_75t_R g1022 ( .A(n_903), .Y(n_1022) );
AND2x4_ASAP7_75t_SL g1023 ( .A(n_937), .B(n_890), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_861), .B(n_909), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_882), .B(n_871), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_925), .B(n_856), .Y(n_1026) );
INVx2_ASAP7_75t_SL g1027 ( .A(n_881), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_836), .Y(n_1028) );
BUFx3_ASAP7_75t_L g1029 ( .A(n_835), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_906), .Y(n_1030) );
INVx2_ASAP7_75t_L g1031 ( .A(n_905), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_868), .B(n_871), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_868), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_887), .B(n_901), .Y(n_1034) );
BUFx2_ASAP7_75t_L g1035 ( .A(n_904), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1005), .B(n_888), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_980), .A2(n_896), .B1(n_862), .B2(n_907), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1005), .B(n_904), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1021), .B(n_879), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_1021), .B(n_896), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1041 ( .A(n_989), .B(n_867), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_955), .B(n_862), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_955), .B(n_957), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_957), .B(n_1025), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1025), .B(n_986), .Y(n_1045) );
INVxp67_ASAP7_75t_SL g1046 ( .A(n_969), .Y(n_1046) );
OAI21xp33_ASAP7_75t_SL g1047 ( .A1(n_1027), .A2(n_976), .B(n_985), .Y(n_1047) );
AOI21xp5_ASAP7_75t_L g1048 ( .A1(n_954), .A2(n_963), .B(n_968), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_952), .Y(n_1049) );
BUFx3_ASAP7_75t_L g1050 ( .A(n_1002), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_989), .B(n_969), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_952), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_959), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_958), .B(n_1003), .Y(n_1054) );
BUFx3_ASAP7_75t_L g1055 ( .A(n_1002), .Y(n_1055) );
OAI211xp5_ASAP7_75t_L g1056 ( .A1(n_970), .A2(n_998), .B(n_988), .C(n_1026), .Y(n_1056) );
NAND2x1_ASAP7_75t_L g1057 ( .A(n_1010), .B(n_1012), .Y(n_1057) );
AND2x4_ASAP7_75t_L g1058 ( .A(n_1010), .B(n_1012), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1003), .B(n_975), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_975), .B(n_984), .Y(n_1060) );
INVx1_ASAP7_75t_SL g1061 ( .A(n_994), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1033), .B(n_982), .Y(n_1062) );
OR2x2_ASAP7_75t_SL g1063 ( .A(n_1016), .B(n_1012), .Y(n_1063) );
OAI31xp33_ASAP7_75t_SL g1064 ( .A1(n_1018), .A2(n_995), .A3(n_1000), .B(n_994), .Y(n_1064) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_1029), .Y(n_1065) );
NOR2x1_ASAP7_75t_SL g1066 ( .A(n_1006), .B(n_1029), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_984), .B(n_1033), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1068 ( .A(n_971), .B(n_960), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_962), .B(n_967), .Y(n_1069) );
BUFx3_ASAP7_75t_L g1070 ( .A(n_1002), .Y(n_1070) );
INVx5_ASAP7_75t_SL g1071 ( .A(n_983), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_962), .B(n_967), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_954), .A2(n_963), .B(n_968), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1014), .B(n_971), .Y(n_1074) );
INVxp67_ASAP7_75t_L g1075 ( .A(n_985), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_972), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_1014), .B(n_1034), .Y(n_1077) );
INVx2_ASAP7_75t_SL g1078 ( .A(n_1002), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_972), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1034), .B(n_964), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_974), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_964), .B(n_977), .Y(n_1082) );
BUFx3_ASAP7_75t_L g1083 ( .A(n_1002), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_974), .B(n_979), .Y(n_1084) );
BUFx2_ASAP7_75t_L g1085 ( .A(n_1008), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1011), .B(n_996), .Y(n_1086) );
AOI221xp5_ASAP7_75t_L g1087 ( .A1(n_1007), .A2(n_1018), .B1(n_1020), .B2(n_995), .C(n_1032), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_977), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_978), .B(n_979), .Y(n_1089) );
INVx2_ASAP7_75t_SL g1090 ( .A(n_1006), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g1091 ( .A(n_1015), .Y(n_1091) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_1004), .A2(n_993), .B1(n_961), .B2(n_1024), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_954), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_996), .B(n_978), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g1095 ( .A1(n_1047), .A2(n_956), .B1(n_981), .B2(n_990), .C(n_992), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1049), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_1060), .B(n_981), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1049), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1052), .Y(n_1099) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1093), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1074), .B(n_1035), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1052), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1053), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1074), .B(n_1035), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1053), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1039), .B(n_1045), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1039), .B(n_1031), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_1068), .B(n_963), .Y(n_1108) );
NAND2xp5_ASAP7_75t_SL g1109 ( .A(n_1064), .B(n_993), .Y(n_1109) );
AND2x2_ASAP7_75t_SL g1110 ( .A(n_1064), .B(n_1023), .Y(n_1110) );
OAI33xp33_ASAP7_75t_L g1111 ( .A1(n_1037), .A2(n_1016), .A3(n_1004), .B1(n_1001), .B2(n_997), .B3(n_1017), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1112 ( .A(n_1043), .B(n_1031), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1059), .B(n_1022), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1080), .B(n_973), .Y(n_1114) );
INVx3_ASAP7_75t_L g1115 ( .A(n_1057), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1080), .B(n_973), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1059), .B(n_1022), .Y(n_1117) );
BUFx3_ASAP7_75t_L g1118 ( .A(n_1085), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1038), .B(n_1022), .Y(n_1119) );
INVx4_ASAP7_75t_L g1120 ( .A(n_1050), .Y(n_1120) );
OAI221xp5_ASAP7_75t_L g1121 ( .A1(n_1056), .A2(n_1047), .B1(n_1087), .B2(n_1054), .C(n_1062), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1038), .B(n_1077), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1082), .B(n_999), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1077), .B(n_1030), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1043), .B(n_999), .Y(n_1125) );
NOR3xp33_ASAP7_75t_SL g1126 ( .A(n_1056), .B(n_1001), .C(n_993), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1069), .B(n_1072), .Y(n_1127) );
INVx1_ASAP7_75t_SL g1128 ( .A(n_1061), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_1051), .B(n_997), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_1091), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1044), .B(n_966), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1044), .B(n_966), .Y(n_1132) );
AND2x4_ASAP7_75t_SL g1133 ( .A(n_1078), .B(n_987), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1036), .B(n_1009), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_1040), .A2(n_1023), .B1(n_1019), .B2(n_1028), .Y(n_1135) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_1054), .A2(n_953), .B1(n_965), .B2(n_961), .C(n_1013), .Y(n_1136) );
HB1xp67_ASAP7_75t_L g1137 ( .A(n_1061), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1127), .B(n_1036), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1127), .B(n_1042), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1122), .B(n_1067), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1130), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1096), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1106), .B(n_1068), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1122), .B(n_1067), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1145 ( .A(n_1113), .B(n_1058), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_1106), .B(n_1068), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1101), .B(n_1084), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1148 ( .A(n_1121), .B(n_1041), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1096), .Y(n_1149) );
INVx1_ASAP7_75t_SL g1150 ( .A(n_1133), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1119), .B(n_1042), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1104), .B(n_1084), .Y(n_1152) );
OR2x2_ASAP7_75t_L g1153 ( .A(n_1125), .B(n_1063), .Y(n_1153) );
INVxp67_ASAP7_75t_L g1154 ( .A(n_1137), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1098), .Y(n_1155) );
OR2x2_ASAP7_75t_L g1156 ( .A(n_1097), .B(n_1046), .Y(n_1156) );
NOR2xp33_ASAP7_75t_L g1157 ( .A(n_1136), .B(n_1041), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1099), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1104), .B(n_1089), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1128), .B(n_1089), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1161 ( .A(n_1113), .B(n_1058), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1123), .B(n_1075), .Y(n_1162) );
NAND4xp25_ASAP7_75t_L g1163 ( .A(n_1095), .B(n_1062), .C(n_1065), .D(n_1086), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1119), .B(n_1058), .Y(n_1164) );
INVx2_ASAP7_75t_SL g1165 ( .A(n_1118), .Y(n_1165) );
NAND2xp33_ASAP7_75t_SL g1166 ( .A(n_1109), .B(n_1085), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1099), .Y(n_1167) );
NOR2xp33_ASAP7_75t_L g1168 ( .A(n_1114), .B(n_1092), .Y(n_1168) );
AOI21xp5_ASAP7_75t_L g1169 ( .A1(n_1111), .A2(n_1066), .B(n_1048), .Y(n_1169) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1100), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1102), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1117), .B(n_1058), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1102), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1103), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1103), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1105), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1141), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1138), .B(n_1117), .Y(n_1178) );
INVx1_ASAP7_75t_SL g1179 ( .A(n_1150), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1139), .B(n_1124), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1138), .B(n_1124), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1142), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1149), .Y(n_1183) );
NAND4xp25_ASAP7_75t_L g1184 ( .A(n_1148), .B(n_1135), .C(n_1086), .D(n_1116), .Y(n_1184) );
NOR2xp33_ASAP7_75t_L g1185 ( .A(n_1148), .B(n_1157), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g1186 ( .A1(n_1157), .A2(n_1110), .B1(n_1126), .B2(n_1120), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1155), .Y(n_1187) );
OAI31xp33_ASAP7_75t_L g1188 ( .A1(n_1166), .A2(n_1133), .A3(n_1019), .B(n_1070), .Y(n_1188) );
NOR3xp33_ASAP7_75t_L g1189 ( .A(n_1163), .B(n_953), .C(n_965), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1140), .B(n_1134), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1158), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1167), .Y(n_1192) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1144), .B(n_1112), .Y(n_1193) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_1154), .B(n_1131), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1170), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1170), .Y(n_1196) );
AOI21xp33_ASAP7_75t_SL g1197 ( .A1(n_1165), .A2(n_1090), .B(n_1129), .Y(n_1197) );
AND2x4_ASAP7_75t_L g1198 ( .A(n_1145), .B(n_1108), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1171), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1147), .B(n_1112), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1173), .Y(n_1201) );
AOI22xp33_ASAP7_75t_SL g1202 ( .A1(n_1185), .A2(n_1120), .B1(n_1168), .B2(n_1066), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1182), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1204 ( .A(n_1185), .B(n_1151), .Y(n_1204) );
XNOR2xp5_ASAP7_75t_L g1205 ( .A(n_1179), .B(n_1186), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1178), .B(n_1143), .Y(n_1206) );
INVx3_ASAP7_75t_L g1207 ( .A(n_1198), .Y(n_1207) );
INVxp67_ASAP7_75t_SL g1208 ( .A(n_1195), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1183), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1196), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1177), .B(n_1151), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1181), .B(n_1143), .Y(n_1212) );
O2A1O1Ixp33_ASAP7_75t_L g1213 ( .A1(n_1189), .A2(n_1169), .B(n_1153), .C(n_1094), .Y(n_1213) );
INVx2_ASAP7_75t_SL g1214 ( .A(n_1198), .Y(n_1214) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1187), .Y(n_1215) );
OAI21xp33_ASAP7_75t_L g1216 ( .A1(n_1189), .A2(n_1146), .B(n_1160), .Y(n_1216) );
XOR2x2_ASAP7_75t_L g1217 ( .A(n_1194), .B(n_1050), .Y(n_1217) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_1202), .A2(n_1197), .B1(n_1193), .B2(n_1190), .Y(n_1218) );
AOI222xp33_ASAP7_75t_L g1219 ( .A1(n_1216), .A2(n_1194), .B1(n_1199), .B2(n_1192), .C1(n_1191), .C2(n_1201), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1203), .Y(n_1220) );
OA21x2_ASAP7_75t_L g1221 ( .A1(n_1205), .A2(n_1196), .B(n_1073), .Y(n_1221) );
AOI222xp33_ASAP7_75t_L g1222 ( .A1(n_1205), .A2(n_1159), .B1(n_1152), .B2(n_1180), .C1(n_1132), .C2(n_1176), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_1207), .A2(n_1184), .B1(n_1188), .B2(n_1107), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1209), .Y(n_1224) );
NAND3xp33_ASAP7_75t_SL g1225 ( .A(n_1213), .B(n_1200), .C(n_1156), .Y(n_1225) );
AOI221xp5_ASAP7_75t_L g1226 ( .A1(n_1204), .A2(n_1162), .B1(n_1175), .B2(n_1174), .C(n_1164), .Y(n_1226) );
AOI31xp33_ASAP7_75t_L g1227 ( .A1(n_1218), .A2(n_1214), .A3(n_1217), .B(n_1208), .Y(n_1227) );
INVx1_ASAP7_75t_SL g1228 ( .A(n_1220), .Y(n_1228) );
NAND4xp25_ASAP7_75t_L g1229 ( .A(n_1223), .B(n_1207), .C(n_1013), .D(n_1083), .Y(n_1229) );
AOI221xp5_ASAP7_75t_L g1230 ( .A1(n_1225), .A2(n_1215), .B1(n_1207), .B2(n_1211), .C(n_1212), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1231 ( .A1(n_1226), .A2(n_1206), .B1(n_1071), .B2(n_1210), .Y(n_1231) );
AOI21xp5_ASAP7_75t_L g1232 ( .A1(n_1219), .A2(n_1221), .B(n_1222), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1224), .Y(n_1233) );
AND2x4_ASAP7_75t_L g1234 ( .A(n_1228), .B(n_993), .Y(n_1234) );
NAND4xp75_ASAP7_75t_L g1235 ( .A(n_1232), .B(n_993), .C(n_1206), .D(n_1090), .Y(n_1235) );
NAND2x1_ASAP7_75t_L g1236 ( .A(n_1227), .B(n_1115), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1233), .B(n_1172), .Y(n_1237) );
AOI21xp5_ASAP7_75t_L g1238 ( .A1(n_1229), .A2(n_1055), .B(n_1070), .Y(n_1238) );
INVx2_ASAP7_75t_L g1239 ( .A(n_1234), .Y(n_1239) );
NAND3xp33_ASAP7_75t_SL g1240 ( .A(n_1236), .B(n_1230), .C(n_1231), .Y(n_1240) );
NOR4xp25_ASAP7_75t_L g1241 ( .A(n_1235), .B(n_1088), .C(n_1076), .D(n_1079), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1237), .B(n_1105), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1239), .B(n_1238), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1242), .Y(n_1244) );
INVx4_ASAP7_75t_L g1245 ( .A(n_1241), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1243), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1244), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1246), .Y(n_1248) );
OAI22x1_ASAP7_75t_L g1249 ( .A1(n_1247), .A2(n_1245), .B1(n_1240), .B2(n_983), .Y(n_1249) );
AOI21xp33_ASAP7_75t_SL g1250 ( .A1(n_1249), .A2(n_983), .B(n_1081), .Y(n_1250) );
AOI22xp5_ASAP7_75t_L g1251 ( .A1(n_1248), .A2(n_983), .B1(n_1083), .B2(n_1055), .Y(n_1251) );
AOI22x1_ASAP7_75t_L g1252 ( .A1(n_1250), .A2(n_987), .B1(n_991), .B2(n_1079), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1253 ( .A1(n_1252), .A2(n_1251), .B1(n_1161), .B2(n_1115), .Y(n_1253) );
endmodule