module fake_jpeg_6858_n_19 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_19;

wire n_13;
wire n_14;
wire n_18;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_7),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_8),
.C(n_10),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_0),
.Y(n_15)
);

FAx1_ASAP7_75t_SL g18 ( 
.A(n_15),
.B(n_16),
.CI(n_17),
.CON(n_18),
.SN(n_18)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_11),
.A2(n_2),
.B(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

AOI21x1_ASAP7_75t_SL g19 ( 
.A1(n_18),
.A2(n_12),
.B(n_9),
.Y(n_19)
);


endmodule