module fake_ibex_1494_n_794 (n_85, n_128, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_106, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_91, n_54, n_19, n_794);

input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_794;

wire n_151;
wire n_599;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_738;
wire n_475;
wire n_166;
wire n_163;
wire n_753;
wire n_747;
wire n_500;
wire n_645;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_383;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_772;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_788;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_706;
wire n_624;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_728;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_159;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_47),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_24),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_15),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_86),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_42),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_7),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_41),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_37),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_9),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_10),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_99),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_23),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_28),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_95),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_115),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_116),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_43),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_54),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_78),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_L g186 ( 
.A(n_121),
.B(n_92),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_117),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_74),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_133),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_94),
.B(n_135),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_62),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_30),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_11),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_72),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_89),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_22),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_88),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_23),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_44),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_68),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_45),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_80),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_35),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_26),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_111),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_46),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_61),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_55),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_131),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_122),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_60),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_113),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_7),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_39),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_66),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_5),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_102),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_4),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_141),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_19),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_2),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_56),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_48),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_69),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_130),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_112),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_27),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_104),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_40),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

OA21x2_ASAP7_75t_L g242 ( 
.A1(n_143),
.A2(n_67),
.B(n_139),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_0),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_166),
.B(n_1),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_148),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_155),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_155),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_144),
.A2(n_70),
.B(n_138),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_155),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_202),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_182),
.B(n_2),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_177),
.A2(n_73),
.B(n_137),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_145),
.A2(n_65),
.B(n_136),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_207),
.B(n_3),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_173),
.B(n_3),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_148),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_148),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_202),
.Y(n_270)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_148),
.Y(n_271)
);

XNOR2x2_ASAP7_75t_R g272 ( 
.A(n_147),
.B(n_6),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_180),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_149),
.A2(n_64),
.B(n_134),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_148),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_178),
.B(n_6),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_176),
.B(n_8),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_193),
.B(n_9),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_147),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_189),
.B(n_12),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_201),
.Y(n_282)
);

OAI22x1_ASAP7_75t_L g283 ( 
.A1(n_222),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_168),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_150),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_206),
.B(n_209),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g288 ( 
.A(n_151),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_169),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_168),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_174),
.Y(n_292)
);

CKINVDCx11_ASAP7_75t_R g293 ( 
.A(n_174),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_152),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_154),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_168),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_156),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_159),
.B(n_16),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_168),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_160),
.B(n_32),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_298),
.A2(n_222),
.B1(n_181),
.B2(n_237),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_293),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_244),
.B(n_175),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g309 ( 
.A1(n_283),
.A2(n_232),
.B1(n_228),
.B2(n_225),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_251),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_246),
.B(n_230),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

NOR2x1p5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_181),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_163),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_249),
.B(n_146),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_300),
.A2(n_204),
.B1(n_239),
.B2(n_164),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_287),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_277),
.B(n_167),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_253),
.A2(n_249),
.B1(n_273),
.B2(n_251),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_263),
.Y(n_331)
);

OR2x6_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_186),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_230),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_293),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_291),
.B(n_172),
.Y(n_341)
);

AND2x4_ASAP7_75t_SL g342 ( 
.A(n_281),
.B(n_240),
.Y(n_342)
);

NAND2xp33_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_190),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_276),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_273),
.A2(n_240),
.B1(n_205),
.B2(n_226),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_288),
.A2(n_226),
.B1(n_205),
.B2(n_203),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_243),
.B(n_157),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_292),
.Y(n_353)
);

AND2x6_ASAP7_75t_L g354 ( 
.A(n_250),
.B(n_179),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_243),
.B(n_162),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_245),
.B(n_195),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_286),
.B(n_196),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_252),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_261),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_269),
.B(n_294),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_R g361 ( 
.A(n_269),
.B(n_153),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_295),
.B(n_198),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_255),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_265),
.Y(n_364)
);

INVx8_ASAP7_75t_L g365 ( 
.A(n_300),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_343),
.C(n_302),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_302),
.A2(n_158),
.B1(n_188),
.B2(n_212),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_347),
.A2(n_300),
.B1(n_283),
.B2(n_224),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_359),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_280),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_360),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_307),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_351),
.A2(n_223),
.B1(n_220),
.B2(n_210),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_360),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_318),
.B(n_217),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_320),
.B(n_194),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_315),
.B(n_262),
.Y(n_384)
);

BUFx4_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_329),
.A2(n_211),
.B1(n_213),
.B2(n_215),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g388 ( 
.A(n_318),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_303),
.B(n_183),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_184),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_336),
.B(n_187),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_306),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_327),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_316),
.B(n_229),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_233),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_274),
.B(n_234),
.C(n_191),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_SL g399 ( 
.A(n_365),
.B(n_214),
.Y(n_399)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_354),
.B(n_216),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_308),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_308),
.Y(n_405)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_354),
.B(n_218),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_313),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_304),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_312),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_354),
.B(n_221),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_355),
.B(n_227),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_231),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_332),
.A2(n_235),
.B1(n_236),
.B2(n_242),
.Y(n_416)
);

AND2x6_ASAP7_75t_SL g417 ( 
.A(n_340),
.B(n_272),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_342),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_356),
.B(n_242),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_242),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_357),
.A2(n_258),
.B1(n_264),
.B2(n_270),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_258),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_L g423 ( 
.A(n_309),
.B(n_272),
.C(n_18),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_319),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_319),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_321),
.Y(n_426)
);

AND2x4_ASAP7_75t_SL g427 ( 
.A(n_332),
.B(n_257),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_330),
.A2(n_309),
.B1(n_344),
.B2(n_346),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_361),
.B(n_17),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_417),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_373),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_388),
.B(n_310),
.Y(n_434)
);

AO21x1_ASAP7_75t_L g435 ( 
.A1(n_420),
.A2(n_419),
.B(n_384),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_400),
.B(n_301),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_372),
.B(n_321),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_382),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_419),
.A2(n_420),
.B(n_422),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_390),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_394),
.B(n_326),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_387),
.B(n_335),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_345),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_333),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_366),
.B(n_339),
.Y(n_446)
);

BUFx5_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_377),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_379),
.B(n_17),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_371),
.B(n_18),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_368),
.B(n_20),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_381),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_20),
.Y(n_456)
);

CKINVDCx8_ASAP7_75t_R g457 ( 
.A(n_385),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_374),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_400),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_429),
.A2(n_406),
.B1(n_380),
.B2(n_413),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_410),
.B(n_21),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_375),
.B(n_24),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_406),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_386),
.B(n_25),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_396),
.A2(n_397),
.B(n_391),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_389),
.B(n_25),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_406),
.A2(n_369),
.B1(n_430),
.B2(n_423),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_402),
.A2(n_259),
.B1(n_260),
.B2(n_270),
.Y(n_470)
);

AO32x1_ASAP7_75t_L g471 ( 
.A1(n_427),
.A2(n_270),
.A3(n_363),
.B1(n_29),
.B2(n_30),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_428),
.Y(n_473)
);

NAND2x1p5_ASAP7_75t_L g474 ( 
.A(n_399),
.B(n_28),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_416),
.A2(n_29),
.B(n_31),
.C(n_33),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_402),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_421),
.A2(n_426),
.B(n_425),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_392),
.Y(n_478)
);

OAI321xp33_ASAP7_75t_L g479 ( 
.A1(n_408),
.A2(n_49),
.A3(n_50),
.B1(n_51),
.B2(n_52),
.C(n_53),
.Y(n_479)
);

AOI33xp33_ASAP7_75t_L g480 ( 
.A1(n_405),
.A2(n_424),
.A3(n_407),
.B1(n_409),
.B2(n_401),
.B3(n_395),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_408),
.A2(n_412),
.B1(n_415),
.B2(n_414),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_412),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_367),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_457),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_444),
.B(n_91),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_431),
.B(n_98),
.Y(n_487)
);

NAND3xp33_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_101),
.C(n_103),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_454),
.Y(n_489)
);

AOI211x1_ASAP7_75t_L g490 ( 
.A1(n_435),
.A2(n_105),
.B(n_106),
.C(n_108),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_432),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_440),
.Y(n_492)
);

CKINVDCx6p67_ASAP7_75t_R g493 ( 
.A(n_462),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_460),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

INVx2_ASAP7_75t_R g496 ( 
.A(n_472),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_455),
.B(n_478),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_474),
.Y(n_498)
);

AND3x1_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_468),
.C(n_461),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_451),
.B(n_449),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_433),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_466),
.Y(n_502)
);

BUFx2_ASAP7_75t_R g503 ( 
.A(n_463),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_456),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_460),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_473),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_447),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_445),
.Y(n_508)
);

NOR4xp25_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_441),
.C(n_442),
.D(n_437),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_434),
.B(n_443),
.Y(n_510)
);

INVx3_ASAP7_75t_SL g511 ( 
.A(n_447),
.Y(n_511)
);

INVx6_ASAP7_75t_L g512 ( 
.A(n_438),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_480),
.A2(n_465),
.B(n_436),
.C(n_453),
.Y(n_513)
);

AOI21x1_ASAP7_75t_L g514 ( 
.A1(n_471),
.A2(n_438),
.B(n_453),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_465),
.A2(n_471),
.B(n_459),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_459),
.A2(n_477),
.B(n_439),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_459),
.A2(n_477),
.B(n_439),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_440),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_439),
.A2(n_467),
.B(n_398),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_444),
.B(n_349),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_440),
.Y(n_522)
);

BUFx2_ASAP7_75t_SL g523 ( 
.A(n_457),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_460),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_440),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_458),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_431),
.B(n_370),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_457),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_431),
.B(n_448),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_458),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_431),
.B(n_370),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_460),
.Y(n_532)
);

CKINVDCx11_ASAP7_75t_R g533 ( 
.A(n_457),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_431),
.B(n_393),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_431),
.B(n_370),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_431),
.B(n_370),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_431),
.B(n_370),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_457),
.B(n_349),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_431),
.B(n_448),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_444),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_431),
.B(n_370),
.Y(n_541)
);

OAI22x1_ASAP7_75t_L g542 ( 
.A1(n_452),
.A2(n_292),
.B1(n_310),
.B2(n_353),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_431),
.B(n_370),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_450),
.Y(n_544)
);

AO31x2_ASAP7_75t_L g545 ( 
.A1(n_435),
.A2(n_439),
.A3(n_398),
.B(n_419),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_458),
.Y(n_546)
);

AO32x2_ASAP7_75t_L g547 ( 
.A1(n_476),
.A2(n_483),
.A3(n_470),
.B1(n_481),
.B2(n_471),
.Y(n_547)
);

AO31x2_ASAP7_75t_L g548 ( 
.A1(n_435),
.A2(n_439),
.A3(n_398),
.B(n_419),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_450),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_450),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_540),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_492),
.B(n_519),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_522),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_525),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_544),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_521),
.B(n_534),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_495),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_527),
.B(n_531),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_526),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_546),
.Y(n_561)
);

INVx6_ASAP7_75t_L g562 ( 
.A(n_485),
.Y(n_562)
);

OA21x2_ASAP7_75t_L g563 ( 
.A1(n_515),
.A2(n_516),
.B(n_514),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_485),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g565 ( 
.A1(n_515),
.A2(n_520),
.B(n_509),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_500),
.A2(n_499),
.B1(n_493),
.B2(n_511),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_529),
.B(n_539),
.Y(n_567)
);

BUFx2_ASAP7_75t_SL g568 ( 
.A(n_484),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_501),
.Y(n_569)
);

BUFx10_ASAP7_75t_L g570 ( 
.A(n_550),
.Y(n_570)
);

NOR2x1_ASAP7_75t_SL g571 ( 
.A(n_524),
.B(n_523),
.Y(n_571)
);

NAND4xp25_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_541),
.C(n_543),
.D(n_535),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_524),
.B(n_498),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_524),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_549),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_536),
.B(n_537),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_499),
.A2(n_502),
.B1(n_504),
.B2(n_486),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_494),
.B(n_508),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_491),
.Y(n_579)
);

INVx8_ASAP7_75t_L g580 ( 
.A(n_528),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_487),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_510),
.B(n_542),
.Y(n_582)
);

BUFx2_ASAP7_75t_R g583 ( 
.A(n_533),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_489),
.Y(n_584)
);

AO21x2_ASAP7_75t_L g585 ( 
.A1(n_509),
.A2(n_513),
.B(n_488),
.Y(n_585)
);

INVx3_ASAP7_75t_SL g586 ( 
.A(n_512),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_532),
.B(n_505),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_503),
.B(n_496),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_490),
.B(n_532),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_548),
.B(n_512),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_547),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_547),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_540),
.B(n_534),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_521),
.B(n_349),
.Y(n_595)
);

AO21x2_ASAP7_75t_L g596 ( 
.A1(n_516),
.A2(n_515),
.B(n_514),
.Y(n_596)
);

OA21x2_ASAP7_75t_L g597 ( 
.A1(n_515),
.A2(n_518),
.B(n_517),
.Y(n_597)
);

CKINVDCx12_ASAP7_75t_R g598 ( 
.A(n_533),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_544),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_492),
.B(n_519),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_506),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_492),
.B(n_519),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_492),
.B(n_519),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_540),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_534),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_534),
.A2(n_455),
.B1(n_497),
.B2(n_431),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_524),
.B(n_450),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_534),
.A2(n_455),
.B1(n_497),
.B2(n_431),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_540),
.B(n_534),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_511),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_534),
.A2(n_455),
.B1(n_497),
.B2(n_431),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_507),
.B(n_460),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_540),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_540),
.B(n_534),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_484),
.Y(n_616)
);

AOI21xp33_ASAP7_75t_SL g617 ( 
.A1(n_542),
.A2(n_349),
.B(n_348),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_540),
.B(n_393),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_533),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_591),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_601),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_601),
.Y(n_622)
);

INVx3_ASAP7_75t_SL g623 ( 
.A(n_567),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_562),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_559),
.B(n_560),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_597),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_562),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_619),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_559),
.B(n_560),
.Y(n_629)
);

BUFx4f_ASAP7_75t_SL g630 ( 
.A(n_579),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_602),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_602),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_553),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_553),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_561),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_558),
.B(n_576),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_595),
.B(n_556),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_573),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_611),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_554),
.B(n_557),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_554),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_572),
.A2(n_577),
.B1(n_605),
.B2(n_609),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_573),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_552),
.B(n_600),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_603),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_569),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_570),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_606),
.B(n_612),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_614),
.B(n_565),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_618),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_594),
.B(n_615),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_551),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_565),
.B(n_593),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_592),
.B(n_593),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_604),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_592),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_584),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_608),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_563),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_563),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_613),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_610),
.B(n_581),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_590),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_596),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_587),
.B(n_590),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_596),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_585),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_566),
.B(n_578),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_574),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_636),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_659),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_657),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_646),
.B(n_582),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_660),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_631),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_620),
.B(n_564),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_651),
.B(n_555),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_652),
.B(n_617),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_655),
.B(n_625),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_664),
.B(n_617),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_655),
.B(n_589),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_665),
.B(n_607),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_642),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_660),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_658),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_651),
.B(n_599),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_650),
.A2(n_575),
.B1(n_607),
.B2(n_568),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_665),
.B(n_613),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_629),
.B(n_570),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_650),
.B(n_586),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_667),
.B(n_571),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_629),
.B(n_616),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_635),
.B(n_580),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_656),
.B(n_583),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_637),
.B(n_580),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_656),
.B(n_580),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_661),
.B(n_579),
.Y(n_699)
);

NOR2x1_ASAP7_75t_L g700 ( 
.A(n_671),
.B(n_598),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_643),
.A2(n_670),
.B1(n_664),
.B2(n_632),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_621),
.B(n_622),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_626),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_661),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_633),
.B(n_641),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_634),
.B(n_640),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_662),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_671),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_674),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_681),
.B(n_669),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_685),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_681),
.B(n_669),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_703),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_683),
.B(n_666),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_708),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_708),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_683),
.B(n_706),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_706),
.B(n_668),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_699),
.B(n_663),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_699),
.B(n_702),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_679),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_679),
.B(n_653),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_709),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_715),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_721),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_720),
.B(n_687),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_717),
.B(n_682),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_711),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_712),
.B(n_688),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_713),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_717),
.B(n_710),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_710),
.B(n_673),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_722),
.B(n_675),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_720),
.B(n_690),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_714),
.B(n_704),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_718),
.B(n_707),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_722),
.B(n_705),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_724),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_723),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_728),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_730),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_726),
.A2(n_720),
.B1(n_696),
.B2(n_680),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_729),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_732),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_726),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_725),
.B(n_716),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_735),
.B(n_736),
.Y(n_747)
);

OAI21xp33_ASAP7_75t_L g748 ( 
.A1(n_742),
.A2(n_727),
.B(n_696),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_741),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_729),
.B1(n_731),
.B2(n_726),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_740),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_738),
.B(n_739),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_743),
.B(n_736),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_743),
.A2(n_734),
.B1(n_697),
.B2(n_672),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_740),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_738),
.A2(n_700),
.B(n_691),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_747),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_747),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_756),
.A2(n_745),
.B(n_734),
.C(n_686),
.Y(n_759)
);

AOI211xp5_ASAP7_75t_SL g760 ( 
.A1(n_748),
.A2(n_630),
.B(n_692),
.C(n_670),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_L g761 ( 
.A1(n_750),
.A2(n_744),
.B1(n_746),
.B2(n_733),
.C(n_737),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_756),
.B(n_628),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_759),
.B(n_757),
.Y(n_763)
);

AOI221xp5_ASAP7_75t_L g764 ( 
.A1(n_761),
.A2(n_752),
.B1(n_754),
.B2(n_758),
.C(n_755),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_760),
.B(n_751),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_765),
.B(n_762),
.C(n_628),
.Y(n_766)
);

AND4x1_ASAP7_75t_L g767 ( 
.A(n_764),
.B(n_689),
.C(n_701),
.D(n_698),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_766),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_767),
.B(n_763),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_768),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_769),
.B(n_753),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_770),
.B(n_649),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_771),
.A2(n_745),
.B1(n_694),
.B2(n_649),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_773),
.A2(n_686),
.B1(n_676),
.B2(n_654),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_SL g775 ( 
.A1(n_772),
.A2(n_676),
.B1(n_624),
.B2(n_627),
.Y(n_775)
);

XOR2xp5_ASAP7_75t_L g776 ( 
.A(n_773),
.B(n_692),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_SL g777 ( 
.A1(n_774),
.A2(n_624),
.B(n_627),
.C(n_695),
.Y(n_777)
);

OA22x2_ASAP7_75t_L g778 ( 
.A1(n_775),
.A2(n_694),
.B1(n_698),
.B2(n_623),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_776),
.Y(n_779)
);

NOR3xp33_ASAP7_75t_L g780 ( 
.A(n_775),
.B(n_648),
.C(n_639),
.Y(n_780)
);

AOI21x1_ASAP7_75t_L g781 ( 
.A1(n_776),
.A2(n_691),
.B(n_645),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_779),
.A2(n_695),
.B(n_647),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_777),
.B(n_648),
.C(n_639),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_781),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_778),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_780),
.A2(n_693),
.B1(n_644),
.B2(n_638),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_779),
.A2(n_693),
.B1(n_677),
.B2(n_749),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_785),
.A2(n_693),
.B1(n_678),
.B2(n_719),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_784),
.B(n_782),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_787),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_790),
.A2(n_783),
.B1(n_786),
.B2(n_684),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_789),
.A2(n_639),
.B(n_648),
.Y(n_792)
);

OR2x6_ASAP7_75t_L g793 ( 
.A(n_792),
.B(n_788),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_793),
.A2(n_791),
.B1(n_684),
.B2(n_734),
.Y(n_794)
);


endmodule