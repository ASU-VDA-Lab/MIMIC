module fake_netlist_6_51_n_2015 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2015);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2015;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_56),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_32),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_121),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_68),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_68),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_39),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_116),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_137),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_36),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_21),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_22),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_8),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_48),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_119),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_130),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_146),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_78),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_8),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_163),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_37),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_115),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_187),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_143),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_1),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_145),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_183),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_76),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_76),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_66),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_127),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_48),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_73),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_18),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_92),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_36),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_60),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_100),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_114),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_107),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_160),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_166),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_171),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_152),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_122),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_154),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_139),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_106),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_108),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_61),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_186),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_61),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_59),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_91),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_58),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_124),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_43),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_30),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_53),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_60),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_193),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_174),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_98),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_189),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_27),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_19),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_63),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_6),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_80),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_141),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_131),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_109),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_84),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_52),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_56),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_142),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_88),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_41),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_15),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_94),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_74),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_63),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_103),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_34),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_1),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_117),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_105),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_102),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_23),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_35),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_136),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_165),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_3),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_132),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_198),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_28),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_134),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_97),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_40),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_62),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_93),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_85),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_155),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_39),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_75),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_49),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_12),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_37),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_49),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_44),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_79),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_28),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_149),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_172),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_15),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_30),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_22),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_44),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_96),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_47),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_144),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_113),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_31),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_6),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_14),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_120),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_101),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_173),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_184),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_133),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_27),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_81),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_194),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_10),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_66),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_75),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_151),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_2),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_157),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_41),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_31),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_95),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_167),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_77),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_50),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_192),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_104),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_50),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_42),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_118),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_23),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_52),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_190),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_54),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_7),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_67),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_125),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_99),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_14),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_53),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_0),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_26),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_170),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_54),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_159),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_135),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_62),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_111),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_162),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_112),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_90),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_24),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_47),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_67),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_9),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_16),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_29),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_29),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_16),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_24),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_180),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_35),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_0),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_18),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_2),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_391),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_200),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_391),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_391),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_201),
.B(n_3),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_202),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_391),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_318),
.B(n_4),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_263),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_204),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_282),
.B(n_4),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_312),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_208),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_209),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_212),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_346),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_282),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_221),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_266),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_266),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_346),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_222),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_301),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_227),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_301),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_199),
.B(n_5),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_326),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_231),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_201),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_213),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_213),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_234),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_240),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_234),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_230),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_210),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_230),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_239),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_232),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_274),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_210),
.B(n_5),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_239),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_216),
.B(n_7),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_235),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_211),
.B(n_9),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_287),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_211),
.B(n_10),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_228),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_242),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_236),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_244),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_242),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_268),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_297),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_268),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_269),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_305),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_269),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_324),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_276),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_219),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_233),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_247),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_223),
.B(n_11),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_203),
.B(n_11),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_276),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_248),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_219),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_350),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_233),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_223),
.B(n_12),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_251),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_350),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_277),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_277),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_252),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_240),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_286),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_298),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_278),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_286),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_254),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_216),
.B(n_13),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_290),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_255),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_290),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_292),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_257),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_292),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_265),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_271),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g490 ( 
.A(n_304),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_304),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_307),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_307),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_298),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_317),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_272),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_280),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_317),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_283),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_404),
.B(n_225),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_431),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_441),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_407),
.B(n_225),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_399),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

NOR2x1_ASAP7_75t_L g508 ( 
.A(n_463),
.B(n_303),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_435),
.B(n_460),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_400),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_403),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_459),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_468),
.B(n_288),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_477),
.B(n_303),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_397),
.B(n_203),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_431),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_414),
.B(n_205),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_403),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_409),
.A2(n_334),
.B(n_320),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_409),
.B(n_220),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_475),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_416),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_466),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_416),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_417),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_291),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_439),
.B(n_220),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_417),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_420),
.Y(n_532)
);

CKINVDCx6p67_ASAP7_75t_R g533 ( 
.A(n_480),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_434),
.A2(n_226),
.B(n_224),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_427),
.B(n_224),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_446),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_422),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_422),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_443),
.B(n_302),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_445),
.B(n_306),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_423),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_423),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_433),
.B(n_206),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_425),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_462),
.B(n_308),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_425),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_433),
.B(n_206),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_469),
.B(n_309),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_401),
.A2(n_229),
.B(n_226),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_427),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_424),
.B(n_241),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_428),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_428),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_429),
.B(n_330),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_429),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_401),
.B(n_241),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_430),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_432),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_413),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

BUFx8_ASAP7_75t_L g564 ( 
.A(n_436),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_440),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_440),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_447),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_447),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_450),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_418),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_451),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_453),
.B(n_323),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_453),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_471),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_456),
.B(n_332),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_398),
.B(n_218),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_456),
.B(n_333),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_557),
.A2(n_408),
.B1(n_328),
.B2(n_371),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_522),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_513),
.B(n_527),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_502),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

NOR2x1p5_ASAP7_75t_L g585 ( 
.A(n_533),
.B(n_323),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_502),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_522),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_522),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_515),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_515),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_513),
.B(n_402),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_508),
.B(n_249),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_522),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_SL g594 ( 
.A(n_500),
.B(n_499),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_543),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_502),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_509),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_515),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_509),
.B(n_406),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_514),
.B(n_458),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_501),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_514),
.B(n_458),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_508),
.B(n_249),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_503),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_528),
.B(n_410),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_549),
.B(n_229),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_503),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_503),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_527),
.B(n_411),
.Y(n_611)
);

CKINVDCx11_ASAP7_75t_R g612 ( 
.A(n_533),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_503),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_528),
.A2(n_359),
.B1(n_342),
.B2(n_334),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_515),
.Y(n_615)
);

BUFx4f_ASAP7_75t_L g616 ( 
.A(n_520),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_515),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_520),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_520),
.Y(n_619)
);

INVxp67_ASAP7_75t_R g620 ( 
.A(n_562),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_520),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_502),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_502),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_502),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_SL g625 ( 
.A(n_500),
.B(n_483),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_502),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_517),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_539),
.B(n_412),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_536),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_536),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_504),
.B(n_415),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_549),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_528),
.A2(n_359),
.B1(n_342),
.B2(n_335),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_528),
.A2(n_335),
.B1(n_363),
.B2(n_320),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_516),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_516),
.Y(n_637)
);

AND3x2_ASAP7_75t_L g638 ( 
.A(n_504),
.B(n_258),
.C(n_530),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_533),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_530),
.B(n_419),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_512),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_562),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_516),
.Y(n_643)
);

AND2x2_ASAP7_75t_SL g644 ( 
.A(n_539),
.B(n_249),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_570),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_540),
.B(n_421),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_540),
.B(n_426),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_570),
.B(n_478),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_517),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_545),
.B(n_437),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_517),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_516),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_517),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_517),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_545),
.B(n_442),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_528),
.A2(n_363),
.B1(n_373),
.B2(n_372),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_549),
.B(n_253),
.Y(n_657)
);

AND3x2_ASAP7_75t_L g658 ( 
.A(n_518),
.B(n_256),
.C(n_253),
.Y(n_658)
);

BUFx4f_ASAP7_75t_L g659 ( 
.A(n_528),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_548),
.B(n_448),
.Y(n_660)
);

BUFx8_ASAP7_75t_SL g661 ( 
.A(n_512),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_517),
.Y(n_662)
);

INVx4_ASAP7_75t_SL g663 ( 
.A(n_528),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_528),
.A2(n_373),
.B1(n_383),
.B2(n_390),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_518),
.B(n_449),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_543),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_528),
.B(n_461),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_514),
.B(n_464),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_543),
.B(n_464),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_528),
.A2(n_378),
.B1(n_372),
.B2(n_383),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_548),
.B(n_465),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_517),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_574),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_516),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_564),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g676 ( 
.A(n_528),
.B(n_470),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_517),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_547),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_564),
.B(n_474),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_501),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_552),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_555),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_501),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_486),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_506),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_506),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_555),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_555),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_512),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_578),
.B(n_496),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_555),
.Y(n_691)
);

CKINVDCx6p67_ASAP7_75t_R g692 ( 
.A(n_524),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_578),
.B(n_488),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_552),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_551),
.B(n_489),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_555),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_564),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_552),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_557),
.A2(n_378),
.B1(n_390),
.B2(n_396),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_555),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_561),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_524),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_L g703 ( 
.A(n_554),
.B(n_249),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_555),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_505),
.A2(n_396),
.B1(n_490),
.B2(n_284),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_561),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_561),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_572),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_524),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_551),
.B(n_497),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_555),
.Y(n_711)
);

BUFx8_ASAP7_75t_SL g712 ( 
.A(n_556),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_505),
.B(n_256),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_535),
.B(n_267),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_547),
.B(n_472),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_572),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_560),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_572),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_560),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_564),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_573),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_564),
.B(n_218),
.Y(n_722)
);

BUFx4f_ASAP7_75t_L g723 ( 
.A(n_560),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_506),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_573),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_554),
.B(n_405),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_534),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_521),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_573),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_507),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_556),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_579),
.A2(n_215),
.B1(n_336),
.B2(n_331),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_589),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_644),
.A2(n_535),
.B1(n_534),
.B2(n_521),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_630),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_600),
.B(n_438),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_693),
.B(n_576),
.C(n_556),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_629),
.B(n_444),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_598),
.B(n_577),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_589),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_582),
.B(n_577),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_647),
.B(n_671),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_690),
.A2(n_455),
.B1(n_457),
.B2(n_452),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_630),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_644),
.B(n_579),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_659),
.B(n_249),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_659),
.B(n_644),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_713),
.A2(n_535),
.B1(n_534),
.B2(n_521),
.Y(n_748)
);

NOR2x2_ASAP7_75t_L g749 ( 
.A(n_713),
.B(n_576),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_631),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_681),
.Y(n_751)
);

NOR2x1p5_ASAP7_75t_L g752 ( 
.A(n_648),
.B(n_692),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_646),
.B(n_558),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_590),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_726),
.A2(n_596),
.B1(n_678),
.B2(n_666),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_642),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_650),
.B(n_558),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_659),
.A2(n_521),
.B(n_535),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_655),
.B(n_558),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_694),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_660),
.B(n_558),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_673),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_590),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_705),
.B(n_574),
.C(n_454),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_636),
.B(n_558),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_636),
.B(n_535),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_673),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_637),
.B(n_535),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_659),
.B(n_294),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_637),
.B(n_560),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_713),
.A2(n_521),
.B1(n_560),
.B2(n_281),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_612),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_713),
.B(n_576),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_595),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_618),
.B(n_619),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_648),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_643),
.B(n_560),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_618),
.A2(n_575),
.B(n_563),
.C(n_567),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_643),
.B(n_560),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_591),
.B(n_250),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_595),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_599),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_652),
.B(n_560),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_620),
.B(n_574),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_694),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_652),
.B(n_521),
.Y(n_786)
);

BUFx4f_ASAP7_75t_L g787 ( 
.A(n_713),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_674),
.B(n_526),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_616),
.B(n_294),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_642),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_698),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_596),
.B(n_563),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_645),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_616),
.B(n_294),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_620),
.B(n_567),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_599),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_611),
.B(n_260),
.Y(n_797)
);

O2A1O1Ixp5_ASAP7_75t_L g798 ( 
.A1(n_616),
.A2(n_507),
.B(n_510),
.C(n_511),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_728),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_698),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_674),
.B(n_526),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_701),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_601),
.B(n_526),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_669),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_669),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_639),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_616),
.B(n_633),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_601),
.B(n_526),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_603),
.B(n_526),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_603),
.B(n_541),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_668),
.B(n_541),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_633),
.B(n_294),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_633),
.B(n_294),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_584),
.B(n_240),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_668),
.B(n_541),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_679),
.B(n_575),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_666),
.B(n_267),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_584),
.A2(n_325),
.B1(n_273),
.B2(n_281),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_678),
.B(n_722),
.Y(n_819)
);

BUFx6f_ASAP7_75t_SL g820 ( 
.A(n_714),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_701),
.B(n_541),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_706),
.B(n_541),
.Y(n_822)
);

AND2x2_ASAP7_75t_SL g823 ( 
.A(n_614),
.B(n_273),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_706),
.B(n_707),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_645),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_665),
.B(n_355),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_615),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_684),
.A2(n_584),
.B1(n_617),
.B2(n_615),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_707),
.B(n_550),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_663),
.B(n_240),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_617),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_708),
.B(n_550),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_728),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_663),
.B(n_240),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_663),
.B(n_240),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_728),
.Y(n_836)
);

OAI221xp5_ASAP7_75t_L g837 ( 
.A1(n_699),
.A2(n_358),
.B1(n_354),
.B2(n_353),
.C(n_299),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_715),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_708),
.B(n_550),
.Y(n_839)
);

AOI221xp5_ASAP7_75t_L g840 ( 
.A1(n_580),
.A2(n_289),
.B1(n_352),
.B2(n_388),
.C(n_321),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_663),
.B(n_240),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_715),
.B(n_284),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_632),
.B(n_207),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_716),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_619),
.A2(n_325),
.B(n_313),
.C(n_314),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_718),
.B(n_553),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_718),
.B(n_553),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_SL g848 ( 
.A(n_641),
.B(n_218),
.Y(n_848)
);

AND2x6_ASAP7_75t_L g849 ( 
.A(n_675),
.B(n_299),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_721),
.B(n_553),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_580),
.B(n_295),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_594),
.A2(n_380),
.B1(n_377),
.B2(n_382),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_663),
.B(n_240),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_721),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_725),
.B(n_553),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_725),
.B(n_559),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_621),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_729),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_731),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_729),
.B(n_559),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_621),
.B(n_559),
.Y(n_861)
);

OAI22xp33_ASAP7_75t_L g862 ( 
.A1(n_607),
.A2(n_313),
.B1(n_314),
.B2(n_322),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_602),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_602),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_627),
.B(n_559),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_627),
.B(n_565),
.Y(n_866)
);

NAND3xp33_ASAP7_75t_SL g867 ( 
.A(n_689),
.B(n_217),
.C(n_214),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_730),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_714),
.B(n_565),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_714),
.B(n_240),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_597),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_640),
.B(n_237),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_714),
.B(n_565),
.Y(n_873)
);

NOR2xp67_ASAP7_75t_L g874 ( 
.A(n_732),
.B(n_525),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_624),
.B(n_565),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_638),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_730),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_583),
.B(n_566),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_583),
.B(n_566),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_695),
.B(n_525),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_680),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_658),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_585),
.B(n_322),
.Y(n_883)
);

BUFx6f_ASAP7_75t_SL g884 ( 
.A(n_592),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_SL g885 ( 
.A(n_702),
.B(n_218),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_597),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_635),
.A2(n_656),
.B1(n_670),
.B2(n_664),
.Y(n_887)
);

NAND2x1p5_ASAP7_75t_L g888 ( 
.A(n_675),
.B(n_337),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_680),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_634),
.A2(n_341),
.B1(n_376),
.B2(n_369),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_607),
.A2(n_341),
.B1(n_376),
.B2(n_369),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_710),
.B(n_238),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_683),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_720),
.B(n_622),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_720),
.B(n_338),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_607),
.A2(n_354),
.B1(n_353),
.B2(n_337),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_583),
.B(n_566),
.Y(n_897)
);

INVx8_ASAP7_75t_L g898 ( 
.A(n_607),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_583),
.B(n_566),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_683),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_677),
.B(n_622),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_677),
.B(n_568),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_744),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_758),
.A2(n_727),
.B(n_723),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_747),
.A2(n_723),
.B(n_667),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_742),
.B(n_625),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_741),
.B(n_592),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_799),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_787),
.B(n_675),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_751),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_805),
.B(n_585),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_747),
.A2(n_794),
.B(n_789),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_739),
.B(n_592),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_744),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_780),
.B(n_592),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_789),
.A2(n_723),
.B(n_676),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_797),
.A2(n_606),
.B(n_703),
.C(n_357),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_750),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_794),
.A2(n_723),
.B(n_586),
.Y(n_919)
);

OAI21xp33_ASAP7_75t_L g920 ( 
.A1(n_840),
.A2(n_245),
.B(n_243),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_751),
.Y(n_921)
);

BUFx4f_ASAP7_75t_L g922 ( 
.A(n_773),
.Y(n_922)
);

NAND2x1_ASAP7_75t_L g923 ( 
.A(n_871),
.B(n_677),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_786),
.A2(n_586),
.B(n_607),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_875),
.A2(n_586),
.B(n_657),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_807),
.A2(n_586),
.B(n_657),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_807),
.A2(n_657),
.B(n_682),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_762),
.B(n_592),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_861),
.A2(n_657),
.B(n_682),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_826),
.A2(n_357),
.B(n_623),
.C(n_626),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_762),
.A2(n_767),
.B(n_845),
.C(n_775),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_865),
.A2(n_866),
.B(n_768),
.Y(n_932)
);

BUFx4f_ASAP7_75t_L g933 ( 
.A(n_773),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_745),
.B(n_697),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_799),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_776),
.B(n_709),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_767),
.B(n_592),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_766),
.A2(n_657),
.B(n_682),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_736),
.B(n_692),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_775),
.A2(n_696),
.B(n_682),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_792),
.B(n_592),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_798),
.A2(n_623),
.B(n_622),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_799),
.B(n_623),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_816),
.A2(n_604),
.B1(n_677),
.B2(n_626),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_735),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_738),
.B(n_685),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_792),
.B(n_604),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_753),
.A2(n_696),
.B(n_608),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_792),
.B(n_604),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_799),
.B(n_757),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_759),
.A2(n_696),
.B(n_608),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_761),
.A2(n_696),
.B(n_608),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_804),
.B(n_604),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_869),
.A2(n_608),
.B(n_597),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_760),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_L g956 ( 
.A(n_867),
.B(n_259),
.C(n_246),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_804),
.B(n_604),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_760),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_756),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_833),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_785),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_803),
.B(n_604),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_859),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_785),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_836),
.B(n_626),
.Y(n_965)
);

CKINVDCx10_ASAP7_75t_R g966 ( 
.A(n_772),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_836),
.B(n_755),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_833),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_873),
.A2(n_777),
.B(n_770),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_L g970 ( 
.A(n_737),
.B(n_262),
.C(n_261),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_887),
.A2(n_818),
.B1(n_819),
.B2(n_734),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_808),
.B(n_604),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_790),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_809),
.B(n_628),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_793),
.B(n_685),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_779),
.A2(n_608),
.B(n_597),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_810),
.B(n_628),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_783),
.A2(n_608),
.B(n_597),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_812),
.A2(n_813),
.B(n_901),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_791),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_791),
.Y(n_981)
);

AO21x1_ASAP7_75t_L g982 ( 
.A1(n_812),
.A2(n_724),
.B(n_686),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_838),
.B(n_472),
.Y(n_983)
);

AOI222xp33_ASAP7_75t_L g984 ( 
.A1(n_851),
.A2(n_366),
.B1(n_295),
.B2(n_349),
.C1(n_347),
.C2(n_345),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_820),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_811),
.B(n_815),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_813),
.A2(n_654),
.B(n_597),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_814),
.A2(n_649),
.B(n_628),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_814),
.A2(n_651),
.B(n_649),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_788),
.A2(n_801),
.B(n_765),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_868),
.B(n_649),
.Y(n_991)
);

NOR2x1p5_ASAP7_75t_L g992 ( 
.A(n_772),
.B(n_661),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_894),
.A2(n_662),
.B(n_654),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_795),
.B(n_473),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_892),
.A2(n_651),
.B(n_653),
.C(n_672),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_894),
.A2(n_662),
.B(n_654),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_871),
.A2(n_662),
.B(n_654),
.Y(n_997)
);

AOI21x1_ASAP7_75t_L g998 ( 
.A1(n_746),
.A2(n_653),
.B(n_651),
.Y(n_998)
);

AO21x1_ASAP7_75t_L g999 ( 
.A1(n_828),
.A2(n_724),
.B(n_686),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_L g1000 ( 
.A(n_825),
.B(n_270),
.C(n_264),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_806),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_746),
.A2(n_672),
.B(n_653),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_823),
.A2(n_295),
.B1(n_366),
.B2(n_381),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_784),
.B(n_473),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_877),
.B(n_672),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_857),
.B(n_654),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_800),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_857),
.B(n_654),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_845),
.A2(n_581),
.B(n_588),
.C(n_587),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_871),
.A2(n_662),
.B(n_719),
.Y(n_1010)
);

AOI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_843),
.A2(n_279),
.B(n_275),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_769),
.A2(n_748),
.B(n_821),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_871),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_800),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_820),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_802),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_824),
.A2(n_662),
.B(n_719),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_802),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_769),
.A2(n_593),
.B(n_587),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_817),
.B(n_662),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_857),
.B(n_593),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_844),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_844),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_854),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_837),
.A2(n_581),
.B(n_587),
.C(n_588),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_817),
.B(n_700),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_733),
.B(n_700),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_830),
.A2(n_688),
.B(n_687),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_878),
.A2(n_688),
.B(n_687),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_740),
.B(n_700),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_817),
.B(n_700),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_778),
.A2(n_581),
.B(n_588),
.C(n_510),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_754),
.B(n_704),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_854),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_879),
.A2(n_719),
.B(n_688),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_819),
.A2(n_711),
.B1(n_691),
.B2(n_687),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_897),
.A2(n_711),
.B(n_691),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_763),
.B(n_774),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_842),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_L g1040 ( 
.A(n_872),
.B(n_293),
.C(n_285),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_820),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_874),
.A2(n_717),
.B(n_711),
.C(n_691),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_858),
.B(n_717),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_781),
.B(n_704),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_891),
.A2(n_717),
.B(n_613),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_898),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_858),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_880),
.A2(n_704),
.B1(n_340),
.B2(n_348),
.Y(n_1048)
);

AO21x1_ASAP7_75t_L g1049 ( 
.A1(n_862),
.A2(n_519),
.B(n_510),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_899),
.A2(n_704),
.B(n_605),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_782),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_863),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_796),
.B(n_568),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_743),
.B(n_295),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_842),
.B(n_366),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_827),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_831),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_819),
.A2(n_339),
.B1(n_343),
.B2(n_344),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_902),
.A2(n_613),
.B(n_610),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_773),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_886),
.A2(n_613),
.B(n_610),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_771),
.B(n_863),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_886),
.A2(n_610),
.B(n_609),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_817),
.B(n_764),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_842),
.B(n_476),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_864),
.B(n_893),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_819),
.A2(n_896),
.B1(n_898),
.B2(n_890),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_823),
.A2(n_366),
.B1(n_381),
.B2(n_568),
.Y(n_1068)
);

AO21x1_ASAP7_75t_L g1069 ( 
.A1(n_895),
.A2(n_511),
.B(n_519),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_773),
.B(n_296),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_882),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_895),
.A2(n_519),
.B(n_511),
.C(n_507),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_864),
.B(n_568),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_893),
.B(n_569),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_886),
.A2(n_609),
.B(n_605),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_900),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_L g1077 ( 
.A(n_898),
.B(n_361),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_898),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_848),
.B(n_476),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_822),
.A2(n_609),
.B(n_605),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_900),
.B(n_569),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_881),
.B(n_889),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_870),
.A2(n_571),
.B(n_569),
.C(n_525),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_852),
.A2(n_870),
.B(n_829),
.C(n_832),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_839),
.A2(n_571),
.B(n_569),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_876),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_846),
.B(n_571),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_847),
.B(n_364),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_850),
.Y(n_1089)
);

CKINVDCx6p67_ASAP7_75t_R g1090 ( 
.A(n_966),
.Y(n_1090)
);

AO32x2_ASAP7_75t_L g1091 ( 
.A1(n_971),
.A2(n_749),
.A3(n_888),
.B1(n_849),
.B2(n_860),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1007),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_906),
.A2(n_885),
.B(n_855),
.C(n_856),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_918),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_921),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_1011),
.B(n_806),
.C(n_830),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_906),
.A2(n_883),
.B1(n_752),
.B2(n_849),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1001),
.Y(n_1098)
);

OAI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1039),
.A2(n_883),
.B1(n_888),
.B2(n_749),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_SL g1100 ( 
.A1(n_939),
.A2(n_883),
.B1(n_315),
.B2(n_385),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1064),
.A2(n_834),
.B(n_853),
.C(n_841),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_963),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_967),
.A2(n_841),
.B(n_853),
.C(n_834),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1007),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1079),
.B(n_883),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_912),
.A2(n_835),
.B(n_884),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_992),
.Y(n_1107)
);

AO22x1_ASAP7_75t_L g1108 ( 
.A1(n_939),
.A2(n_1040),
.B1(n_936),
.B2(n_1054),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_914),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_916),
.A2(n_884),
.B(n_849),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_932),
.A2(n_904),
.B(n_986),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_958),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_946),
.B(n_849),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_946),
.A2(n_849),
.B1(n_392),
.B2(n_368),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_967),
.A2(n_532),
.B(n_537),
.C(n_538),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_914),
.Y(n_1116)
);

OAI21xp33_ASAP7_75t_L g1117 ( 
.A1(n_920),
.A2(n_393),
.B(n_310),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1047),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_936),
.B(n_712),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1047),
.Y(n_1120)
);

AO22x1_ASAP7_75t_L g1121 ( 
.A1(n_970),
.A2(n_386),
.B1(n_394),
.B2(n_375),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_905),
.A2(n_529),
.B(n_544),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_979),
.A2(n_529),
.B(n_544),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_924),
.A2(n_529),
.B(n_544),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_1064),
.A2(n_532),
.B(n_537),
.C(n_538),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_938),
.A2(n_925),
.B(n_929),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_961),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_970),
.A2(n_374),
.B1(n_379),
.B2(n_381),
.Y(n_1128)
);

CKINVDCx8_ASAP7_75t_R g1129 ( 
.A(n_911),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_969),
.A2(n_544),
.B(n_529),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_931),
.A2(n_532),
.B(n_538),
.C(n_537),
.Y(n_1131)
);

NOR3xp33_ASAP7_75t_L g1132 ( 
.A(n_956),
.B(n_498),
.C(n_495),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1013),
.Y(n_1133)
);

BUFx2_ASAP7_75t_SL g1134 ( 
.A(n_959),
.Y(n_1134)
);

AO21x2_ASAP7_75t_L g1135 ( 
.A1(n_999),
.A2(n_492),
.B(n_479),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_994),
.B(n_531),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1012),
.A2(n_387),
.B1(n_311),
.B2(n_316),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1065),
.A2(n_381),
.B1(n_542),
.B2(n_523),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_907),
.A2(n_531),
.B(n_542),
.Y(n_1139)
);

BUFx8_ASAP7_75t_L g1140 ( 
.A(n_903),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_994),
.B(n_300),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1065),
.A2(n_546),
.B1(n_542),
.B2(n_523),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_945),
.B(n_973),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_945),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1004),
.A2(n_1067),
.B1(n_1000),
.B2(n_1070),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_910),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_955),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1014),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1038),
.A2(n_1089),
.B(n_1084),
.C(n_1051),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_973),
.B(n_319),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1004),
.B(n_327),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_960),
.B(n_329),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_975),
.B(n_351),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1056),
.A2(n_531),
.B(n_482),
.C(n_484),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1013),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_964),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_968),
.Y(n_1157)
);

AND2x2_ASAP7_75t_SL g1158 ( 
.A(n_922),
.B(n_482),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_1077),
.B(n_356),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1016),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_1046),
.B(n_523),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1057),
.A2(n_360),
.B(n_362),
.C(n_365),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_SL g1163 ( 
.A1(n_1003),
.A2(n_367),
.B1(n_370),
.B2(n_384),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_975),
.B(n_546),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1022),
.Y(n_1165)
);

BUFx8_ASAP7_75t_L g1166 ( 
.A(n_1060),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1023),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_984),
.A2(n_546),
.B1(n_542),
.B2(n_523),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_913),
.A2(n_389),
.B(n_395),
.C(n_492),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_915),
.A2(n_546),
.B1(n_542),
.B2(n_523),
.Y(n_1170)
);

INVx5_ASAP7_75t_L g1171 ( 
.A(n_1013),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_1071),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_980),
.Y(n_1173)
);

OR2x6_ASAP7_75t_L g1174 ( 
.A(n_985),
.B(n_1015),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_1013),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_950),
.A2(n_546),
.B(n_542),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_L g1177 ( 
.A(n_956),
.B(n_484),
.C(n_485),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1028),
.A2(n_485),
.B(n_498),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_922),
.B(n_546),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1055),
.B(n_983),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1024),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_983),
.B(n_495),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_908),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_908),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1034),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_933),
.A2(n_546),
.B1(n_542),
.B2(n_523),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_985),
.B(n_493),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_981),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1018),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1052),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1076),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1071),
.B(n_17),
.Y(n_1192)
);

O2A1O1Ixp5_ASAP7_75t_L g1193 ( 
.A1(n_1069),
.A2(n_493),
.B(n_491),
.C(n_487),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_1015),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1070),
.B(n_1086),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1026),
.A2(n_491),
.B(n_487),
.C(n_542),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_968),
.B(n_523),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1003),
.A2(n_523),
.B1(n_19),
.B2(n_20),
.C(n_21),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_998),
.A2(n_197),
.B(n_195),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_974),
.B(n_17),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_911),
.B(n_20),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1020),
.B(n_25),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1020),
.B(n_25),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1082),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_SL g1205 ( 
.A1(n_1042),
.A2(n_188),
.B(n_185),
.C(n_181),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1026),
.A2(n_26),
.B(n_32),
.C(n_33),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1031),
.B(n_33),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_935),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_933),
.B(n_178),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1041),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1031),
.B(n_34),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_926),
.A2(n_38),
.B(n_40),
.C(n_42),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_950),
.A2(n_138),
.B(n_169),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_R g1214 ( 
.A(n_1041),
.B(n_176),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_935),
.B(n_168),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_927),
.A2(n_126),
.B(n_158),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1066),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1088),
.B(n_38),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1046),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1000),
.B(n_43),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1078),
.B(n_164),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1078),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_941),
.A2(n_156),
.B1(n_150),
.B2(n_147),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_909),
.B(n_129),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_990),
.B(n_45),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_930),
.A2(n_45),
.B(n_46),
.C(n_51),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1053),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_917),
.A2(n_46),
.B(n_51),
.C(n_55),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_919),
.A2(n_87),
.B(n_86),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1062),
.A2(n_55),
.B(n_57),
.C(n_58),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1068),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1058),
.B(n_64),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_948),
.A2(n_89),
.B(n_83),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_947),
.B(n_82),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_949),
.B(n_65),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1087),
.B(n_991),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1005),
.B(n_69),
.Y(n_1237)
);

INVxp33_ASAP7_75t_SL g1238 ( 
.A(n_1048),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1068),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_951),
.A2(n_69),
.B(n_70),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_934),
.A2(n_74),
.B1(n_71),
.B2(n_72),
.Y(n_1241)
);

BUFx10_ASAP7_75t_L g1242 ( 
.A(n_1049),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_952),
.A2(n_70),
.B(n_71),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_977),
.B(n_72),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_977),
.A2(n_73),
.B(n_943),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_953),
.A2(n_957),
.B1(n_1062),
.B2(n_937),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1111),
.A2(n_940),
.B(n_909),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1144),
.B(n_1066),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1191),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1124),
.A2(n_942),
.B(n_978),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1204),
.B(n_1030),
.Y(n_1251)
);

AO21x1_ASAP7_75t_L g1252 ( 
.A1(n_1225),
.A2(n_1036),
.B(n_1072),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1126),
.A2(n_982),
.A3(n_995),
.B(n_1017),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1190),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1239),
.A2(n_1027),
.B1(n_944),
.B2(n_928),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1246),
.A2(n_987),
.A3(n_976),
.B(n_993),
.Y(n_1256)
);

NAND2xp33_ASAP7_75t_SL g1257 ( 
.A(n_1231),
.B(n_923),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1145),
.A2(n_962),
.B(n_972),
.C(n_1032),
.Y(n_1258)
);

NOR2x1_ASAP7_75t_R g1259 ( 
.A(n_1098),
.B(n_943),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1095),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1093),
.A2(n_988),
.B(n_989),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_SL g1262 ( 
.A(n_1090),
.B(n_1027),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1232),
.A2(n_1083),
.B(n_1043),
.C(n_1033),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_SL g1264 ( 
.A(n_1134),
.B(n_1044),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1180),
.B(n_965),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1236),
.A2(n_954),
.B(n_1008),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1149),
.A2(n_1006),
.B(n_996),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1174),
.B(n_965),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1153),
.B(n_1074),
.Y(n_1269)
);

AOI221xp5_ASAP7_75t_SL g1270 ( 
.A1(n_1198),
.A2(n_1025),
.B1(n_1009),
.B2(n_1043),
.C(n_1085),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1158),
.B(n_1045),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_SL g1272 ( 
.A1(n_1149),
.A2(n_1002),
.B(n_1081),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1112),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1219),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1127),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1108),
.B(n_1073),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1238),
.A2(n_1195),
.B1(n_1163),
.B2(n_1220),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1148),
.Y(n_1278)
);

NOR4xp25_ASAP7_75t_L g1279 ( 
.A(n_1230),
.B(n_1019),
.C(n_1021),
.D(n_1037),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1124),
.A2(n_1029),
.A3(n_1035),
.B(n_1050),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1105),
.B(n_1059),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1110),
.A2(n_997),
.B(n_1010),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1143),
.B(n_1080),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1110),
.A2(n_1061),
.B(n_1063),
.Y(n_1284)
);

AOI222xp33_ASAP7_75t_L g1285 ( 
.A1(n_1100),
.A2(n_1075),
.B1(n_1182),
.B2(n_1121),
.C1(n_1137),
.C2(n_1119),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1102),
.B(n_1109),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1113),
.A2(n_1097),
.B1(n_1114),
.B2(n_1157),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1106),
.A2(n_1101),
.B(n_1103),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1174),
.B(n_1210),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1116),
.B(n_1150),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1106),
.A2(n_1103),
.B(n_1164),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1216),
.A2(n_1227),
.B(n_1179),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1216),
.A2(n_1171),
.B(n_1130),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1171),
.A2(n_1233),
.B(n_1229),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1133),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1171),
.A2(n_1233),
.B(n_1229),
.Y(n_1296)
);

AOI221x1_ASAP7_75t_L g1297 ( 
.A1(n_1212),
.A2(n_1243),
.B1(n_1240),
.B2(n_1228),
.C(n_1203),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1096),
.B(n_1094),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1096),
.B(n_1200),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1207),
.B(n_1211),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1171),
.A2(n_1197),
.B(n_1234),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1170),
.A2(n_1122),
.A3(n_1169),
.B(n_1196),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1140),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1240),
.A2(n_1243),
.A3(n_1139),
.B(n_1123),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1123),
.A2(n_1176),
.A3(n_1244),
.B(n_1186),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1131),
.A2(n_1136),
.B(n_1218),
.Y(n_1306)
);

NAND3xp33_ASAP7_75t_L g1307 ( 
.A(n_1128),
.B(n_1177),
.C(n_1132),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1131),
.A2(n_1209),
.B(n_1237),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1241),
.A2(n_1187),
.B1(n_1201),
.B2(n_1099),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1213),
.A2(n_1205),
.B(n_1215),
.Y(n_1310)
);

AOI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1176),
.A2(n_1202),
.B(n_1213),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1199),
.A2(n_1193),
.B(n_1217),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1172),
.B(n_1151),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1192),
.A2(n_1132),
.B1(n_1177),
.B2(n_1235),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1160),
.A2(n_1167),
.B(n_1181),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1157),
.B(n_1185),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_SL g1317 ( 
.A1(n_1206),
.A2(n_1221),
.B(n_1125),
.C(n_1162),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1193),
.A2(n_1165),
.B(n_1168),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1161),
.A2(n_1224),
.B(n_1219),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1194),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1188),
.B(n_1156),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1161),
.A2(n_1224),
.B(n_1222),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1146),
.A2(n_1173),
.B(n_1189),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1147),
.Y(n_1324)
);

BUFx2_ASAP7_75t_R g1325 ( 
.A(n_1107),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1183),
.A2(n_1184),
.B(n_1208),
.Y(n_1326)
);

O2A1O1Ixp33_ASAP7_75t_SL g1327 ( 
.A1(n_1230),
.A2(n_1223),
.B(n_1152),
.C(n_1226),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1208),
.A2(n_1120),
.B(n_1092),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1133),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1141),
.A2(n_1117),
.B1(n_1187),
.B2(n_1242),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1226),
.A2(n_1154),
.B(n_1138),
.C(n_1118),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1135),
.A2(n_1115),
.B(n_1175),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1104),
.A2(n_1154),
.B(n_1142),
.Y(n_1333)
);

OAI22x1_ASAP7_75t_L g1334 ( 
.A1(n_1091),
.A2(n_1175),
.B1(n_1242),
.B2(n_1129),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1133),
.A2(n_1155),
.B(n_1187),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1091),
.A2(n_1174),
.B(n_1155),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1155),
.A2(n_1091),
.B1(n_1159),
.B2(n_1214),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1091),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1140),
.B(n_1166),
.Y(n_1339)
);

OA22x2_ASAP7_75t_L g1340 ( 
.A1(n_1166),
.A2(n_1231),
.B1(n_1239),
.B2(n_580),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1204),
.B(n_742),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1126),
.A2(n_999),
.A3(n_1069),
.B(n_982),
.Y(n_1342)
);

AO32x2_ASAP7_75t_L g1343 ( 
.A1(n_1231),
.A2(n_1137),
.A3(n_1246),
.B1(n_971),
.B2(n_1036),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1204),
.B(n_742),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1102),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1204),
.B(n_742),
.Y(n_1346)
);

AO21x1_ASAP7_75t_L g1347 ( 
.A1(n_1225),
.A2(n_742),
.B(n_906),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_L g1349 ( 
.A1(n_1108),
.A2(n_840),
.B1(n_518),
.B2(n_693),
.C(n_736),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1180),
.B(n_630),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1110),
.A2(n_934),
.B(n_1245),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1153),
.B(n_742),
.C(n_906),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_SL g1353 ( 
.A1(n_1149),
.A2(n_931),
.B(n_1213),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1116),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1093),
.A2(n_742),
.B(n_906),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1180),
.B(n_630),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1180),
.B(n_630),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1124),
.A2(n_1178),
.B(n_1122),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1145),
.A2(n_742),
.B(n_906),
.C(n_797),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1095),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1124),
.A2(n_1178),
.B(n_1122),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1126),
.A2(n_999),
.A3(n_1069),
.B(n_982),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1239),
.A2(n_742),
.B1(n_736),
.B2(n_738),
.Y(n_1366)
);

INVx4_ASAP7_75t_L g1367 ( 
.A(n_1171),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1239),
.A2(n_742),
.B1(n_736),
.B2(n_738),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1191),
.Y(n_1369)
);

AO21x1_ASAP7_75t_L g1370 ( 
.A1(n_1225),
.A2(n_742),
.B(n_906),
.Y(n_1370)
);

OAI22x1_ASAP7_75t_L g1371 ( 
.A1(n_1239),
.A2(n_1145),
.B1(n_1232),
.B2(n_693),
.Y(n_1371)
);

BUFx8_ASAP7_75t_L g1372 ( 
.A(n_1210),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1373)
);

O2A1O1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1232),
.A2(n_742),
.B(n_906),
.C(n_736),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1232),
.A2(n_742),
.B(n_906),
.C(n_736),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1180),
.B(n_1174),
.Y(n_1376)
);

AO31x2_ASAP7_75t_L g1377 ( 
.A1(n_1126),
.A2(n_999),
.A3(n_1069),
.B(n_982),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1239),
.B(n_742),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1095),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1116),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1158),
.B(n_631),
.Y(n_1381)
);

BUFx10_ASAP7_75t_L g1382 ( 
.A(n_1150),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1204),
.B(n_742),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1090),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1145),
.A2(n_742),
.B(n_906),
.C(n_797),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_SL g1387 ( 
.A(n_1090),
.B(n_631),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1239),
.B(n_742),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1204),
.B(n_742),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1116),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1239),
.A2(n_742),
.B1(n_1231),
.B2(n_1232),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1095),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1239),
.A2(n_742),
.B1(n_1231),
.B2(n_1232),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1158),
.B(n_631),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1239),
.A2(n_742),
.B1(n_736),
.B2(n_738),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1145),
.A2(n_742),
.B(n_906),
.C(n_797),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1095),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1111),
.A2(n_742),
.B(n_659),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1095),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1180),
.B(n_630),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1126),
.A2(n_999),
.A3(n_1069),
.B(n_982),
.Y(n_1406)
);

AO21x1_ASAP7_75t_L g1407 ( 
.A1(n_1225),
.A2(n_742),
.B(n_906),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1194),
.Y(n_1408)
);

CKINVDCx11_ASAP7_75t_R g1409 ( 
.A(n_1320),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1340),
.A2(n_1389),
.B1(n_1378),
.B2(n_1368),
.Y(n_1410)
);

BUFx8_ASAP7_75t_L g1411 ( 
.A(n_1408),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1366),
.A2(n_1399),
.B1(n_1349),
.B2(n_1371),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1384),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1300),
.B(n_1360),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1307),
.A2(n_1352),
.B1(n_1397),
.B2(n_1393),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1307),
.A2(n_1352),
.B1(n_1290),
.B2(n_1382),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1260),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1314),
.B2(n_1277),
.Y(n_1418)
);

CKINVDCx11_ASAP7_75t_R g1419 ( 
.A(n_1345),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1374),
.B(n_1375),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1277),
.A2(n_1314),
.B1(n_1344),
.B2(n_1341),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1346),
.A2(n_1391),
.B1(n_1383),
.B2(n_1385),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1273),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1249),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1286),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1330),
.A2(n_1387),
.B1(n_1262),
.B2(n_1271),
.Y(n_1426)
);

INVx6_ASAP7_75t_L g1427 ( 
.A(n_1372),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1372),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1354),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1309),
.A2(n_1285),
.B1(n_1299),
.B2(n_1298),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1382),
.A2(n_1271),
.B1(n_1337),
.B2(n_1355),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1381),
.B(n_1398),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1350),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1288),
.A2(n_1283),
.B1(n_1353),
.B2(n_1343),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1376),
.B(n_1289),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1295),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1281),
.A2(n_1257),
.B1(n_1265),
.B2(n_1330),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1369),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1265),
.A2(n_1287),
.B1(n_1308),
.B2(n_1376),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1275),
.Y(n_1440)
);

INVx6_ASAP7_75t_L g1441 ( 
.A(n_1367),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1401),
.A2(n_1251),
.B1(n_1396),
.B2(n_1361),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1357),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1254),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1324),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1278),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1379),
.A2(n_1402),
.B1(n_1404),
.B2(n_1269),
.Y(n_1447)
);

OAI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1276),
.A2(n_1297),
.B1(n_1248),
.B2(n_1392),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1313),
.A2(n_1380),
.B1(n_1268),
.B2(n_1407),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1316),
.A2(n_1331),
.B1(n_1289),
.B2(n_1321),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1358),
.B(n_1405),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1268),
.A2(n_1264),
.B1(n_1255),
.B2(n_1327),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1315),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1318),
.A2(n_1258),
.B1(n_1338),
.B2(n_1306),
.Y(n_1454)
);

BUFx2_ASAP7_75t_SL g1455 ( 
.A(n_1303),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1325),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1318),
.A2(n_1261),
.B1(n_1335),
.B2(n_1343),
.Y(n_1457)
);

CKINVDCx11_ASAP7_75t_R g1458 ( 
.A(n_1295),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1347),
.A2(n_1370),
.B1(n_1334),
.B2(n_1252),
.Y(n_1459)
);

INVx8_ASAP7_75t_L g1460 ( 
.A(n_1329),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1343),
.A2(n_1292),
.B1(n_1310),
.B2(n_1291),
.Y(n_1461)
);

INVx6_ASAP7_75t_L g1462 ( 
.A(n_1329),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1329),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1328),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1339),
.Y(n_1465)
);

NAND2x1p5_ASAP7_75t_L g1466 ( 
.A(n_1274),
.B(n_1326),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1323),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1259),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1274),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1348),
.B(n_1394),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1336),
.A2(n_1296),
.B1(n_1294),
.B2(n_1247),
.Y(n_1471)
);

BUFx12f_ASAP7_75t_L g1472 ( 
.A(n_1317),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1263),
.A2(n_1364),
.B(n_1403),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1356),
.A2(n_1386),
.B1(n_1400),
.B2(n_1395),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1333),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1365),
.A2(n_1390),
.B1(n_1388),
.B2(n_1373),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1311),
.A2(n_1293),
.B(n_1301),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1304),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1304),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1266),
.B(n_1279),
.Y(n_1480)
);

BUFx12f_ASAP7_75t_L g1481 ( 
.A(n_1272),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1279),
.B(n_1267),
.Y(n_1482)
);

INVx6_ASAP7_75t_L g1483 ( 
.A(n_1319),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1305),
.B(n_1406),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1332),
.A2(n_1250),
.B(n_1270),
.Y(n_1485)
);

INVx5_ASAP7_75t_L g1486 ( 
.A(n_1322),
.Y(n_1486)
);

INVx6_ASAP7_75t_L g1487 ( 
.A(n_1351),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1312),
.A2(n_1282),
.B1(n_1362),
.B2(n_1359),
.Y(n_1488)
);

BUFx2_ASAP7_75t_SL g1489 ( 
.A(n_1284),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1270),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1305),
.A2(n_1302),
.B1(n_1406),
.B2(n_1342),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1256),
.Y(n_1492)
);

OAI21xp33_ASAP7_75t_L g1493 ( 
.A1(n_1363),
.A2(n_1377),
.B(n_1302),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1363),
.A2(n_1377),
.B1(n_1253),
.B2(n_1256),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1377),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1256),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1253),
.A2(n_1371),
.B1(n_742),
.B2(n_1349),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1253),
.A2(n_1393),
.B1(n_1397),
.B2(n_1239),
.Y(n_1498)
);

INVx11_ASAP7_75t_L g1499 ( 
.A(n_1280),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1280),
.A2(n_1371),
.B1(n_742),
.B2(n_1349),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1280),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1300),
.B(n_1360),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1239),
.B2(n_742),
.Y(n_1503)
);

BUFx12f_ASAP7_75t_L g1504 ( 
.A(n_1320),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1345),
.Y(n_1505)
);

CKINVDCx11_ASAP7_75t_R g1506 ( 
.A(n_1320),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1239),
.B2(n_742),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1340),
.A2(n_1239),
.B1(n_1231),
.B2(n_742),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1340),
.A2(n_1239),
.B1(n_1231),
.B2(n_742),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1295),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1345),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1260),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1260),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1516)
);

OAI22x1_ASAP7_75t_L g1517 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1277),
.B2(n_1314),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1260),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1393),
.A2(n_742),
.B1(n_1397),
.B2(n_1239),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1372),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1286),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1286),
.Y(n_1522)
);

INVx8_ASAP7_75t_L g1523 ( 
.A(n_1295),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1260),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1340),
.A2(n_1239),
.B1(n_1231),
.B2(n_742),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1239),
.B2(n_742),
.Y(n_1529)
);

CKINVDCx11_ASAP7_75t_R g1530 ( 
.A(n_1320),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1239),
.B2(n_742),
.Y(n_1532)
);

AO22x1_ASAP7_75t_L g1533 ( 
.A1(n_1378),
.A2(n_742),
.B1(n_693),
.B2(n_939),
.Y(n_1533)
);

INVx4_ASAP7_75t_R g1534 ( 
.A(n_1345),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1286),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1260),
.Y(n_1536)
);

INVx8_ASAP7_75t_L g1537 ( 
.A(n_1295),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1300),
.B(n_1360),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1300),
.B(n_1360),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1367),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1239),
.B2(n_742),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1260),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1372),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1260),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1239),
.B2(n_742),
.Y(n_1546)
);

INVx6_ASAP7_75t_L g1547 ( 
.A(n_1372),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1300),
.B(n_1360),
.Y(n_1548)
);

INVx6_ASAP7_75t_L g1549 ( 
.A(n_1372),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1371),
.A2(n_742),
.B1(n_1349),
.B2(n_1366),
.Y(n_1550)
);

CKINVDCx16_ASAP7_75t_R g1551 ( 
.A(n_1387),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1372),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1260),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1393),
.A2(n_1397),
.B1(n_1239),
.B2(n_742),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1384),
.Y(n_1555)
);

BUFx12f_ASAP7_75t_L g1556 ( 
.A(n_1320),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1260),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1453),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1481),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1434),
.B(n_1484),
.Y(n_1560)
);

AOI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1420),
.A2(n_1482),
.B(n_1470),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1517),
.A2(n_1418),
.B1(n_1415),
.B2(n_1430),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1478),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1521),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1451),
.B(n_1433),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1479),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1447),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1503),
.A2(n_1529),
.B1(n_1554),
.B2(n_1532),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1522),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1446),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1473),
.A2(n_1485),
.B(n_1480),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1421),
.B(n_1422),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1495),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1434),
.B(n_1500),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1555),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1483),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1501),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1475),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1447),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1483),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1493),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1470),
.A2(n_1476),
.B(n_1474),
.Y(n_1582)
);

AO31x2_ASAP7_75t_L g1583 ( 
.A1(n_1461),
.A2(n_1454),
.A3(n_1491),
.B(n_1457),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1491),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1496),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_SL g1586 ( 
.A(n_1472),
.B(n_1442),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1425),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1456),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1499),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1487),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1492),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1487),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1454),
.Y(n_1593)
);

AO32x2_ASAP7_75t_L g1594 ( 
.A1(n_1457),
.A2(n_1498),
.A3(n_1461),
.B1(n_1492),
.B2(n_1503),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1486),
.B(n_1464),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1509),
.A2(n_1510),
.B1(n_1527),
.B2(n_1410),
.Y(n_1596)
);

AO21x2_ASAP7_75t_L g1597 ( 
.A1(n_1485),
.A2(n_1477),
.B(n_1502),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1508),
.A2(n_1546),
.B1(n_1529),
.B2(n_1554),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1459),
.B(n_1497),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1535),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1423),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1440),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1443),
.Y(n_1603)
);

INVx11_ASAP7_75t_L g1604 ( 
.A(n_1411),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1442),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1467),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1486),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1422),
.B(n_1533),
.Y(n_1608)
);

AO21x1_ASAP7_75t_SL g1609 ( 
.A1(n_1414),
.A2(n_1548),
.B(n_1502),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1416),
.B(n_1429),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1508),
.A2(n_1546),
.B1(n_1541),
.B2(n_1532),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1494),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1498),
.B(n_1490),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1414),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1538),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1538),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1412),
.B(n_1410),
.Y(n_1617)
);

OAI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1466),
.A2(n_1548),
.B(n_1539),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1448),
.B(n_1539),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1486),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1514),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1439),
.A2(n_1450),
.B(n_1452),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1551),
.B(n_1519),
.Y(n_1623)
);

AO21x1_ASAP7_75t_L g1624 ( 
.A1(n_1541),
.A2(n_1426),
.B(n_1450),
.Y(n_1624)
);

AND2x4_ASAP7_75t_SL g1625 ( 
.A(n_1437),
.B(n_1435),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1515),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1507),
.A2(n_1512),
.B1(n_1516),
.B2(n_1550),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1469),
.A2(n_1488),
.B(n_1553),
.Y(n_1628)
);

AO21x2_ASAP7_75t_L g1629 ( 
.A1(n_1518),
.A2(n_1557),
.B(n_1545),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1536),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1417),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1525),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1542),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1489),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1424),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_SL g1636 ( 
.A1(n_1520),
.A2(n_1552),
.B(n_1432),
.C(n_1540),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1438),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1435),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1471),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1444),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1445),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1524),
.B(n_1526),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1431),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1449),
.Y(n_1644)
);

INVx6_ASAP7_75t_L g1645 ( 
.A(n_1463),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1528),
.B(n_1531),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1544),
.B(n_1509),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1510),
.B(n_1527),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1441),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1465),
.B(n_1505),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1462),
.A2(n_1523),
.B(n_1537),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1436),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1458),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1511),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1513),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1462),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1460),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1537),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1427),
.Y(n_1659)
);

OAI222xp33_ASAP7_75t_L g1660 ( 
.A1(n_1428),
.A2(n_1468),
.B1(n_1534),
.B2(n_1549),
.C1(n_1547),
.C2(n_1427),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1455),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1419),
.A2(n_1549),
.B(n_1547),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1427),
.A2(n_1549),
.B(n_1547),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1543),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1543),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1543),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1411),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1613),
.B(n_1413),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1613),
.B(n_1504),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1570),
.B(n_1556),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1559),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1589),
.B(n_1409),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1560),
.B(n_1506),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1560),
.B(n_1530),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1596),
.A2(n_1617),
.B1(n_1572),
.B2(n_1627),
.C(n_1562),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1601),
.Y(n_1676)
);

NOR2x1_ASAP7_75t_SL g1677 ( 
.A(n_1609),
.B(n_1619),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_SL g1678 ( 
.A(n_1609),
.B(n_1619),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1617),
.B(n_1608),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1564),
.B(n_1587),
.Y(n_1680)
);

O2A1O1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1642),
.A2(n_1646),
.B(n_1648),
.C(n_1624),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1586),
.A2(n_1582),
.B(n_1620),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1594),
.B(n_1571),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1614),
.B(n_1615),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1568),
.B(n_1598),
.C(n_1611),
.D(n_1647),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1594),
.B(n_1571),
.Y(n_1687)
);

NOR2x1_ASAP7_75t_SL g1688 ( 
.A(n_1634),
.B(n_1597),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1622),
.A2(n_1647),
.B(n_1610),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1643),
.A2(n_1644),
.B1(n_1661),
.B2(n_1569),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1594),
.B(n_1571),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1624),
.A2(n_1574),
.B1(n_1599),
.B2(n_1644),
.C(n_1567),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1580),
.B(n_1663),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1614),
.B(n_1615),
.Y(n_1694)
);

OAI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1579),
.A2(n_1599),
.B(n_1605),
.C(n_1639),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1622),
.A2(n_1639),
.B(n_1605),
.C(n_1593),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1616),
.B(n_1631),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1663),
.B(n_1576),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1593),
.A2(n_1616),
.B(n_1625),
.C(n_1618),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1625),
.A2(n_1618),
.B(n_1594),
.C(n_1581),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1636),
.A2(n_1660),
.B(n_1661),
.C(n_1600),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1633),
.B(n_1635),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1655),
.A2(n_1625),
.B1(n_1664),
.B2(n_1603),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1602),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1629),
.Y(n_1705)
);

OAI211xp5_ASAP7_75t_SL g1706 ( 
.A1(n_1662),
.A2(n_1650),
.B(n_1667),
.C(n_1565),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1594),
.B(n_1612),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1597),
.A2(n_1586),
.B(n_1634),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1612),
.A2(n_1584),
.B1(n_1597),
.B2(n_1606),
.C(n_1621),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1654),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1590),
.B(n_1607),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1583),
.B(n_1602),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1559),
.B(n_1561),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1559),
.A2(n_1584),
.B(n_1659),
.C(n_1664),
.Y(n_1714)
);

INVxp33_ASAP7_75t_SL g1715 ( 
.A(n_1588),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1664),
.A2(n_1667),
.B1(n_1659),
.B2(n_1666),
.Y(n_1716)
);

BUFx4f_ASAP7_75t_SL g1717 ( 
.A(n_1653),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1651),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1637),
.B(n_1640),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1558),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1628),
.A2(n_1591),
.B(n_1595),
.Y(n_1721)
);

AO21x2_ASAP7_75t_L g1722 ( 
.A1(n_1628),
.A2(n_1577),
.B(n_1578),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1575),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1656),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1656),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1626),
.B(n_1630),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1583),
.B(n_1578),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1632),
.B(n_1641),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1651),
.Y(n_1729)
);

O2A1O1Ixp33_ASAP7_75t_L g1730 ( 
.A1(n_1665),
.A2(n_1666),
.B(n_1659),
.C(n_1649),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1683),
.B(n_1583),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1698),
.B(n_1595),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1712),
.B(n_1583),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1683),
.B(n_1583),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1687),
.B(n_1585),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1720),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1729),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1712),
.B(n_1707),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1687),
.B(n_1566),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1718),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1705),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1722),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1718),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1595),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1707),
.B(n_1629),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1691),
.B(n_1573),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1727),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1700),
.B(n_1563),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1688),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1675),
.A2(n_1659),
.B1(n_1638),
.B2(n_1645),
.Y(n_1750)
);

OAI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1681),
.A2(n_1592),
.B(n_1591),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1676),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1704),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1726),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1728),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1682),
.Y(n_1756)
);

OAI211xp5_ASAP7_75t_L g1757 ( 
.A1(n_1751),
.A2(n_1692),
.B(n_1686),
.C(n_1689),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1745),
.B(n_1709),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1753),
.Y(n_1759)
);

AOI31xp33_ASAP7_75t_L g1760 ( 
.A1(n_1751),
.A2(n_1673),
.A3(n_1674),
.B(n_1672),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1753),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1736),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1753),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1751),
.A2(n_1678),
.B1(n_1677),
.B2(n_1695),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1750),
.A2(n_1706),
.B1(n_1685),
.B2(n_1679),
.Y(n_1765)
);

INVx4_ASAP7_75t_L g1766 ( 
.A(n_1743),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_L g1767 ( 
.A(n_1750),
.B(n_1685),
.C(n_1679),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1752),
.Y(n_1768)
);

AOI211xp5_ASAP7_75t_L g1769 ( 
.A1(n_1748),
.A2(n_1701),
.B(n_1690),
.C(n_1674),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1732),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1745),
.B(n_1696),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1734),
.A2(n_1716),
.B1(n_1703),
.B2(n_1671),
.Y(n_1772)
);

INVxp67_ASAP7_75t_SL g1773 ( 
.A(n_1741),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1737),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1745),
.B(n_1754),
.Y(n_1775)
);

AO21x2_ASAP7_75t_L g1776 ( 
.A1(n_1742),
.A2(n_1708),
.B(n_1721),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1747),
.B(n_1680),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1752),
.Y(n_1778)
);

AOI222xp33_ASAP7_75t_L g1779 ( 
.A1(n_1750),
.A2(n_1673),
.B1(n_1672),
.B2(n_1717),
.C1(n_1669),
.C2(n_1668),
.Y(n_1779)
);

BUFx3_ASAP7_75t_L g1780 ( 
.A(n_1737),
.Y(n_1780)
);

OAI31xp33_ASAP7_75t_L g1781 ( 
.A1(n_1748),
.A2(n_1714),
.A3(n_1699),
.B(n_1696),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1736),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1747),
.B(n_1711),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1747),
.B(n_1711),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1735),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1747),
.B(n_1739),
.Y(n_1786)
);

OAI33xp33_ASAP7_75t_L g1787 ( 
.A1(n_1733),
.A2(n_1702),
.A3(n_1719),
.B1(n_1697),
.B2(n_1684),
.B3(n_1694),
.Y(n_1787)
);

OAI33xp33_ASAP7_75t_L g1788 ( 
.A1(n_1733),
.A2(n_1710),
.A3(n_1725),
.B1(n_1724),
.B2(n_1730),
.B3(n_1652),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1754),
.B(n_1713),
.Y(n_1789)
);

OAI211xp5_ASAP7_75t_L g1790 ( 
.A1(n_1733),
.A2(n_1699),
.B(n_1713),
.C(n_1714),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1740),
.B(n_1693),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1732),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1770),
.B(n_1731),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1771),
.B(n_1734),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1758),
.B(n_1731),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1792),
.B(n_1732),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1758),
.B(n_1731),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1759),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1792),
.B(n_1732),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1759),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1786),
.B(n_1732),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_SL g1802 ( 
.A(n_1774),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1774),
.B(n_1744),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1761),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1771),
.B(n_1738),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1762),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1786),
.B(n_1744),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1761),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1775),
.B(n_1738),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1791),
.B(n_1744),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1791),
.B(n_1744),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1763),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1774),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1789),
.B(n_1754),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1791),
.B(n_1744),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1767),
.B(n_1715),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1763),
.Y(n_1817)
);

CKINVDCx16_ASAP7_75t_R g1818 ( 
.A(n_1780),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1762),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1780),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_R g1821 ( 
.A(n_1765),
.B(n_1723),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1775),
.B(n_1738),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1780),
.B(n_1744),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1762),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1789),
.B(n_1746),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1773),
.B(n_1755),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1767),
.B(n_1715),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1777),
.B(n_1746),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1798),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1802),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1793),
.B(n_1785),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1802),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1793),
.B(n_1783),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1806),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1801),
.B(n_1784),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1806),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1798),
.Y(n_1837)
);

OAI21xp33_ASAP7_75t_L g1838 ( 
.A1(n_1821),
.A2(n_1757),
.B(n_1764),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1800),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1800),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1813),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1794),
.B(n_1782),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1795),
.B(n_1768),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1816),
.B(n_1757),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1804),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1795),
.B(n_1768),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1796),
.B(n_1803),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1794),
.B(n_1782),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1806),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1804),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1819),
.Y(n_1851)
);

INVxp33_ASAP7_75t_L g1852 ( 
.A(n_1827),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1819),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1819),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1807),
.B(n_1791),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1797),
.B(n_1778),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1805),
.B(n_1782),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1824),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1824),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1824),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1805),
.B(n_1787),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1796),
.B(n_1766),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1813),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1808),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1797),
.B(n_1778),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1809),
.B(n_1822),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1820),
.Y(n_1867)
);

NOR2xp67_ASAP7_75t_L g1868 ( 
.A(n_1803),
.B(n_1790),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1796),
.B(n_1799),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1796),
.B(n_1799),
.Y(n_1870)
);

OAI21xp33_ASAP7_75t_L g1871 ( 
.A1(n_1838),
.A2(n_1769),
.B(n_1760),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1866),
.B(n_1814),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1844),
.B(n_1814),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1844),
.B(n_1769),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1863),
.Y(n_1875)
);

AND4x1_ASAP7_75t_L g1876 ( 
.A(n_1838),
.B(n_1779),
.C(n_1781),
.D(n_1788),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1863),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1850),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1850),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1863),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1861),
.B(n_1818),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1861),
.B(n_1818),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1830),
.B(n_1810),
.Y(n_1883)
);

OAI211xp5_ASAP7_75t_SL g1884 ( 
.A1(n_1830),
.A2(n_1779),
.B(n_1781),
.C(n_1790),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1832),
.B(n_1826),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1841),
.Y(n_1886)
);

INVxp67_ASAP7_75t_L g1887 ( 
.A(n_1832),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1852),
.B(n_1604),
.Y(n_1888)
);

NAND2x1p5_ASAP7_75t_L g1889 ( 
.A(n_1868),
.B(n_1820),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1834),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1866),
.B(n_1809),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1829),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1866),
.B(n_1822),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1829),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1868),
.B(n_1810),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1867),
.B(n_1820),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1841),
.B(n_1825),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1829),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1834),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1837),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1847),
.B(n_1811),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1837),
.Y(n_1902)
);

CKINVDCx16_ASAP7_75t_R g1903 ( 
.A(n_1867),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_SL g1904 ( 
.A(n_1867),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1857),
.B(n_1825),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1847),
.B(n_1811),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1852),
.B(n_1833),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1837),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1874),
.A2(n_1760),
.B1(n_1772),
.B2(n_1737),
.Y(n_1909)
);

INVxp67_ASAP7_75t_L g1910 ( 
.A(n_1904),
.Y(n_1910)
);

CKINVDCx16_ASAP7_75t_R g1911 ( 
.A(n_1903),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1883),
.B(n_1815),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1896),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1871),
.A2(n_1672),
.B(n_1670),
.Y(n_1914)
);

OR2x6_ASAP7_75t_L g1915 ( 
.A(n_1887),
.B(n_1645),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1877),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1877),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1881),
.A2(n_1828),
.B1(n_1671),
.B2(n_1749),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1883),
.B(n_1815),
.Y(n_1919)
);

OAI21xp33_ASAP7_75t_L g1920 ( 
.A1(n_1882),
.A2(n_1846),
.B(n_1843),
.Y(n_1920)
);

OAI22x1_ASAP7_75t_L g1921 ( 
.A1(n_1876),
.A2(n_1847),
.B1(n_1803),
.B2(n_1823),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1884),
.A2(n_1840),
.B1(n_1845),
.B2(n_1839),
.C(n_1864),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1888),
.B(n_1604),
.Y(n_1923)
);

OAI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1889),
.A2(n_1847),
.B1(n_1823),
.B2(n_1803),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1889),
.B(n_1847),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1875),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1888),
.A2(n_1823),
.B1(n_1847),
.B2(n_1831),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1901),
.Y(n_1928)
);

OAI32xp33_ASAP7_75t_L g1929 ( 
.A1(n_1889),
.A2(n_1857),
.A3(n_1842),
.B1(n_1848),
.B2(n_1831),
.Y(n_1929)
);

OAI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1873),
.A2(n_1828),
.B1(n_1671),
.B2(n_1749),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1907),
.A2(n_1895),
.B1(n_1885),
.B2(n_1886),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1875),
.Y(n_1932)
);

O2A1O1Ixp33_ASAP7_75t_L g1933 ( 
.A1(n_1880),
.A2(n_1864),
.B(n_1839),
.C(n_1840),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1895),
.A2(n_1823),
.B1(n_1831),
.B2(n_1862),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1892),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1911),
.A2(n_1896),
.B1(n_1901),
.B2(n_1906),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1926),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1932),
.Y(n_1938)
);

OAI31xp33_ASAP7_75t_L g1939 ( 
.A1(n_1909),
.A2(n_1896),
.A3(n_1897),
.B(n_1879),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1931),
.B(n_1897),
.Y(n_1940)
);

OAI21xp33_ASAP7_75t_L g1941 ( 
.A1(n_1921),
.A2(n_1878),
.B(n_1891),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1913),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1935),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1910),
.A2(n_1898),
.B(n_1894),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1925),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1916),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1917),
.B(n_1891),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1909),
.A2(n_1906),
.B1(n_1893),
.B2(n_1776),
.Y(n_1948)
);

OAI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1914),
.A2(n_1893),
.B(n_1872),
.Y(n_1949)
);

O2A1O1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1929),
.A2(n_1908),
.B(n_1900),
.C(n_1902),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1933),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1914),
.B(n_1872),
.Y(n_1952)
);

INVxp67_ASAP7_75t_L g1953 ( 
.A(n_1915),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1928),
.A2(n_1776),
.B1(n_1862),
.B2(n_1749),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1927),
.A2(n_1862),
.B(n_1905),
.Y(n_1955)
);

INVxp67_ASAP7_75t_SL g1956 ( 
.A(n_1924),
.Y(n_1956)
);

OAI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1922),
.A2(n_1905),
.B1(n_1756),
.B2(n_1839),
.C(n_1864),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1947),
.Y(n_1958)
);

NOR2x1_ASAP7_75t_L g1959 ( 
.A(n_1951),
.B(n_1915),
.Y(n_1959)
);

A2O1A1Ixp33_ASAP7_75t_SL g1960 ( 
.A1(n_1953),
.A2(n_1939),
.B(n_1957),
.C(n_1946),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1937),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1938),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1942),
.B(n_1915),
.Y(n_1963)
);

NAND3xp33_ASAP7_75t_L g1964 ( 
.A(n_1940),
.B(n_1920),
.C(n_1934),
.Y(n_1964)
);

AO22x2_ASAP7_75t_L g1965 ( 
.A1(n_1944),
.A2(n_1890),
.B1(n_1899),
.B2(n_1845),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1936),
.B(n_1923),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_SL g1967 ( 
.A1(n_1949),
.A2(n_1919),
.B1(n_1912),
.B2(n_1776),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1945),
.B(n_1855),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1956),
.A2(n_1918),
.B1(n_1930),
.B2(n_1776),
.Y(n_1969)
);

NAND3xp33_ASAP7_75t_L g1970 ( 
.A(n_1960),
.B(n_1964),
.C(n_1959),
.Y(n_1970)
);

NAND4xp25_ASAP7_75t_L g1971 ( 
.A(n_1966),
.B(n_1941),
.C(n_1944),
.D(n_1948),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1963),
.B(n_1952),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1968),
.B(n_1955),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1958),
.B(n_1943),
.Y(n_1974)
);

OAI211xp5_ASAP7_75t_L g1975 ( 
.A1(n_1967),
.A2(n_1957),
.B(n_1950),
.C(n_1954),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1965),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1961),
.B(n_1835),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1969),
.B(n_1840),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1962),
.B(n_1835),
.Y(n_1979)
);

AOI211xp5_ASAP7_75t_L g1980 ( 
.A1(n_1970),
.A2(n_1965),
.B(n_1899),
.C(n_1890),
.Y(n_1980)
);

AOI211xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1975),
.A2(n_1723),
.B(n_1845),
.C(n_1857),
.Y(n_1981)
);

AOI211xp5_ASAP7_75t_L g1982 ( 
.A1(n_1971),
.A2(n_1836),
.B(n_1834),
.C(n_1849),
.Y(n_1982)
);

NOR2x1_ASAP7_75t_L g1983 ( 
.A(n_1976),
.B(n_1834),
.Y(n_1983)
);

OAI21xp33_ASAP7_75t_L g1984 ( 
.A1(n_1972),
.A2(n_1849),
.B(n_1836),
.Y(n_1984)
);

AOI211xp5_ASAP7_75t_SL g1985 ( 
.A1(n_1974),
.A2(n_1848),
.B(n_1842),
.C(n_1836),
.Y(n_1985)
);

NAND4xp75_ASAP7_75t_L g1986 ( 
.A(n_1983),
.B(n_1973),
.C(n_1978),
.D(n_1979),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1980),
.A2(n_1977),
.B1(n_1848),
.B2(n_1842),
.Y(n_1987)
);

OAI211xp5_ASAP7_75t_L g1988 ( 
.A1(n_1981),
.A2(n_1836),
.B(n_1860),
.C(n_1849),
.Y(n_1988)
);

AOI21xp33_ASAP7_75t_L g1989 ( 
.A1(n_1984),
.A2(n_1851),
.B(n_1849),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1982),
.A2(n_1858),
.B1(n_1853),
.B2(n_1851),
.C(n_1860),
.Y(n_1990)
);

O2A1O1Ixp33_ASAP7_75t_L g1991 ( 
.A1(n_1985),
.A2(n_1854),
.B(n_1859),
.C(n_1858),
.Y(n_1991)
);

BUFx2_ASAP7_75t_L g1992 ( 
.A(n_1983),
.Y(n_1992)
);

NAND5xp2_ASAP7_75t_L g1993 ( 
.A(n_1988),
.B(n_1870),
.C(n_1869),
.D(n_1855),
.E(n_1645),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1992),
.Y(n_1994)
);

NAND2xp33_ASAP7_75t_SL g1995 ( 
.A(n_1987),
.B(n_1855),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1986),
.B(n_1843),
.Y(n_1996)
);

NAND2x1p5_ASAP7_75t_L g1997 ( 
.A(n_1989),
.B(n_1658),
.Y(n_1997)
);

NOR2xp67_ASAP7_75t_L g1998 ( 
.A(n_1991),
.B(n_1851),
.Y(n_1998)
);

OAI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1996),
.A2(n_1990),
.B1(n_1853),
.B2(n_1854),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1994),
.Y(n_2000)
);

NOR2x1p5_ASAP7_75t_L g2001 ( 
.A(n_1993),
.B(n_1851),
.Y(n_2001)
);

NAND3xp33_ASAP7_75t_L g2002 ( 
.A(n_1995),
.B(n_1854),
.C(n_1853),
.Y(n_2002)
);

O2A1O1Ixp33_ASAP7_75t_L g2003 ( 
.A1(n_2000),
.A2(n_1997),
.B(n_1998),
.C(n_1854),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_2003),
.Y(n_2004)
);

OR3x1_ASAP7_75t_L g2005 ( 
.A(n_2004),
.B(n_2001),
.C(n_1999),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_2004),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_2005),
.A2(n_2002),
.B1(n_1853),
.B2(n_1858),
.Y(n_2007)
);

AOI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_2006),
.A2(n_1858),
.B1(n_1860),
.B2(n_1859),
.Y(n_2008)
);

OAI21xp33_ASAP7_75t_L g2009 ( 
.A1(n_2008),
.A2(n_1860),
.B(n_1859),
.Y(n_2009)
);

XNOR2xp5_ASAP7_75t_L g2010 ( 
.A(n_2007),
.B(n_1869),
.Y(n_2010)
);

OAI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_2010),
.A2(n_1859),
.B(n_1856),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_2011),
.B(n_2009),
.Y(n_2012)
);

OAI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_2012),
.A2(n_1645),
.B1(n_1846),
.B2(n_1865),
.Y(n_2013)
);

OAI221xp5_ASAP7_75t_R g2014 ( 
.A1(n_2013),
.A2(n_1865),
.B1(n_1856),
.B2(n_1808),
.C(n_1812),
.Y(n_2014)
);

AOI211xp5_ASAP7_75t_L g2015 ( 
.A1(n_2014),
.A2(n_1658),
.B(n_1657),
.C(n_1817),
.Y(n_2015)
);


endmodule