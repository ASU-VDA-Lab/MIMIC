module real_jpeg_20822_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_314, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_314;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_51),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_20),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_1),
.B(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_71),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_1),
.A2(n_10),
.B(n_45),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_1),
.B(n_54),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_1),
.A2(n_24),
.B(n_56),
.C(n_204),
.Y(n_203)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_3),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_3),
.A2(n_22),
.B1(n_45),
.B2(n_46),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_3),
.A2(n_22),
.B1(n_39),
.B2(n_40),
.Y(n_246)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_4),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_4),
.B(n_154),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_6),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_119),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_119),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_119),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_20),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_9),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_9),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_10),
.A2(n_39),
.B(n_43),
.C(n_44),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_10),
.B(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_11),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_97),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_95),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_82),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_15),
.B(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_69),
.C(n_77),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_16),
.A2(n_17),
.B1(n_69),
.B2(n_300),
.Y(n_306)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_34),
.B1(n_35),
.B2(n_68),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_23),
.B(n_27),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_19),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_23),
.B(n_30),
.C(n_31),
.Y(n_29)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_23),
.B(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_23),
.A2(n_29),
.B(n_75),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_24),
.A2(n_55),
.B(n_56),
.C(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_24),
.B(n_26),
.Y(n_140)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_25),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_28),
.B(n_117),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_29),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_31),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_36),
.B(n_67),
.C(n_68),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_36),
.A2(n_66),
.B1(n_120),
.B2(n_121),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_36),
.A2(n_66),
.B1(n_78),
.B2(n_303),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_48),
.B(n_49),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_37),
.A2(n_112),
.B(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_38),
.B(n_50),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_38),
.B(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_38),
.B(n_113),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_40),
.B1(n_56),
.B2(n_58),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_39),
.A2(n_51),
.B(n_58),
.Y(n_204)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_40),
.A2(n_47),
.B(n_51),
.C(n_169),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_44),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_44),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_44),
.B(n_50),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_46),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_48),
.B(n_51),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_48),
.A2(n_209),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_51),
.B(n_107),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_60),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_53),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_54),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_65),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_62),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_55),
.A2(n_60),
.B(n_80),
.Y(n_283)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_59),
.B(n_61),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_79),
.B(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_62),
.B(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_69),
.C(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_116),
.C(n_120),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_69),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_69),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_71),
.B(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_75),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_77),
.B(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_78),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_81),
.B(n_131),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_81),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_91),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_86),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_89),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_89),
.A2(n_91),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_91),
.B(n_248),
.C(n_251),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_297),
.A3(n_307),
.B1(n_310),
.B2(n_311),
.C(n_314),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_276),
.B(n_296),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_255),
.B(n_275),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_156),
.B(n_238),
.C(n_254),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_143),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_102),
.B(n_143),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_124),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_104),
.B(n_115),
.C(n_124),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_111),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_105),
.B(n_111),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_106),
.A2(n_107),
.B(n_155),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_108),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_112),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_114),
.B(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_125),
.Y(n_252)
);

FAx1_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.CI(n_133),
.CON(n_125),
.SN(n_125)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_127),
.B(n_265),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_136),
.B(n_195),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_137),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_165),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_147),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_144),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_235),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_146),
.Y(n_235)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.C(n_151),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_149),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_150),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_237),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_231),
.B(n_236),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_216),
.B(n_230),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_197),
.B(n_215),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_185),
.B(n_196),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_174),
.B(n_184),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_166),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_170),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_187),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_199),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_206),
.B1(n_207),
.B2(n_214),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_200),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_201),
.A2(n_202),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_201),
.A2(n_202),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_201),
.A2(n_289),
.B(n_291),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_203),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_202),
.B(n_272),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_209),
.B(n_226),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_218),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_225),
.C(n_229),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_227),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_240),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_252),
.B2(n_253),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_247),
.C(n_253),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_245),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_257),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_274),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_270),
.B2(n_271),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_271),
.C(n_274),
.Y(n_277)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_263),
.C(n_269),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_267),
.B2(n_269),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_267),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_272),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_278),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_294),
.B2(n_295),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_285),
.B1(n_292),
.B2(n_293),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_293),
.C(n_295),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B(n_284),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_283),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_299),
.C(n_304),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_284),
.B(n_299),
.CI(n_304),
.CON(n_309),
.SN(n_309)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_290),
.B2(n_291),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_286),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_287),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_305),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_305),
.Y(n_311)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_309),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_309),
.Y(n_312)
);


endmodule