module fake_jpeg_4552_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_41),
.B1(n_24),
.B2(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_17),
.Y(n_45)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_44),
.B(n_51),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_17),
.B1(n_32),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_26),
.B1(n_24),
.B2(n_16),
.Y(n_90)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_19),
.B(n_18),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_22),
.B(n_32),
.C(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_61),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_60),
.A2(n_63),
.B1(n_24),
.B2(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_21),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_16),
.C(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_77),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_41),
.B1(n_35),
.B2(n_38),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_77),
.B1(n_53),
.B2(n_67),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_82),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_87),
.B(n_23),
.Y(n_101)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_38),
.B1(n_35),
.B2(n_26),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_94),
.B(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_96),
.Y(n_141)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_103),
.B1(n_104),
.B2(n_113),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_101),
.B1(n_114),
.B2(n_75),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_69),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_111),
.C(n_22),
.Y(n_137)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_69),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_108),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_107),
.B1(n_59),
.B2(n_97),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_35),
.B1(n_61),
.B2(n_66),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_72),
.B(n_47),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_92),
.B(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_47),
.B1(n_31),
.B2(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_42),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_43),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_118),
.Y(n_121)
);

BUFx2_ASAP7_75t_SL g120 ( 
.A(n_76),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_128),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_70),
.B1(n_86),
.B2(n_78),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_134),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_70),
.B1(n_78),
.B2(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_99),
.B1(n_119),
.B2(n_95),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

AOI22x1_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_47),
.B1(n_46),
.B2(n_56),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_68),
.B1(n_65),
.B2(n_55),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_98),
.B1(n_96),
.B2(n_103),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_80),
.B1(n_73),
.B2(n_55),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_145),
.C(n_109),
.Y(n_162)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_138),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_28),
.B(n_25),
.C(n_27),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_112),
.B(n_58),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_102),
.B(n_112),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_58),
.C(n_43),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_109),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_153),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_155),
.B1(n_169),
.B2(n_173),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_140),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_159),
.B(n_165),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_109),
.B(n_20),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_42),
.C(n_84),
.Y(n_192)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_124),
.B(n_118),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_174),
.B(n_19),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_43),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_43),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_146),
.B1(n_145),
.B2(n_135),
.Y(n_173)
);

AOI32xp33_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_84),
.A3(n_43),
.B1(n_42),
.B2(n_19),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_190),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_124),
.B1(n_136),
.B2(n_138),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_194),
.B1(n_165),
.B2(n_161),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_184),
.B(n_186),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_196),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_124),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_0),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_84),
.B(n_42),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_121),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_121),
.B(n_127),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_197),
.C(n_199),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_123),
.B(n_27),
.C(n_33),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_123),
.B1(n_25),
.B2(n_28),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_149),
.A2(n_19),
.B(n_20),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_0),
.Y(n_220)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_132),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_155),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_198),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_132),
.C(n_142),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_183),
.A2(n_170),
.B1(n_163),
.B2(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_152),
.B1(n_168),
.B2(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_161),
.B1(n_152),
.B2(n_148),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_213),
.B1(n_181),
.B2(n_187),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_165),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_210),
.B(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_214),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_154),
.B1(n_156),
.B2(n_33),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_186),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_192),
.C(n_191),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_218),
.C(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_33),
.C(n_20),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_1),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_225),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_175),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_232),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_185),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_209),
.C(n_223),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_209),
.B(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_185),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_242),
.Y(n_262)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_243),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_182),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_210),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_204),
.A2(n_187),
.B1(n_176),
.B2(n_180),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_213),
.B1(n_207),
.B2(n_189),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_248),
.B(n_254),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_227),
.A2(n_212),
.B(n_180),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_261),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_203),
.C(n_214),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_263),
.C(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_220),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_205),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_230),
.B1(n_235),
.B2(n_228),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_244),
.CI(n_236),
.CON(n_267),
.SN(n_267)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_10),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_273),
.B(n_275),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_237),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_5),
.Y(n_289)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

OA21x2_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_239),
.B(n_226),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_278),
.B1(n_276),
.B2(n_264),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_222),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_258),
.C(n_3),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_189),
.B1(n_240),
.B2(n_222),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_9),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_262),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_282),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_262),
.Y(n_280)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_281),
.A2(n_270),
.B(n_8),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_291),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_265),
.B(n_5),
.Y(n_291)
);

AOI31xp33_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_273),
.A3(n_267),
.B(n_275),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_298),
.B(n_300),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_270),
.B1(n_8),
.B2(n_11),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_299),
.Y(n_306)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_15),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_290),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_279),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_282),
.Y(n_307)
);

AOI31xp33_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_308),
.A3(n_309),
.B(n_12),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_298),
.B(n_294),
.C(n_11),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_7),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_313),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_312),
.B1(n_314),
.B2(n_306),
.Y(n_317)
);

AOI221xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_315),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_15),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_13),
.Y(n_320)
);


endmodule