module fake_jpeg_17727_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_73),
.Y(n_79)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_64),
.Y(n_81)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_52),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_47),
.B(n_54),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_95),
.B(n_0),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_57),
.B1(n_59),
.B2(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_53),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_54),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_62),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_59),
.B1(n_61),
.B2(n_65),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_67),
.B1(n_66),
.B2(n_50),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_109),
.B1(n_111),
.B2(n_117),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_119),
.B1(n_120),
.B2(n_6),
.Y(n_124)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_104),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_118),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_52),
.B1(n_49),
.B2(n_61),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_55),
.Y(n_115)
);

NOR2x1_ASAP7_75t_R g131 ( 
.A(n_115),
.B(n_122),
.Y(n_131)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_1),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_3),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_107),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_28),
.B(n_43),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_135),
.B1(n_10),
.B2(n_11),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_132),
.B1(n_115),
.B2(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_27),
.B1(n_42),
.B2(n_41),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_125),
.B(n_132),
.Y(n_145)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_141),
.B(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_145),
.A2(n_131),
.B(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_151),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_146),
.A2(n_139),
.B1(n_131),
.B2(n_126),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_134),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_130),
.B1(n_133),
.B2(n_114),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_143),
.B1(n_135),
.B2(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_156),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_153),
.B1(n_155),
.B2(n_12),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g161 ( 
.A(n_159),
.B(n_33),
.CON(n_161),
.SN(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_34),
.B(n_39),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_160),
.C(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_31),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_30),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_32),
.B(n_45),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_23),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_22),
.C(n_38),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_14),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_37),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_121),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_173),
.B(n_101),
.CI(n_112),
.CON(n_174),
.SN(n_174)
);


endmodule