module fake_netlist_5_1391_n_82 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_82);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_82;

wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_81;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_8),
.A2(n_6),
.B1(n_1),
.B2(n_7),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_10),
.Y(n_25)
);

AND2x6_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_7),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_17),
.A2(n_8),
.B1(n_15),
.B2(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_2),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_0),
.A2(n_3),
.B1(n_18),
.B2(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_26),
.Y(n_41)
);

OR2x6_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_28),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_24),
.B1(n_28),
.B2(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_30),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_32),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_42),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_23),
.C(n_35),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_26),
.B1(n_23),
.B2(n_35),
.Y(n_56)
);

NAND2x1p5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_26),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_49),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_60),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_50),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NAND4xp25_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_34),
.C(n_53),
.D(n_54),
.Y(n_69)
);

NOR4xp25_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_53),
.C(n_54),
.D(n_59),
.Y(n_70)
);

AOI211xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_29),
.B(n_50),
.C(n_35),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_50),
.B(n_56),
.C(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_47),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_66),
.B1(n_47),
.B2(n_65),
.Y(n_75)
);

NOR4xp25_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_65),
.C(n_26),
.D(n_23),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_26),
.C(n_73),
.Y(n_77)
);

NOR4xp25_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_40),
.C(n_44),
.D(n_34),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_75),
.B1(n_78),
.B2(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

OR2x6_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_79),
.Y(n_82)
);


endmodule