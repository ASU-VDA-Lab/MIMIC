module fake_jpeg_7235_n_258 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_37),
.Y(n_55)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_29),
.B1(n_34),
.B2(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_37),
.Y(n_74)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_23),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_62),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_28),
.B1(n_26),
.B2(n_22),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_32),
.B1(n_24),
.B2(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_27),
.B1(n_20),
.B2(n_33),
.Y(n_63)
);

NAND2x1_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_64),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_27),
.B1(n_20),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_17),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_27),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_81),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_26),
.B(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_87),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_17),
.B(n_19),
.Y(n_81)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_57),
.B1(n_37),
.B2(n_48),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_113),
.B1(n_35),
.B2(n_75),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_107),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_98),
.A2(n_93),
.B(n_87),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_49),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_106),
.Y(n_125)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_37),
.B1(n_65),
.B2(n_47),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_84),
.B1(n_75),
.B2(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_67),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_118),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_35),
.B1(n_36),
.B2(n_31),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_17),
.B1(n_19),
.B2(n_31),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_54),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_130),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_115),
.B1(n_35),
.B2(n_99),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_70),
.B1(n_88),
.B2(n_72),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_142),
.B1(n_95),
.B2(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_126),
.B(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_88),
.B(n_89),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_129),
.A2(n_139),
.B(n_116),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_88),
.B(n_76),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_141),
.B(n_99),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_98),
.A2(n_114),
.B1(n_118),
.B2(n_109),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_143),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_146),
.C(n_164),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_148),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_150),
.A2(n_159),
.B(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_157),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_122),
.B1(n_151),
.B2(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_160),
.B1(n_168),
.B2(n_138),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_128),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_95),
.A3(n_104),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_10),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_163),
.B1(n_122),
.B2(n_30),
.C(n_23),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_104),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_103),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_120),
.C(n_103),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_SL g192 ( 
.A(n_169),
.B(n_183),
.C(n_187),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_146),
.C(n_166),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_168),
.B1(n_161),
.B2(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_167),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_136),
.B1(n_140),
.B2(n_137),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_78),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_83),
.B1(n_120),
.B2(n_36),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_159),
.C(n_103),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_19),
.B(n_30),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_147),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_186),
.B(n_190),
.C(n_21),
.Y(n_200)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_159),
.A2(n_23),
.B(n_21),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVxp33_ASAP7_75t_SL g206 ( 
.A(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_144),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_196),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_204),
.B1(n_205),
.B2(n_190),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_178),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_201),
.C(n_203),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_36),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_22),
.C(n_21),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_187),
.B(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_54),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_188),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_53),
.C(n_52),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_53),
.C(n_52),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_78),
.B1(n_53),
.B2(n_52),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_85),
.B1(n_60),
.B2(n_6),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_184),
.C(n_170),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_214),
.C(n_222),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_213),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_183),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_177),
.B1(n_185),
.B2(n_171),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_16),
.B1(n_8),
.B2(n_10),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_219),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_200),
.B1(n_60),
.B2(n_7),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_170),
.C(n_60),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_197),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_226),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_192),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_207),
.C(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_230),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_231),
.B1(n_11),
.B2(n_12),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_200),
.C(n_5),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

OAI221xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_214),
.B1(n_221),
.B2(n_209),
.C(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_217),
.B1(n_209),
.B2(n_212),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_236),
.B(n_238),
.Y(n_242)
);

NOR2xp67_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_4),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_12),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_240),
.B(n_11),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_245),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_235),
.A2(n_230),
.B1(n_226),
.B2(n_227),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_238),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_247),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_12),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_SL g253 ( 
.A1(n_251),
.A2(n_242),
.B(n_14),
.C(n_15),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_253),
.A2(n_249),
.B1(n_14),
.B2(n_15),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_249),
.B(n_250),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_255),
.A2(n_256),
.B1(n_254),
.B2(n_13),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_13),
.Y(n_258)
);


endmodule