module fake_jpeg_4120_n_325 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_38),
.B(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_44),
.B1(n_52),
.B2(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_21),
.Y(n_57)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_48),
.Y(n_100)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_51),
.Y(n_87)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_14),
.C(n_21),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_57),
.B(n_58),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_35),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_35),
.B1(n_34),
.B2(n_31),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

OR2x2_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_11),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_62),
.B(n_70),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_64),
.Y(n_106)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_22),
.B1(n_18),
.B2(n_26),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_66),
.A2(n_83),
.B1(n_23),
.B2(n_29),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_49),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_79),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_76),
.Y(n_127)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_78),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_90),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_37),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_43),
.B(n_20),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_43),
.B(n_23),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_19),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_128),
.B1(n_24),
.B2(n_15),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_121),
.B(n_24),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_17),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_17),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_30),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_63),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_83),
.A2(n_29),
.B1(n_24),
.B2(n_30),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_67),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_137),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_118),
.B1(n_105),
.B2(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_141),
.B1(n_148),
.B2(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_143),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_62),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_147),
.B(n_171),
.Y(n_178)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_131),
.Y(n_140)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_60),
.B1(n_66),
.B2(n_83),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_67),
.B1(n_74),
.B2(n_88),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_142),
.A2(n_158),
.B1(n_163),
.B2(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_78),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_146),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_115),
.A2(n_54),
.B1(n_81),
.B2(n_84),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_149),
.B(n_153),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_68),
.B1(n_54),
.B2(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_59),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_164),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_154),
.B(n_155),
.Y(n_205)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_80),
.B(n_101),
.C(n_87),
.D(n_55),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_97),
.C(n_101),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_108),
.C(n_111),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_87),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_129),
.B1(n_126),
.B2(n_103),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_123),
.B(n_69),
.Y(n_159)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_114),
.A2(n_65),
.B1(n_30),
.B2(n_15),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_85),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_130),
.A2(n_94),
.B1(n_89),
.B2(n_71),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_85),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_0),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_94),
.B1(n_71),
.B2(n_99),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_3),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_106),
.B(n_76),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_108),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_99),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_177),
.C(n_186),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_110),
.B(n_129),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_179),
.A2(n_180),
.B(n_182),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_110),
.B(n_111),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_107),
.B1(n_102),
.B2(n_103),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_7),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_125),
.B(n_107),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_189),
.B(n_166),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_125),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_195),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_102),
.B(n_2),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_119),
.C(n_2),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_198),
.C(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_1),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_119),
.C(n_9),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_119),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_202),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_1),
.C(n_2),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_144),
.B(n_5),
.C(n_7),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_9),
.C(n_10),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_5),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_217),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_176),
.B(n_165),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_176),
.B(n_153),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_173),
.A2(n_141),
.B1(n_139),
.B2(n_162),
.Y(n_213)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_155),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_231),
.C(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_224),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_146),
.B1(n_135),
.B2(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_138),
.Y(n_222)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_140),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_180),
.B1(n_185),
.B2(n_189),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_7),
.B(n_8),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_234),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_229),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_230),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_174),
.C(n_198),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_10),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_11),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_12),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_236),
.B(n_238),
.Y(n_270)
);

A2O1A1O1Ixp25_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_186),
.B(n_192),
.C(n_179),
.D(n_205),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_219),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_249),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_209),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_251),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_228),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_249),
.B1(n_244),
.B2(n_245),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_257),
.C(n_215),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_177),
.C(n_191),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_265),
.C(n_268),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_240),
.Y(n_286)
);

AOI221xp5_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_218),
.B1(n_224),
.B2(n_210),
.C(n_211),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_267),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_266),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_211),
.C(n_223),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_224),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_242),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_258),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_206),
.B1(n_217),
.B2(n_182),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_223),
.C(n_212),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_241),
.C(n_245),
.Y(n_280)
);

OAI321xp33_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_202),
.A3(n_193),
.B1(n_226),
.B2(n_216),
.C(n_196),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_282),
.C(n_284),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_243),
.C(n_234),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_193),
.C(n_222),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_236),
.B1(n_196),
.B2(n_199),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_289),
.B(n_199),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_287),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_260),
.B(n_237),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_227),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_298),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_267),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_248),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_272),
.C(n_268),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_270),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_264),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_240),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_197),
.B1(n_190),
.B2(n_214),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_288),
.B(n_279),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_302),
.C(n_309),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_238),
.B1(n_252),
.B2(n_239),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_230),
.B1(n_220),
.B2(n_214),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_307),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_292),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_291),
.B(n_201),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_301),
.C(n_294),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_313),
.C(n_314),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_292),
.B1(n_279),
.B2(n_190),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_316),
.B1(n_197),
.B2(n_184),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_291),
.C(n_231),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_310),
.C(n_308),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_184),
.C(n_12),
.Y(n_321)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_318),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_315),
.B(n_184),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_322),
.Y(n_325)
);


endmodule