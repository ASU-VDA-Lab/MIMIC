module fake_jpeg_25502_n_33 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_1),
.A2(n_5),
.B1(n_0),
.B2(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_19),
.B1(n_22),
.B2(n_13),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_3),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_14),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_16),
.Y(n_23)
);

AOI322xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_18),
.A3(n_22),
.B1(n_19),
.B2(n_21),
.C1(n_14),
.C2(n_12),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_22),
.Y(n_28)
);

A2O1A1O1Ixp25_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_23),
.B(n_26),
.C(n_24),
.D(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_14),
.B1(n_9),
.B2(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_29),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_25),
.C1(n_30),
.C2(n_29),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);


endmodule