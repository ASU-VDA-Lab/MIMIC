module fake_ariane_1435_n_272 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_272);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_272;

wire n_83;
wire n_233;
wire n_56;
wire n_60;
wire n_190;
wire n_170;
wire n_160;
wire n_64;
wire n_179;
wire n_240;
wire n_124;
wire n_119;
wire n_180;
wire n_167;
wire n_90;
wire n_195;
wire n_213;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_221;
wire n_86;
wire n_269;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_158;
wire n_237;
wire n_172;
wire n_69;
wire n_259;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_203;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_242;
wire n_260;
wire n_115;
wire n_133;
wire n_66;
wire n_205;
wire n_236;
wire n_265;
wire n_71;
wire n_267;
wire n_109;
wire n_208;
wire n_245;
wire n_96;
wire n_156;
wire n_209;
wire n_49;
wire n_262;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_210;
wire n_147;
wire n_204;
wire n_225;
wire n_235;
wire n_200;
wire n_51;
wire n_166;
wire n_253;
wire n_76;
wire n_218;
wire n_103;
wire n_79;
wire n_246;
wire n_226;
wire n_244;
wire n_271;
wire n_46;
wire n_220;
wire n_84;
wire n_247;
wire n_261;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_217;
wire n_44;
wire n_224;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_263;
wire n_201;
wire n_229;
wire n_70;
wire n_250;
wire n_222;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_256;
wire n_214;
wire n_227;
wire n_48;
wire n_101;
wire n_94;
wire n_243;
wire n_134;
wire n_188;
wire n_185;
wire n_249;
wire n_58;
wire n_65;
wire n_123;
wire n_212;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_264;
wire n_129;
wire n_126;
wire n_137;
wire n_255;
wire n_122;
wire n_268;
wire n_257;
wire n_266;
wire n_198;
wire n_148;
wire n_232;
wire n_164;
wire n_52;
wire n_157;
wire n_248;
wire n_184;
wire n_177;
wire n_135;
wire n_258;
wire n_73;
wire n_77;
wire n_171;
wire n_228;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_206;
wire n_207;
wire n_241;
wire n_254;
wire n_238;
wire n_41;
wire n_219;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_231;
wire n_192;
wire n_80;
wire n_146;
wire n_234;
wire n_230;
wire n_211;
wire n_270;
wire n_194;
wire n_97;
wire n_154;
wire n_215;
wire n_252;
wire n_142;
wire n_251;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_202;
wire n_145;
wire n_78;
wire n_193;
wire n_63;
wire n_59;
wire n_99;
wire n_216;
wire n_155;
wire n_127;
wire n_239;
wire n_223;
wire n_54;

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g57 ( 
.A(n_12),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_14),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_29),
.Y(n_66)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_0),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_1),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_1),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_2),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_53),
.B(n_3),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_58),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_44),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_57),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_50),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_45),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_41),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_4),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_48),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_114)
);

O2A1O1Ixp5_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_81),
.B(n_77),
.C(n_74),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_104),
.B(n_111),
.C(n_114),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_110),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_87),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_87),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_103),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_81),
.Y(n_132)
);

NOR2x2_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_97),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_109),
.B(n_75),
.C(n_77),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_109),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_129),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_124),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_132),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_107),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_98),
.B1(n_105),
.B2(n_94),
.Y(n_149)
);

AND2x4_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_75),
.Y(n_151)
);

NAND2x1p5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_73),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_86),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_125),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_69),
.B(n_92),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

OR2x6_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_119),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

AO21x2_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_73),
.B(n_133),
.Y(n_161)
);

BUFx2_ASAP7_75t_SL g162 ( 
.A(n_137),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_144),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_69),
.B(n_25),
.Y(n_167)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_69),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_24),
.B(n_38),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_152),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_140),
.B1(n_138),
.B2(n_147),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_138),
.Y(n_183)
);

OAI211xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_149),
.B(n_145),
.C(n_139),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_142),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_142),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_139),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_164),
.B1(n_159),
.B2(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_170),
.C(n_153),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_165),
.Y(n_196)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

OAI222xp33_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_159),
.B1(n_152),
.B2(n_172),
.C1(n_150),
.C2(n_164),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_171),
.B1(n_159),
.B2(n_137),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_159),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_137),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_206),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_186),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

OR2x6_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_214),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_197),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_192),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_174),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_234),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_167),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_167),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_195),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_220),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_214),
.Y(n_244)
);

NOR2x1p5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_173),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_233),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_231),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_231),
.C(n_230),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_173),
.C(n_193),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_155),
.C(n_198),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_231),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_242),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_245),
.B(n_247),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_244),
.B1(n_177),
.B2(n_192),
.Y(n_257)
);

AOI221xp5_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_243),
.B1(n_239),
.B2(n_237),
.C(n_151),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_254),
.B(n_253),
.C(n_250),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_258),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_257),
.Y(n_262)
);

AND3x1_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_237),
.C(n_239),
.Y(n_263)
);

NAND4xp75_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_169),
.C(n_167),
.D(n_172),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_SL g265 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_265)
);

AOI321xp33_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_180),
.A3(n_185),
.B1(n_166),
.B2(n_181),
.C(n_154),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_266),
.A2(n_169),
.B(n_162),
.Y(n_267)
);

OAI211xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_137),
.B(n_10),
.C(n_11),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_19),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_31),
.B(n_33),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

OR2x6_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_270),
.Y(n_272)
);


endmodule