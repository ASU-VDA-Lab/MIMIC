module fake_jpeg_1686_n_396 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_6),
.B(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_54),
.B(n_60),
.Y(n_159)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_6),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_63),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_68),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_78),
.Y(n_118)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_76),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_21),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_79),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_81),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_87),
.Y(n_128)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_4),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_29),
.A2(n_34),
.B1(n_53),
.B2(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_88),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_24),
.B(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_89),
.B(n_91),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_28),
.B(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_92),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_13),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_15),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_16),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_96),
.B(n_47),
.Y(n_146)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_25),
.B(n_16),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_98),
.B(n_99),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_25),
.B(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_107),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_40),
.B(n_16),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_109),
.Y(n_141)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_20),
.B1(n_30),
.B2(n_51),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_111),
.A2(n_166),
.B1(n_172),
.B2(n_122),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_51),
.B1(n_50),
.B2(n_45),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_57),
.A2(n_44),
.B1(n_39),
.B2(n_47),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_115),
.A2(n_135),
.B1(n_147),
.B2(n_160),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_30),
.B1(n_20),
.B2(n_44),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g194 ( 
.A1(n_119),
.A2(n_160),
.A3(n_147),
.B1(n_115),
.B2(n_124),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_41),
.B(n_48),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_125),
.B(n_143),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_50),
.B1(n_31),
.B2(n_38),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_130),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_75),
.A2(n_39),
.B1(n_48),
.B2(n_46),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_31),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_144),
.B(n_145),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_61),
.B(n_45),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_61),
.B(n_0),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_0),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_152),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_85),
.A2(n_69),
.B1(n_107),
.B2(n_76),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_151),
.A2(n_173),
.B1(n_155),
.B2(n_124),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_58),
.B(n_2),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_64),
.B(n_2),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_67),
.B(n_2),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_77),
.A2(n_86),
.B1(n_104),
.B2(n_103),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_55),
.A2(n_80),
.B1(n_95),
.B2(n_102),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_68),
.B(n_70),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_148),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_71),
.B(n_106),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_172),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_81),
.A2(n_93),
.B1(n_88),
.B2(n_43),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_186),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_180),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_182),
.A2(n_214),
.B1(n_205),
.B2(n_232),
.Y(n_234)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_114),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_187),
.B(n_196),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_128),
.A2(n_139),
.B1(n_119),
.B2(n_126),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_194),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_113),
.B(n_173),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_191),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_159),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_116),
.B(n_120),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_117),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_223),
.C(n_227),
.Y(n_250)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_118),
.B(n_157),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_201),
.B(n_216),
.Y(n_238)
);

BUFx8_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_202),
.B(n_215),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_168),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_206),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_119),
.A2(n_135),
.B1(n_142),
.B2(n_127),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_205),
.A2(n_221),
.B1(n_232),
.B2(n_225),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_164),
.B(n_167),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_148),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_130),
.B(n_134),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_209),
.B(n_229),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_127),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_132),
.A2(n_140),
.B1(n_142),
.B2(n_134),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_211),
.A2(n_212),
.B1(n_221),
.B2(n_200),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_132),
.A2(n_140),
.B1(n_112),
.B2(n_138),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_112),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_129),
.B(n_169),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_219),
.B(n_215),
.Y(n_255)
);

INVx4_ASAP7_75t_SL g220 ( 
.A(n_169),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_224),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_174),
.A2(n_138),
.B1(n_165),
.B2(n_110),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_153),
.A2(n_165),
.B(n_156),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_110),
.B(n_156),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_153),
.A2(n_131),
.B(n_174),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_231),
.B(n_177),
.C(n_223),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_131),
.A2(n_141),
.B(n_128),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_146),
.B(n_136),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_183),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_137),
.B(n_150),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_137),
.B(n_150),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_202),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_128),
.A2(n_136),
.B(n_143),
.C(n_141),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_111),
.A2(n_88),
.B1(n_166),
.B2(n_137),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_234),
.A2(n_256),
.B1(n_259),
.B2(n_271),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_182),
.B1(n_222),
.B2(n_209),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_239),
.A2(n_241),
.B1(n_237),
.B2(n_247),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_226),
.B1(n_189),
.B2(n_194),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_199),
.A2(n_226),
.B(n_185),
.C(n_188),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_243),
.A2(n_237),
.B(n_241),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_196),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_202),
.C(n_250),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_227),
.B(n_231),
.CI(n_178),
.CON(n_253),
.SN(n_253)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_253),
.B(n_263),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_229),
.A2(n_230),
.B1(n_179),
.B2(n_181),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_187),
.B(n_203),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_217),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_268),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_220),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_197),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_193),
.A2(n_195),
.B1(n_184),
.B2(n_192),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_245),
.B(n_180),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_273),
.B(n_291),
.Y(n_304)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_242),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_284),
.Y(n_313)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_282),
.A2(n_284),
.B(n_301),
.Y(n_314)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_260),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_285),
.A2(n_240),
.B(n_253),
.Y(n_311)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_254),
.Y(n_286)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_250),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_288),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_235),
.B(n_238),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_235),
.B(n_238),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_296),
.Y(n_317)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_270),
.C(n_233),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_298),
.Y(n_319)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_246),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_236),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_301),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_264),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_234),
.B(n_247),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_302),
.B(n_262),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_256),
.B1(n_243),
.B2(n_249),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_305),
.A2(n_320),
.B1(n_277),
.B2(n_291),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_274),
.A2(n_243),
.B1(n_253),
.B2(n_240),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_322),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_311),
.A2(n_324),
.B(n_325),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_314),
.B(n_282),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_274),
.A2(n_271),
.B1(n_262),
.B2(n_252),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_263),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_285),
.A2(n_262),
.B(n_258),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_289),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_278),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_287),
.C(n_280),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_334),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_302),
.B(n_300),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_330),
.A2(n_341),
.B(n_304),
.Y(n_353)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_333),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_297),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_335),
.B(n_336),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_306),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_273),
.C(n_288),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_337),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_272),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_272),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_305),
.A2(n_277),
.B1(n_303),
.B2(n_279),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_306),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_305),
.A2(n_275),
.B1(n_293),
.B2(n_292),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_342),
.A2(n_304),
.B1(n_315),
.B2(n_321),
.Y(n_352)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_343),
.A2(n_344),
.B1(n_315),
.B2(n_318),
.Y(n_357)
);

NOR3xp33_ASAP7_75t_SL g344 ( 
.A(n_308),
.B(n_292),
.C(n_281),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_331),
.A2(n_309),
.B1(n_310),
.B2(n_320),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_346),
.A2(n_349),
.B1(n_352),
.B2(n_357),
.Y(n_363)
);

AOI322xp5_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_314),
.A3(n_308),
.B1(n_319),
.B2(n_322),
.C1(n_324),
.C2(n_310),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_347),
.A2(n_351),
.B(n_353),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_330),
.A2(n_320),
.B1(n_326),
.B2(n_275),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_328),
.A2(n_325),
.B(n_317),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_328),
.A2(n_317),
.B(n_321),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_358),
.B(n_343),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_350),
.B(n_334),
.Y(n_359)
);

NAND3xp33_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_362),
.C(n_345),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_327),
.C(n_337),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_365),
.C(n_366),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_339),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_368),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_350),
.B(n_344),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_356),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_356),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_338),
.C(n_329),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_342),
.C(n_340),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_333),
.C(n_307),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_358),
.C(n_351),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_377),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_369),
.A2(n_349),
.B1(n_346),
.B2(n_352),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_353),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_375),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_360),
.B(n_357),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_376),
.B(n_365),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_368),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_379),
.A2(n_371),
.B(n_372),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_380),
.B(n_382),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_361),
.Y(n_382)
);

AOI21x1_ASAP7_75t_L g389 ( 
.A1(n_384),
.A2(n_388),
.B(n_367),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_381),
.A2(n_379),
.B(n_378),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_387),
.C(n_348),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_372),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_378),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_391),
.B(n_390),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_363),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_390),
.B(n_386),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_393),
.C(n_307),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_332),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_316),
.Y(n_396)
);


endmodule