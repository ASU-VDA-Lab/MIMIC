module fake_jpeg_28844_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_5),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_0),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_54),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_78),
.Y(n_84)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_70),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_57),
.B1(n_55),
.B2(n_51),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_87),
.B1(n_76),
.B2(n_77),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_68),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_57),
.B1(n_64),
.B2(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_62),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_71),
.A2(n_65),
.B(n_59),
.C(n_64),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_93),
.B(n_82),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_64),
.CON(n_93),
.SN(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_93),
.B1(n_83),
.B2(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_98),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_58),
.C(n_60),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_8),
.C(n_10),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_67),
.Y(n_98)
);

NOR2x1_ASAP7_75t_R g127 ( 
.A(n_99),
.B(n_16),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_61),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_103),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_63),
.B1(n_3),
.B2(n_4),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_63),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_0),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_108),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_1),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_24),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_2),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_115),
.B1(n_123),
.B2(n_100),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_6),
.B(n_7),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_122),
.B(n_113),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_28),
.C(n_46),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_8),
.B(n_11),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_127),
.A2(n_104),
.B(n_97),
.Y(n_131)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NAND2x1p5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_17),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_38),
.B(n_39),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_136),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_25),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_31),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_33),
.B(n_34),
.Y(n_141)
);

NOR2xp67_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_36),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_130),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_146),
.A2(n_135),
.B1(n_134),
.B2(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_125),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_154),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_142),
.C(n_140),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_152),
.B(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_154),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_156),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_149),
.B(n_142),
.C(n_151),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_148),
.B(n_120),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_148),
.Y(n_162)
);


endmodule