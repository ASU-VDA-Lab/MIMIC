module fake_jpeg_14309_n_482 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_482);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_482;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_66),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_73),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_0),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_63),
.B(n_80),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_16),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_17),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_75),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_31),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_82),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_2),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_41),
.C(n_44),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_18),
.B(n_2),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_18),
.B(n_2),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_84),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_3),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_37),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_21),
.B(n_3),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_95),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_22),
.B(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_56),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_109),
.A2(n_46),
.B1(n_36),
.B2(n_30),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_37),
.B(n_40),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_111),
.B(n_148),
.C(n_39),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_31),
.B1(n_34),
.B2(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_118),
.B1(n_144),
.B2(n_147),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_50),
.A2(n_24),
.B1(n_41),
.B2(n_34),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_49),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_123),
.Y(n_173)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_125),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_25),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_138),
.B(n_39),
.Y(n_155)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_145),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_72),
.A2(n_41),
.B1(n_37),
.B2(n_48),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_78),
.A2(n_37),
.B1(n_32),
.B2(n_48),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_91),
.A2(n_32),
.B1(n_47),
.B2(n_23),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_55),
.B1(n_93),
.B2(n_92),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_40),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_155),
.B(n_163),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_119),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_75),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_160),
.B(n_161),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_106),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_117),
.B(n_52),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_120),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_87),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_165),
.B(n_169),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_83),
.B(n_76),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_166),
.A2(n_29),
.B(n_28),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_66),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_168),
.B(n_177),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_102),
.B(n_60),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_181),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_69),
.B1(n_65),
.B2(n_68),
.Y(n_215)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_176),
.B(n_180),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_54),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_108),
.B(n_61),
.C(n_86),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_113),
.B(n_85),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_115),
.B(n_77),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_110),
.B(n_71),
.C(n_93),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_121),
.B(n_29),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_146),
.A3(n_136),
.B1(n_104),
.B2(n_126),
.Y(n_206)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_57),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_187),
.Y(n_233)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_64),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_188),
.Y(n_208)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_28),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_30),
.Y(n_235)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_101),
.B1(n_143),
.B2(n_112),
.Y(n_230)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_104),
.A2(n_53),
.B1(n_51),
.B2(n_32),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_70),
.B1(n_101),
.B2(n_99),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_172),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_211),
.B(n_235),
.Y(n_243)
);

AO21x2_ASAP7_75t_L g212 ( 
.A1(n_166),
.A2(n_144),
.B(n_147),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_212),
.A2(n_220),
.B(n_175),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_172),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_67),
.B1(n_131),
.B2(n_126),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_222),
.B1(n_230),
.B2(n_180),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_156),
.A2(n_131),
.B1(n_146),
.B2(n_149),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_157),
.A2(n_107),
.B(n_22),
.C(n_25),
.Y(n_225)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_170),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_236),
.B(n_237),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_153),
.B1(n_159),
.B2(n_179),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_238),
.A2(n_253),
.B1(n_112),
.B2(n_143),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_182),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_184),
.B1(n_153),
.B2(n_178),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_240),
.A2(n_246),
.B1(n_215),
.B2(n_209),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_161),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_247),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_159),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_256),
.C(n_257),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_252),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_181),
.B(n_188),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_264),
.B(n_269),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_172),
.B1(n_151),
.B2(n_154),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_173),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_248),
.A2(n_231),
.B1(n_205),
.B2(n_120),
.Y(n_295)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_251),
.B(n_255),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_220),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_180),
.B1(n_167),
.B2(n_154),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_199),
.B(n_167),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_170),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_186),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_185),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_158),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_169),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_209),
.A2(n_195),
.B1(n_152),
.B2(n_183),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_213),
.B(n_129),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_266),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_190),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_238),
.A2(n_212),
.B1(n_215),
.B2(n_206),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_272),
.A2(n_279),
.B1(n_298),
.B2(n_300),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_219),
.C(n_222),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_256),
.C(n_245),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_237),
.A2(n_212),
.B1(n_215),
.B2(n_225),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_243),
.B(n_262),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_281),
.B(n_282),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_208),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_234),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_284),
.B(n_293),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_285),
.A2(n_296),
.B1(n_274),
.B2(n_294),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_239),
.B(n_221),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_258),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_301),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_295),
.A2(n_254),
.B(n_249),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_240),
.B(n_207),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_296),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_236),
.A2(n_194),
.B1(n_140),
.B2(n_229),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_258),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_205),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_303),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_249),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_251),
.B(n_232),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_227),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_306),
.B(n_319),
.Y(n_352)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_271),
.Y(n_307)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_284),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_308),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_272),
.A2(n_292),
.B1(n_279),
.B2(n_298),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_325),
.B1(n_334),
.B2(n_286),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_302),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_312),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_257),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_316),
.C(n_322),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_269),
.B1(n_246),
.B2(n_248),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_314),
.A2(n_326),
.B1(n_278),
.B2(n_301),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_275),
.B(n_253),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_317),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_303),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_304),
.A2(n_260),
.B(n_248),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_321),
.A2(n_328),
.B(n_330),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_266),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g323 ( 
.A(n_273),
.B(n_265),
.Y(n_323)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_260),
.B1(n_261),
.B2(n_268),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_232),
.C(n_201),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_331),
.C(n_293),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_275),
.A2(n_296),
.B(n_292),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_273),
.B(n_201),
.Y(n_329)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_329),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_274),
.A2(n_204),
.B(n_207),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_196),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_300),
.A2(n_229),
.B1(n_202),
.B2(n_162),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_336),
.B(n_227),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_322),
.B(n_313),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_341),
.B(n_348),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_343),
.A2(n_311),
.B1(n_329),
.B2(n_325),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_281),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_356),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_278),
.B1(n_287),
.B2(n_277),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_345),
.A2(n_346),
.B1(n_349),
.B2(n_315),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_326),
.A2(n_277),
.B1(n_283),
.B2(n_289),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_331),
.B(n_291),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_283),
.B1(n_289),
.B2(n_291),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_329),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_351),
.A2(n_353),
.B1(n_355),
.B2(n_306),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_305),
.A2(n_276),
.B1(n_290),
.B2(n_299),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_276),
.B1(n_299),
.B2(n_297),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_297),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_323),
.B(n_189),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_359),
.B(n_317),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_204),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_366),
.C(n_328),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_319),
.Y(n_373)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_364),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_221),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_369),
.A2(n_376),
.B1(n_174),
.B2(n_140),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_372),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_371),
.Y(n_396)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_317),
.C(n_309),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_378),
.C(n_385),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_379),
.B1(n_23),
.B2(n_4),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_309),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_360),
.A2(n_308),
.B1(n_312),
.B2(n_307),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_365),
.A2(n_330),
.B(n_321),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_380),
.B(n_381),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_338),
.B(n_332),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_348),
.B(n_332),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_386),
.Y(n_410)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

O2A1O1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_363),
.A2(n_365),
.B(n_343),
.C(n_337),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_47),
.B(n_43),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_318),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_342),
.B(n_335),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_361),
.C(n_356),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_388),
.C(n_390),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_357),
.A2(n_324),
.B1(n_320),
.B2(n_334),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_389),
.A2(n_347),
.B1(n_346),
.B2(n_363),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_202),
.C(n_162),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_349),
.Y(n_391)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

XNOR2x1_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_127),
.Y(n_392)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_392),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_393),
.A2(n_398),
.B1(n_411),
.B2(n_412),
.Y(n_421)
);

NOR3xp33_ASAP7_75t_SL g394 ( 
.A(n_377),
.B(n_337),
.C(n_354),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_401),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_339),
.Y(n_397)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_397),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_390),
.A2(n_339),
.B1(n_358),
.B2(n_366),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_404),
.A2(n_407),
.B1(n_402),
.B2(n_396),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_372),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_408),
.B(n_413),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_409),
.B(n_4),
.Y(n_425)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_387),
.C(n_378),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_415),
.B(n_418),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_385),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_417),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_367),
.C(n_368),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_367),
.C(n_368),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_382),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_419),
.B(n_426),
.Y(n_431)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_420),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_392),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_422),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_370),
.C(n_127),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_427),
.C(n_399),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_393),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_127),
.C(n_58),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_46),
.C(n_36),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_410),
.B(n_6),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_409),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_46),
.Y(n_430)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_430),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_438),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_436),
.A2(n_429),
.B(n_428),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_424),
.A2(n_401),
.B(n_397),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_444),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_399),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_427),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_414),
.A2(n_402),
.B(n_404),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_10),
.C(n_11),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_422),
.A2(n_394),
.B(n_8),
.Y(n_442)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_46),
.C(n_36),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_46),
.C(n_36),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_36),
.C(n_12),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_437),
.B(n_425),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_448),
.B(n_455),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_459),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_433),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_452),
.A2(n_434),
.B1(n_435),
.B2(n_431),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_436),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_454),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_438),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_30),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_457),
.B(n_11),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_464),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_450),
.B(n_443),
.Y(n_465)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_465),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_440),
.Y(n_466)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_466),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_432),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_467),
.A2(n_456),
.B(n_453),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_474),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_441),
.C(n_445),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_462),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_460),
.A2(n_458),
.B(n_454),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_475),
.A2(n_470),
.B(n_473),
.Y(n_478)
);

AOI321xp33_ASAP7_75t_L g477 ( 
.A1(n_469),
.A2(n_467),
.A3(n_468),
.B1(n_444),
.B2(n_452),
.C(n_459),
.Y(n_477)
);

AOI321xp33_ASAP7_75t_L g479 ( 
.A1(n_477),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_475),
.C(n_462),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_478),
.A2(n_479),
.B(n_476),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_480),
.B(n_13),
.C(n_14),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g482 ( 
.A(n_481),
.Y(n_482)
);


endmodule