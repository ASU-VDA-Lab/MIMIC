module fake_ariane_900_n_897 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_897);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_897;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_819;
wire n_189;
wire n_717;
wire n_706;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_705;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_847;
wire n_772;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_97),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_10),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_47),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_39),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_136),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_61),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_38),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_44),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_67),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_23),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_1),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_54),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_12),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_56),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_36),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_100),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_5),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_26),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_116),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_53),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_79),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_156),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_64),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_112),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_167),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_13),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_57),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_122),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_4),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_14),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_51),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_92),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_35),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_27),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_164),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_121),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_29),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_91),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_71),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_40),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_98),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_43),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_160),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_139),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_68),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_130),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_171),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_8),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_155),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_66),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_52),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_135),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_28),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_83),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_175),
.Y(n_261)
);

NOR2xp67_ASAP7_75t_L g262 ( 
.A(n_37),
.B(n_17),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_173),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_58),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_55),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_19),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_105),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

BUFx8_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_224),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_211),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_198),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_0),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_185),
.B(n_187),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_261),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_191),
.B(n_2),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

BUFx8_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_205),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_229),
.B(n_3),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_225),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_188),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_3),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_194),
.B(n_4),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_195),
.B(n_196),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_188),
.A2(n_95),
.B(n_183),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_225),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_200),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_233),
.B(n_5),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_204),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_217),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_253),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_204),
.A2(n_96),
.B(n_182),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_228),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_304)
);

NOR2x1_ASAP7_75t_L g305 ( 
.A(n_201),
.B(n_20),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_208),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_203),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_208),
.B(n_6),
.Y(n_308)
);

CKINVDCx11_ASAP7_75t_R g309 ( 
.A(n_235),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_207),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_212),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_220),
.Y(n_313)
);

BUFx12f_ASAP7_75t_L g314 ( 
.A(n_186),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_244),
.B(n_255),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_225),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_225),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_234),
.A2(n_99),
.B(n_181),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_237),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_269),
.A2(n_236),
.B1(n_192),
.B2(n_266),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_270),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_276),
.B(n_241),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_241),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_276),
.B(n_197),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_245),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_280),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_276),
.B(n_250),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_270),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_271),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_271),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_308),
.B(n_193),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_271),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_292),
.B(n_199),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_271),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_279),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_265),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_281),
.B(n_213),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_283),
.B(n_202),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_271),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_283),
.B(n_254),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_318),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_SL g357 ( 
.A(n_287),
.B(n_291),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_281),
.B(n_206),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_285),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_285),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_287),
.B(n_256),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_284),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_284),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_289),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_286),
.B(n_210),
.Y(n_370)
);

OR2x6_ASAP7_75t_L g371 ( 
.A(n_273),
.B(n_257),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_290),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_289),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_284),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_315),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_300),
.B(n_263),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_352),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_349),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_349),
.Y(n_379)
);

OR2x6_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_268),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_365),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_283),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_365),
.A2(n_304),
.B1(n_291),
.B2(n_298),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_328),
.B(n_297),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_357),
.A2(n_351),
.B1(n_328),
.B2(n_339),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_340),
.B(n_297),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_340),
.B(n_312),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_340),
.B(n_312),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_360),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_274),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_314),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_331),
.B(n_274),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_376),
.B(n_278),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_288),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_278),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_324),
.B(n_322),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_288),
.Y(n_406)
);

O2A1O1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_339),
.A2(n_298),
.B(n_320),
.C(n_313),
.Y(n_407)
);

OAI22xp33_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_286),
.B1(n_268),
.B2(n_323),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_357),
.A2(n_323),
.B1(n_307),
.B2(n_311),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_L g410 ( 
.A1(n_371),
.A2(n_314),
.B1(n_319),
.B2(n_306),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_331),
.B(n_306),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_355),
.B(n_269),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_351),
.B(n_306),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_345),
.A2(n_296),
.B(n_295),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_345),
.A2(n_294),
.B(n_303),
.C(n_321),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_356),
.B(n_295),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_326),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_353),
.B(n_269),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_347),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_325),
.B(n_215),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_337),
.B(n_216),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_346),
.B(n_319),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_346),
.B(n_319),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_346),
.B(n_290),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_326),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_344),
.B(n_218),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_333),
.B(n_290),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_341),
.B(n_290),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_341),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_342),
.B(n_219),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g437 ( 
.A(n_342),
.B(n_305),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_343),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_371),
.A2(n_264),
.B1(n_222),
.B2(n_252),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_343),
.B(n_296),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_348),
.B(n_302),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_354),
.A2(n_258),
.B1(n_227),
.B2(n_231),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_354),
.B(n_290),
.Y(n_444)
);

CKINVDCx10_ASAP7_75t_R g445 ( 
.A(n_380),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_383),
.B(n_299),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_383),
.B(n_299),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_394),
.B(n_223),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_395),
.B(n_299),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_402),
.A2(n_303),
.B(n_294),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_402),
.A2(n_321),
.B(n_369),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_406),
.A2(n_405),
.B(n_421),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_388),
.B(n_238),
.Y(n_454)
);

AOI21x1_ASAP7_75t_L g455 ( 
.A1(n_417),
.A2(n_302),
.B(n_316),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_412),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_418),
.A2(n_407),
.B(n_406),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_405),
.A2(n_373),
.B(n_369),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_429),
.A2(n_373),
.B(n_368),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_384),
.B(n_239),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_424),
.A2(n_317),
.B(n_316),
.C(n_363),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_389),
.A2(n_368),
.B(n_364),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_392),
.B(n_299),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_393),
.A2(n_364),
.B(n_363),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_392),
.B(n_299),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_409),
.B(n_310),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_427),
.A2(n_362),
.B(n_361),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_444),
.Y(n_468)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_440),
.A2(n_317),
.B(n_361),
.Y(n_469)
);

BUFx2_ASAP7_75t_SL g470 ( 
.A(n_396),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_403),
.A2(n_362),
.B(n_359),
.C(n_358),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_L g472 ( 
.A(n_377),
.B(n_310),
.Y(n_472)
);

AOI21x1_ASAP7_75t_L g473 ( 
.A1(n_440),
.A2(n_359),
.B(n_358),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_398),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_426),
.A2(n_344),
.B(n_248),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_386),
.A2(n_425),
.B1(n_419),
.B2(n_382),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_399),
.B(n_309),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_415),
.A2(n_344),
.B(n_247),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_416),
.B(n_310),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_420),
.A2(n_246),
.B(n_242),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_386),
.A2(n_310),
.B1(n_309),
.B2(n_259),
.Y(n_482)
);

A2O1A1Ixp33_ASAP7_75t_L g483 ( 
.A1(n_439),
.A2(n_310),
.B(n_251),
.C(n_243),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_397),
.B(n_240),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_404),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_423),
.B(n_7),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_414),
.B(n_9),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_442),
.A2(n_289),
.B(n_101),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_401),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_379),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_94),
.B(n_180),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_385),
.A2(n_387),
.B(n_428),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_410),
.B(n_9),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_380),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_400),
.Y(n_499)
);

O2A1O1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_411),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_380),
.B(n_408),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_422),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_437),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_443),
.B(n_435),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_434),
.A2(n_103),
.B(n_179),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_437),
.B(n_11),
.Y(n_508)
);

O2A1O1Ixp33_ASAP7_75t_L g509 ( 
.A1(n_431),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_509)
);

AOI21xp33_ASAP7_75t_L g510 ( 
.A1(n_432),
.A2(n_15),
.B(n_16),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_17),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_433),
.A2(n_106),
.B(n_21),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_441),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_437),
.B(n_18),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_438),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_L g516 ( 
.A1(n_488),
.A2(n_436),
.B(n_413),
.C(n_18),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_451),
.A2(n_413),
.B(n_24),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_506),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_455),
.A2(n_452),
.B(n_473),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_477),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g521 ( 
.A1(n_457),
.A2(n_184),
.B(n_25),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_469),
.A2(n_22),
.B(n_30),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_453),
.A2(n_31),
.B(n_33),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_474),
.B(n_446),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_L g525 ( 
.A1(n_456),
.A2(n_178),
.B(n_41),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_485),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_457),
.A2(n_34),
.B(n_42),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_467),
.A2(n_45),
.B(n_46),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_490),
.A2(n_48),
.B(n_49),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_474),
.B(n_177),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_501),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_486),
.B(n_487),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_459),
.A2(n_50),
.B(n_60),
.Y(n_533)
);

NAND2x1_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_62),
.Y(n_534)
);

AOI21x1_ASAP7_75t_SL g535 ( 
.A1(n_508),
.A2(n_63),
.B(n_65),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_462),
.A2(n_69),
.B(n_70),
.Y(n_536)
);

NAND2x1_ASAP7_75t_L g537 ( 
.A(n_506),
.B(n_176),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_446),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_446),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_492),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_478),
.B(n_482),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_493),
.Y(n_542)
);

AOI211x1_ASAP7_75t_L g543 ( 
.A1(n_510),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_464),
.A2(n_496),
.B(n_458),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_499),
.B(n_75),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_447),
.A2(n_76),
.B(n_77),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_492),
.Y(n_547)
);

OAI21x1_ASAP7_75t_SL g548 ( 
.A1(n_511),
.A2(n_78),
.B(n_81),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_480),
.A2(n_82),
.B(n_84),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_494),
.Y(n_550)
);

O2A1O1Ixp5_ASAP7_75t_L g551 ( 
.A1(n_454),
.A2(n_85),
.B(n_86),
.C(n_87),
.Y(n_551)
);

AO31x2_ASAP7_75t_L g552 ( 
.A1(n_471),
.A2(n_88),
.A3(n_89),
.B(n_90),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_502),
.B(n_102),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_L g554 ( 
.A(n_504),
.B(n_172),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_470),
.B(n_104),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_491),
.A2(n_107),
.B(n_108),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_484),
.B(n_109),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_448),
.A2(n_110),
.B(n_111),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_498),
.B(n_113),
.Y(n_559)
);

AOI211x1_ASAP7_75t_L g560 ( 
.A1(n_510),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_560)
);

A2O1A1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_489),
.A2(n_120),
.B(n_123),
.C(n_124),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_445),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_495),
.A2(n_125),
.B(n_126),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_481),
.A2(n_127),
.B(n_132),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_449),
.A2(n_134),
.B(n_137),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_468),
.B(n_138),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_479),
.A2(n_140),
.B(n_144),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_505),
.B(n_145),
.Y(n_569)
);

A2O1A1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_497),
.A2(n_146),
.B(n_147),
.C(n_148),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_466),
.A2(n_150),
.B(n_151),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_503),
.Y(n_572)
);

NAND2x1p5_ASAP7_75t_L g573 ( 
.A(n_472),
.B(n_157),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_514),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_450),
.A2(n_161),
.B(n_162),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_572),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_538),
.B(n_476),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_539),
.Y(n_578)
);

AOI21x1_ASAP7_75t_L g579 ( 
.A1(n_569),
.A2(n_475),
.B(n_513),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

INVx8_ASAP7_75t_L g581 ( 
.A(n_545),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_541),
.B(n_463),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_532),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_569),
.A2(n_460),
.B(n_465),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_531),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_519),
.A2(n_517),
.B(n_544),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_520),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_550),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_522),
.A2(n_507),
.B(n_512),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_526),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_527),
.A2(n_461),
.B(n_483),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_562),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_536),
.A2(n_515),
.B(n_509),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_542),
.Y(n_595)
);

OR2x6_ASAP7_75t_L g596 ( 
.A(n_538),
.B(n_515),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_567),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_540),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_553),
.B(n_500),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_538),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_528),
.A2(n_163),
.B(n_166),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_552),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_524),
.B(n_168),
.Y(n_603)
);

OAI21x1_ASAP7_75t_L g604 ( 
.A1(n_571),
.A2(n_169),
.B(n_170),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_518),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_518),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_558),
.A2(n_533),
.B(n_535),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_574),
.B(n_559),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_552),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_563),
.A2(n_523),
.B(n_549),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_518),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_556),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_SL g615 ( 
.A1(n_557),
.A2(n_561),
.B(n_570),
.C(n_525),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_540),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_530),
.B(n_566),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_547),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_547),
.A2(n_566),
.B1(n_560),
.B2(n_543),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_547),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_551),
.A2(n_516),
.B(n_564),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_555),
.B(n_566),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_554),
.B(n_543),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_573),
.Y(n_624)
);

AO21x2_ASAP7_75t_L g625 ( 
.A1(n_525),
.A2(n_521),
.B(n_554),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_580),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_585),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_576),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_577),
.A2(n_565),
.B1(n_548),
.B2(n_529),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_588),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_587),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_592),
.Y(n_633)
);

OAI321xp33_ASAP7_75t_L g634 ( 
.A1(n_599),
.A2(n_560),
.A3(n_546),
.B1(n_575),
.B2(n_534),
.C(n_537),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_583),
.B(n_568),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_593),
.B(n_581),
.Y(n_636)
);

AO21x2_ASAP7_75t_L g637 ( 
.A1(n_602),
.A2(n_611),
.B(n_609),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_582),
.B(n_593),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_577),
.B(n_596),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_587),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_590),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_590),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_581),
.A2(n_603),
.B1(n_622),
.B2(n_617),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_595),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_618),
.B(n_596),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_618),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_595),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_602),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_581),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_606),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_609),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_608),
.A2(n_586),
.B(n_612),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_578),
.B(n_606),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_615),
.A2(n_584),
.B(n_621),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_600),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_611),
.Y(n_656)
);

O2A1O1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_615),
.A2(n_623),
.B(n_619),
.C(n_597),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_622),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_594),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_610),
.A2(n_603),
.B1(n_622),
.B2(n_617),
.Y(n_660)
);

OA21x2_ASAP7_75t_L g661 ( 
.A1(n_614),
.A2(n_589),
.B(n_579),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_SL g662 ( 
.A1(n_622),
.A2(n_625),
.B1(n_624),
.B2(n_598),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_600),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_605),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_614),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_613),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_622),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_601),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_591),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_592),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_591),
.Y(n_671)
);

NAND2x1_ASAP7_75t_L g672 ( 
.A(n_658),
.B(n_591),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_658),
.B(n_598),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_665),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_626),
.B(n_620),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_627),
.B(n_616),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_665),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_639),
.B(n_607),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_638),
.B(n_619),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_653),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_648),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_648),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_658),
.B(n_596),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_651),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_639),
.B(n_650),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_651),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_656),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_667),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_667),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_667),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_638),
.B(n_607),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_650),
.B(n_625),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_659),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_653),
.B(n_645),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_655),
.B(n_624),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_645),
.B(n_604),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_663),
.B(n_666),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_664),
.B(n_645),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_628),
.B(n_629),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_628),
.B(n_629),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_646),
.B(n_631),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_669),
.B(n_671),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_632),
.B(n_641),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_646),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_640),
.B(n_647),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_637),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_637),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_637),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_636),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_635),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_642),
.B(n_644),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_667),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_661),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_667),
.B(n_660),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_643),
.B(n_657),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_649),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_661),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_649),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_662),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_680),
.B(n_670),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_710),
.B(n_659),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_715),
.B(n_649),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_697),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_697),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_703),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_701),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_709),
.B(n_633),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_674),
.Y(n_729)
);

BUFx2_ASAP7_75t_L g730 ( 
.A(n_704),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_691),
.B(n_694),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_674),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_677),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_677),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_681),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_675),
.B(n_633),
.Y(n_736)
);

NAND2x1_ASAP7_75t_L g737 ( 
.A(n_673),
.B(n_654),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_685),
.B(n_652),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_675),
.B(n_649),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_685),
.B(n_652),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_703),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_705),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_692),
.B(n_668),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_681),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_676),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_686),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_705),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_686),
.Y(n_748)
);

AND2x4_ASAP7_75t_SL g749 ( 
.A(n_688),
.B(n_649),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_711),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_692),
.B(n_668),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_676),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_698),
.B(n_630),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_687),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_698),
.B(n_634),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_711),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_695),
.B(n_678),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_695),
.B(n_678),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_699),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_690),
.B(n_716),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_679),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_699),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_700),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_729),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_745),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_738),
.B(n_693),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_729),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_732),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_752),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_726),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_760),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_732),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_741),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_727),
.B(n_679),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_731),
.B(n_724),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_725),
.B(n_715),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_742),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_747),
.B(n_704),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_733),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_743),
.B(n_693),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_750),
.Y(n_781)
);

AND2x4_ASAP7_75t_SL g782 ( 
.A(n_761),
.B(n_688),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_756),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_730),
.B(n_696),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_760),
.B(n_723),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_759),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_757),
.B(n_718),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_721),
.B(n_673),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_762),
.Y(n_789)
);

INVxp67_ASAP7_75t_R g790 ( 
.A(n_755),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_738),
.B(n_713),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_740),
.B(n_713),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_758),
.B(n_714),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_728),
.B(n_690),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_740),
.B(n_719),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_721),
.Y(n_796)
);

O2A1O1Ixp5_ASAP7_75t_L g797 ( 
.A1(n_785),
.A2(n_723),
.B(n_737),
.C(n_755),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_765),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_769),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_786),
.Y(n_800)
);

AOI21xp33_ASAP7_75t_SL g801 ( 
.A1(n_778),
.A2(n_736),
.B(n_739),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_793),
.B(n_743),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_784),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_796),
.B(n_716),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_789),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_770),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_773),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_766),
.B(n_751),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_777),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_771),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_781),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_766),
.B(n_751),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_764),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_764),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_767),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_783),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_767),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_813),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_798),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_810),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_803),
.A2(n_774),
.B1(n_776),
.B2(n_785),
.Y(n_821)
);

OAI32xp33_ASAP7_75t_L g822 ( 
.A1(n_803),
.A2(n_788),
.A3(n_775),
.B1(n_787),
.B2(n_780),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_801),
.B(n_794),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_802),
.B(n_792),
.Y(n_824)
);

AOI21xp33_ASAP7_75t_SL g825 ( 
.A1(n_799),
.A2(n_788),
.B(n_792),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_800),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_797),
.B(n_791),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_808),
.B(n_791),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_812),
.B(n_795),
.Y(n_829)
);

INVx3_ASAP7_75t_SL g830 ( 
.A(n_805),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_821),
.B(n_827),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_830),
.B(n_804),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_823),
.A2(n_797),
.B(n_804),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_820),
.B(n_795),
.Y(n_834)
);

OAI221xp5_ASAP7_75t_L g835 ( 
.A1(n_825),
.A2(n_811),
.B1(n_816),
.B2(n_806),
.C(n_807),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_826),
.Y(n_836)
);

NAND2x1_ASAP7_75t_L g837 ( 
.A(n_819),
.B(n_809),
.Y(n_837)
);

OA21x2_ASAP7_75t_L g838 ( 
.A1(n_818),
.A2(n_815),
.B(n_814),
.Y(n_838)
);

A2O1A1O1Ixp25_ASAP7_75t_L g839 ( 
.A1(n_831),
.A2(n_835),
.B(n_833),
.C(n_832),
.D(n_836),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_837),
.B(n_824),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_834),
.B(n_822),
.Y(n_841)
);

AOI221xp5_ASAP7_75t_L g842 ( 
.A1(n_838),
.A2(n_825),
.B1(n_817),
.B2(n_829),
.C(n_828),
.Y(n_842)
);

NAND4xp25_ASAP7_75t_L g843 ( 
.A(n_838),
.B(n_753),
.C(n_722),
.D(n_780),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_831),
.A2(n_790),
.B1(n_720),
.B2(n_714),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_836),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_839),
.B(n_722),
.C(n_753),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_841),
.A2(n_782),
.B(n_720),
.Y(n_847)
);

NAND3xp33_ASAP7_75t_L g848 ( 
.A(n_842),
.B(n_672),
.C(n_815),
.Y(n_848)
);

NOR4xp25_ASAP7_75t_L g849 ( 
.A(n_845),
.B(n_814),
.C(n_813),
.D(n_779),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_840),
.B(n_782),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_844),
.B(n_749),
.Y(n_851)
);

NOR3xp33_ASAP7_75t_SL g852 ( 
.A(n_850),
.B(n_846),
.C(n_848),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_847),
.B(n_843),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_851),
.Y(n_854)
);

NAND4xp75_ASAP7_75t_L g855 ( 
.A(n_849),
.B(n_689),
.C(n_712),
.D(n_763),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_R g856 ( 
.A(n_854),
.B(n_690),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_852),
.Y(n_857)
);

NOR3xp33_ASAP7_75t_L g858 ( 
.A(n_853),
.B(n_672),
.C(n_712),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_855),
.Y(n_859)
);

XOR2x2_ASAP7_75t_L g860 ( 
.A(n_857),
.B(n_683),
.Y(n_860)
);

AND3x4_ASAP7_75t_L g861 ( 
.A(n_858),
.B(n_683),
.C(n_673),
.Y(n_861)
);

INVxp33_ASAP7_75t_L g862 ( 
.A(n_856),
.Y(n_862)
);

NOR2x1_ASAP7_75t_L g863 ( 
.A(n_859),
.B(n_683),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_857),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_859),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_864),
.A2(n_683),
.B1(n_673),
.B2(n_689),
.Y(n_866)
);

AOI222xp33_ASAP7_75t_L g867 ( 
.A1(n_865),
.A2(n_779),
.B1(n_772),
.B2(n_768),
.C1(n_734),
.C2(n_733),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_862),
.B(n_772),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_863),
.B(n_749),
.Y(n_869)
);

XOR2xp5_ASAP7_75t_L g870 ( 
.A(n_860),
.B(n_688),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_861),
.B(n_768),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_864),
.B(n_734),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_864),
.A2(n_719),
.B(n_717),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_868),
.A2(n_717),
.B(n_748),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_872),
.B(n_688),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_872),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_870),
.Y(n_877)
);

XNOR2xp5_ASAP7_75t_L g878 ( 
.A(n_866),
.B(n_700),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_R g879 ( 
.A(n_869),
.B(n_688),
.Y(n_879)
);

XNOR2xp5_ASAP7_75t_L g880 ( 
.A(n_877),
.B(n_876),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_879),
.B(n_873),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_875),
.A2(n_871),
.B1(n_867),
.B2(n_754),
.Y(n_882)
);

OAI22x1_ASAP7_75t_L g883 ( 
.A1(n_878),
.A2(n_754),
.B1(n_748),
.B2(n_746),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_879),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_884),
.B(n_874),
.Y(n_885)
);

OA22x2_ASAP7_75t_L g886 ( 
.A1(n_880),
.A2(n_682),
.B1(n_684),
.B2(n_707),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_881),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_SL g888 ( 
.A1(n_882),
.A2(n_682),
.B1(n_684),
.B2(n_707),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_883),
.Y(n_889)
);

INVxp67_ASAP7_75t_SL g890 ( 
.A(n_887),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_885),
.A2(n_889),
.B(n_888),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_886),
.A2(n_746),
.B(n_744),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_890),
.A2(n_744),
.B(n_735),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_891),
.B(n_735),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_894),
.A2(n_892),
.B1(n_706),
.B2(n_708),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_893),
.B(n_702),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_895),
.A2(n_896),
.B(n_706),
.Y(n_897)
);


endmodule