module real_aes_4510_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_936;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_926;
wire n_922;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_0), .A2(n_41), .B1(n_697), .B2(n_700), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_1), .A2(n_102), .B1(n_335), .B2(n_388), .Y(n_547) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_2), .Y(n_655) );
AND2x4_ASAP7_75t_L g670 ( .A(n_2), .B(n_671), .Y(n_670) );
AND2x4_ASAP7_75t_L g680 ( .A(n_2), .B(n_240), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_3), .A2(n_204), .B1(n_383), .B2(n_386), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_4), .A2(n_150), .B1(n_525), .B2(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g304 ( .A(n_5), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_6), .A2(n_50), .B1(n_347), .B2(n_436), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_7), .A2(n_30), .B1(n_368), .B2(n_370), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_8), .A2(n_247), .B1(n_293), .B2(n_475), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_9), .B(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_10), .A2(n_21), .B1(n_447), .B2(n_534), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_11), .A2(n_189), .B1(n_357), .B2(n_436), .Y(n_900) );
AOI21xp33_ASAP7_75t_L g495 ( .A1(n_12), .A2(n_418), .B(n_496), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_13), .A2(n_99), .B1(n_442), .B2(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_14), .A2(n_170), .B1(n_408), .B2(n_409), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_15), .A2(n_109), .B1(n_385), .B2(n_546), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_16), .A2(n_633), .B(n_634), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_17), .A2(n_220), .B1(n_357), .B2(n_379), .Y(n_378) );
XOR2xp5_ASAP7_75t_L g255 ( .A(n_18), .B(n_256), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_18), .A2(n_69), .B1(n_690), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_19), .A2(n_146), .B1(n_402), .B2(n_403), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_20), .A2(n_128), .B1(n_375), .B2(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g677 ( .A(n_22), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_23), .A2(n_195), .B1(n_593), .B2(n_637), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g549 ( .A1(n_24), .A2(n_40), .B1(n_460), .B2(n_550), .C(n_551), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_25), .A2(n_68), .B1(n_683), .B2(n_713), .Y(n_763) );
INVx1_ASAP7_75t_SL g746 ( .A(n_26), .Y(n_746) );
INVx1_ASAP7_75t_L g888 ( .A(n_27), .Y(n_888) );
INVx1_ASAP7_75t_L g552 ( .A(n_28), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_29), .A2(n_163), .B1(n_445), .B2(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g279 ( .A(n_31), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_31), .B(n_192), .Y(n_326) );
INVxp67_ASAP7_75t_L g355 ( .A(n_31), .Y(n_355) );
OA22x2_ASAP7_75t_L g395 ( .A1(n_32), .A2(n_396), .B1(n_420), .B2(n_421), .Y(n_395) );
INVx1_ASAP7_75t_L g421 ( .A(n_32), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_32), .A2(n_73), .B1(n_667), .B2(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_33), .A2(n_194), .B1(n_415), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_34), .A2(n_108), .B1(n_386), .B2(n_536), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_35), .A2(n_47), .B1(n_402), .B2(n_403), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_36), .B(n_372), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_37), .A2(n_91), .B1(n_287), .B2(n_936), .Y(n_935) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_38), .B(n_264), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_39), .A2(n_216), .B1(n_447), .B2(n_534), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_42), .A2(n_239), .B1(n_357), .B2(n_379), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_43), .A2(n_214), .B1(n_385), .B2(n_386), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_44), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_45), .A2(n_248), .B1(n_679), .B2(n_714), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_46), .A2(n_86), .B1(n_436), .B2(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g517 ( .A(n_48), .Y(n_517) );
INVxp67_ASAP7_75t_R g681 ( .A(n_49), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_51), .A2(n_232), .B1(n_332), .B2(n_335), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_52), .A2(n_124), .B1(n_447), .B2(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_53), .A2(n_153), .B1(n_452), .B2(n_898), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_54), .A2(n_100), .B1(n_377), .B2(n_902), .Y(n_901) );
INVx2_ASAP7_75t_L g653 ( .A(n_55), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_56), .A2(n_89), .B1(n_287), .B2(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g513 ( .A(n_57), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_58), .A2(n_119), .B1(n_287), .B2(n_293), .Y(n_286) );
INVx1_ASAP7_75t_L g669 ( .A(n_59), .Y(n_669) );
AND2x4_ASAP7_75t_L g674 ( .A(n_59), .B(n_653), .Y(n_674) );
INVx1_ASAP7_75t_SL g691 ( .A(n_59), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_60), .A2(n_182), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_61), .A2(n_885), .B(n_887), .Y(n_884) );
INVx1_ASAP7_75t_L g466 ( .A(n_62), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_63), .A2(n_159), .B1(n_568), .B2(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g364 ( .A(n_64), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_64), .A2(n_186), .B1(n_690), .B2(n_704), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_65), .A2(n_226), .B1(n_332), .B2(n_335), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_66), .A2(n_168), .B1(n_923), .B2(n_926), .Y(n_922) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_67), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_70), .A2(n_178), .B1(n_335), .B2(n_388), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_71), .A2(n_244), .B1(n_282), .B2(n_293), .Y(n_469) );
INVx1_ASAP7_75t_L g919 ( .A(n_72), .Y(n_919) );
CKINVDCx16_ASAP7_75t_R g675 ( .A(n_74), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_75), .A2(n_156), .B1(n_667), .B2(n_765), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_76), .A2(n_155), .B1(n_382), .B2(n_383), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_77), .A2(n_123), .B1(n_382), .B2(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_78), .A2(n_215), .B1(n_405), .B2(n_406), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_79), .A2(n_238), .B1(n_287), .B2(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g265 ( .A(n_80), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_80), .B(n_191), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_81), .A2(n_167), .B1(n_587), .B2(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g318 ( .A(n_82), .Y(n_318) );
OAI22x1_ASAP7_75t_L g623 ( .A1(n_83), .A2(n_624), .B1(n_629), .B2(n_642), .Y(n_623) );
NAND5xp2_ASAP7_75t_SL g624 ( .A(n_83), .B(n_625), .C(n_626), .D(n_627), .E(n_628), .Y(n_624) );
AO22x1_ASAP7_75t_L g434 ( .A1(n_84), .A2(n_105), .B1(n_370), .B2(n_379), .Y(n_434) );
XNOR2x1_ASAP7_75t_L g489 ( .A(n_85), .B(n_490), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_87), .A2(n_141), .B1(n_614), .B2(n_616), .C(n_618), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_88), .B(n_460), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_90), .A2(n_134), .B1(n_411), .B2(n_419), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_92), .A2(n_242), .B1(n_399), .B2(n_400), .Y(n_398) );
INVx2_ASAP7_75t_R g507 ( .A(n_93), .Y(n_507) );
AOI221xp5_ASAP7_75t_SL g410 ( .A1(n_94), .A2(n_222), .B1(n_314), .B2(n_411), .C(n_412), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_95), .A2(n_116), .B1(n_345), .B2(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_96), .A2(n_140), .B1(n_472), .B2(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g692 ( .A(n_97), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_98), .A2(n_158), .B1(n_713), .B2(n_714), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_101), .A2(n_172), .B1(n_450), .B2(n_536), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_103), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_104), .A2(n_165), .B1(n_415), .B2(n_416), .C(n_417), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_106), .A2(n_218), .B1(n_400), .B2(n_405), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_107), .A2(n_433), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_110), .B(n_314), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_111), .A2(n_132), .B1(n_332), .B2(n_563), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_112), .A2(n_145), .B1(n_408), .B2(n_409), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_113), .A2(n_161), .B1(n_679), .B2(n_683), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_113), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_113), .A2(n_910), .B1(n_912), .B2(n_937), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_114), .A2(n_148), .B1(n_259), .B2(n_382), .Y(n_930) );
INVx1_ASAP7_75t_L g497 ( .A(n_115), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_117), .A2(n_225), .B1(n_287), .B2(n_452), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_118), .A2(n_173), .B1(n_335), .B2(n_534), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_120), .A2(n_205), .B1(n_382), .B2(n_454), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_121), .A2(n_133), .B1(n_338), .B2(n_340), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_122), .A2(n_184), .B1(n_377), .B2(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_125), .A2(n_157), .B1(n_345), .B2(n_347), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_126), .A2(n_162), .B1(n_471), .B2(n_472), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_127), .A2(n_231), .B1(n_399), .B2(n_411), .Y(n_501) );
INVx1_ASAP7_75t_L g635 ( .A(n_129), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_130), .A2(n_213), .B1(n_259), .B2(n_450), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_131), .A2(n_199), .B1(n_415), .B2(n_419), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_135), .A2(n_183), .B1(n_282), .B2(n_454), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_136), .A2(n_171), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_137), .A2(n_236), .B1(n_332), .B2(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_138), .A2(n_228), .B1(n_385), .B2(n_546), .Y(n_607) );
INVx1_ASAP7_75t_L g511 ( .A(n_139), .Y(n_511) );
INVx1_ASAP7_75t_L g695 ( .A(n_142), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_143), .A2(n_221), .B1(n_697), .B2(n_700), .Y(n_709) );
AO22x1_ASAP7_75t_L g417 ( .A1(n_144), .A2(n_212), .B1(n_418), .B2(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g693 ( .A(n_147), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_149), .A2(n_237), .B1(n_338), .B2(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_151), .A2(n_185), .B1(n_565), .B2(n_566), .Y(n_564) );
XNOR2x1_ASAP7_75t_L g456 ( .A(n_152), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g518 ( .A(n_154), .Y(n_518) );
XOR2xp5_ASAP7_75t_L g912 ( .A(n_160), .B(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_164), .A2(n_200), .B1(n_406), .B2(n_416), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_166), .A2(n_219), .B1(n_436), .B2(n_437), .Y(n_435) );
OA22x2_ASAP7_75t_L g269 ( .A1(n_169), .A2(n_192), .B1(n_264), .B2(n_268), .Y(n_269) );
INVx1_ASAP7_75t_L g300 ( .A(n_169), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_174), .A2(n_201), .B1(n_357), .B2(n_359), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_175), .A2(n_575), .B(n_578), .Y(n_574) );
AOI221x1_ASAP7_75t_L g917 ( .A1(n_176), .A2(n_209), .B1(n_577), .B2(n_641), .C(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_177), .A2(n_229), .B1(n_259), .B2(n_382), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_179), .A2(n_187), .B1(n_450), .B2(n_536), .Y(n_931) );
INVx1_ASAP7_75t_L g585 ( .A(n_180), .Y(n_585) );
INVx1_ASAP7_75t_L g581 ( .A(n_181), .Y(n_581) );
CKINVDCx6p67_ASAP7_75t_R g672 ( .A(n_188), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_190), .Y(n_427) );
INVx1_ASAP7_75t_L g281 ( .A(n_191), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_191), .B(n_298), .Y(n_329) );
OAI21xp33_ASAP7_75t_L g301 ( .A1(n_192), .A2(n_202), .B(n_302), .Y(n_301) );
AO22x2_ASAP7_75t_L g559 ( .A1(n_193), .A2(n_560), .B1(n_594), .B2(n_595), .Y(n_559) );
INVx1_ASAP7_75t_L g595 ( .A(n_193), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_196), .A2(n_208), .B1(n_667), .B2(n_716), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_197), .A2(n_206), .B1(n_441), .B2(n_442), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_198), .A2(n_224), .B1(n_450), .B2(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g267 ( .A(n_202), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_202), .B(n_233), .Y(n_327) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_203), .A2(n_314), .B(n_317), .Y(n_313) );
INVx1_ASAP7_75t_L g619 ( .A(n_207), .Y(n_619) );
INVx1_ASAP7_75t_L g747 ( .A(n_210), .Y(n_747) );
XNOR2x1_ASAP7_75t_L g602 ( .A(n_211), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g521 ( .A(n_217), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_223), .A2(n_227), .B1(n_571), .B2(n_572), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_230), .A2(n_235), .B1(n_259), .B2(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_233), .B(n_273), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_234), .A2(n_241), .B1(n_259), .B2(n_282), .Y(n_258) );
INVx1_ASAP7_75t_L g671 ( .A(n_240), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_243), .B(n_639), .Y(n_638) );
XNOR2x1_ASAP7_75t_L g540 ( .A(n_245), .B(n_541), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_246), .A2(n_431), .B(n_434), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_482), .B(n_648), .C(n_656), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_250), .A2(n_482), .B(n_649), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_423), .B1(n_480), .B2(n_481), .Y(n_250) );
INVx1_ASAP7_75t_L g480 ( .A(n_251), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_392), .B1(n_393), .B2(n_422), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g422 ( .A(n_253), .Y(n_422) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
XNOR2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_362), .Y(n_254) );
NAND4xp75_ASAP7_75t_L g256 ( .A(n_257), .B(n_303), .C(n_330), .D(n_343), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_286), .Y(n_257) );
BUFx3_ASAP7_75t_L g571 ( .A(n_259), .Y(n_571) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx8_ASAP7_75t_L g454 ( .A(n_260), .Y(n_454) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_270), .Y(n_260) );
AND2x4_ASAP7_75t_L g283 ( .A(n_261), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g309 ( .A(n_261), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g358 ( .A(n_261), .B(n_334), .Y(n_358) );
AND2x4_ASAP7_75t_L g399 ( .A(n_261), .B(n_270), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_261), .B(n_292), .Y(n_400) );
AND2x4_ASAP7_75t_L g415 ( .A(n_261), .B(n_334), .Y(n_415) );
AND2x2_ASAP7_75t_L g418 ( .A(n_261), .B(n_310), .Y(n_418) );
AND2x2_ASAP7_75t_L g473 ( .A(n_261), .B(n_270), .Y(n_473) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_269), .Y(n_261) );
INVx1_ASAP7_75t_L g290 ( .A(n_262), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
NAND2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g268 ( .A(n_264), .Y(n_268) );
INVx3_ASAP7_75t_L g273 ( .A(n_264), .Y(n_273) );
NAND2xp33_ASAP7_75t_L g280 ( .A(n_264), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g302 ( .A(n_264), .Y(n_302) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_264), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_265), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_267), .A2(n_302), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
AND2x2_ASAP7_75t_L g316 ( .A(n_269), .B(n_290), .Y(n_316) );
AND2x2_ASAP7_75t_L g353 ( .A(n_269), .B(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g339 ( .A(n_270), .B(n_289), .Y(n_339) );
AND2x4_ASAP7_75t_L g342 ( .A(n_270), .B(n_296), .Y(n_342) );
AND2x4_ASAP7_75t_L g405 ( .A(n_270), .B(n_289), .Y(n_405) );
AND2x4_ASAP7_75t_L g408 ( .A(n_270), .B(n_296), .Y(n_408) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .Y(n_270) );
OR2x2_ASAP7_75t_L g285 ( .A(n_271), .B(n_276), .Y(n_285) );
INVx2_ASAP7_75t_L g311 ( .A(n_271), .Y(n_311) );
AND2x4_ASAP7_75t_L g334 ( .A(n_271), .B(n_312), .Y(n_334) );
AND2x2_ASAP7_75t_L g350 ( .A(n_271), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_273), .B(n_279), .Y(n_278) );
INVxp67_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g328 ( .A(n_274), .B(n_297), .C(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
BUFx3_ASAP7_75t_L g572 ( .A(n_282), .Y(n_572) );
BUFx12f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_283), .Y(n_382) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_283), .Y(n_606) );
BUFx3_ASAP7_75t_L g898 ( .A(n_283), .Y(n_898) );
AND2x4_ASAP7_75t_L g406 ( .A(n_284), .B(n_289), .Y(n_406) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g292 ( .A(n_285), .Y(n_292) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_288), .Y(n_386) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_288), .Y(n_475) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
AND2x4_ASAP7_75t_L g333 ( .A(n_289), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g336 ( .A(n_289), .B(n_310), .Y(n_336) );
AND2x4_ASAP7_75t_L g402 ( .A(n_289), .B(n_334), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_289), .B(n_310), .Y(n_403) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x4_ASAP7_75t_L g295 ( .A(n_292), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g409 ( .A(n_292), .B(n_296), .Y(n_409) );
INVx5_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g383 ( .A(n_294), .Y(n_383) );
INVx1_ASAP7_75t_L g531 ( .A(n_294), .Y(n_531) );
INVx1_ASAP7_75t_L g936 ( .A(n_294), .Y(n_936) );
INVx6_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx12f_ASAP7_75t_L g452 ( .A(n_295), .Y(n_452) );
AND2x4_ASAP7_75t_L g361 ( .A(n_296), .B(n_310), .Y(n_361) );
AND2x4_ASAP7_75t_L g419 ( .A(n_296), .B(n_310), .Y(n_419) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OA21x2_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_313), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g577 ( .A(n_307), .Y(n_577) );
INVx2_ASAP7_75t_L g639 ( .A(n_307), .Y(n_639) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx3_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
BUFx3_ASAP7_75t_L g433 ( .A(n_309), .Y(n_433) );
AND2x4_ASAP7_75t_L g315 ( .A(n_310), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g373 ( .A(n_315), .Y(n_373) );
BUFx8_ASAP7_75t_SL g460 ( .A(n_315), .Y(n_460) );
INVx2_ASAP7_75t_L g615 ( .A(n_315), .Y(n_615) );
BUFx3_ASAP7_75t_L g902 ( .A(n_315), .Y(n_902) );
AND2x4_ASAP7_75t_L g346 ( .A(n_316), .B(n_334), .Y(n_346) );
AND2x4_ASAP7_75t_L g411 ( .A(n_316), .B(n_334), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_319), .B(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g370 ( .A(n_321), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_321), .B(n_413), .Y(n_412) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_321), .Y(n_467) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx3_ASAP7_75t_L g499 ( .A(n_322), .Y(n_499) );
AO21x2_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B(n_328), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_324), .B(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_325), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_337), .Y(n_330) );
BUFx12f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx3_ASAP7_75t_L g389 ( .A(n_333), .Y(n_389) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_333), .Y(n_534) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx5_ASAP7_75t_L g447 ( .A(n_336), .Y(n_447) );
BUFx3_ASAP7_75t_L g477 ( .A(n_336), .Y(n_477) );
BUFx2_ASAP7_75t_SL g568 ( .A(n_338), .Y(n_568) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_339), .Y(n_385) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_339), .Y(n_536) );
INVx4_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g391 ( .A(n_341), .Y(n_391) );
INVx4_ASAP7_75t_L g450 ( .A(n_341), .Y(n_450) );
INVx2_ASAP7_75t_L g471 ( .A(n_341), .Y(n_471) );
INVx2_ASAP7_75t_SL g546 ( .A(n_341), .Y(n_546) );
INVx8_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_356), .Y(n_343) );
BUFx2_ASAP7_75t_L g590 ( .A(n_345), .Y(n_590) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g376 ( .A(n_346), .Y(n_376) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_346), .Y(n_436) );
BUFx3_ASAP7_75t_L g633 ( .A(n_346), .Y(n_633) );
INVx2_ASAP7_75t_L g889 ( .A(n_347), .Y(n_889) );
INVx4_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g580 ( .A(n_348), .Y(n_580) );
INVx2_ASAP7_75t_L g609 ( .A(n_348), .Y(n_609) );
INVx2_ASAP7_75t_L g637 ( .A(n_348), .Y(n_637) );
INVx3_ASAP7_75t_L g926 ( .A(n_348), .Y(n_926) );
INVx5_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g379 ( .A(n_349), .Y(n_379) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_349), .Y(n_525) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_353), .Y(n_349) );
AND2x2_ASAP7_75t_L g416 ( .A(n_350), .B(n_353), .Y(n_416) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g439 ( .A(n_358), .Y(n_439) );
BUFx3_ASAP7_75t_L g593 ( .A(n_358), .Y(n_593) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx3_ASAP7_75t_L g377 ( .A(n_360), .Y(n_377) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_361), .Y(n_442) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_361), .Y(n_463) );
XNOR2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_364), .Y(n_363) );
NOR2x1_ASAP7_75t_L g365 ( .A(n_366), .B(n_380), .Y(n_365) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_367), .B(n_371), .C(n_374), .D(n_378), .Y(n_366) );
INVx2_ASAP7_75t_L g886 ( .A(n_368), .Y(n_886) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g523 ( .A(n_369), .Y(n_523) );
INVx2_ASAP7_75t_L g550 ( .A(n_369), .Y(n_550) );
INVx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g441 ( .A(n_373), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_373), .A2(n_517), .B1(n_518), .B2(n_519), .Y(n_516) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND4xp25_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .C(n_387), .D(n_390), .Y(n_380) );
BUFx12f_ASAP7_75t_L g449 ( .A(n_385), .Y(n_449) );
BUFx3_ASAP7_75t_L g565 ( .A(n_386), .Y(n_565) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g446 ( .A(n_389), .Y(n_446) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
BUFx4_ASAP7_75t_R g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g420 ( .A(n_396), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_410), .C(n_414), .Y(n_396) );
AND4x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_401), .C(n_404), .D(n_407), .Y(n_397) );
INVx2_ASAP7_75t_L g617 ( .A(n_418), .Y(n_617) );
INVx1_ASAP7_75t_L g481 ( .A(n_423), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_455), .B1(n_478), .B2(n_479), .Y(n_423) );
INVx1_ASAP7_75t_L g478 ( .A(n_424), .Y(n_478) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
XNOR2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NOR2xp67_ASAP7_75t_L g428 ( .A(n_429), .B(n_443), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_435), .C(n_440), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx4_ASAP7_75t_L g512 ( .A(n_436), .Y(n_512) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g515 ( .A(n_438), .Y(n_515) );
INVx2_ASAP7_75t_L g555 ( .A(n_438), .Y(n_555) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g925 ( .A(n_439), .Y(n_925) );
INVx4_ASAP7_75t_L g519 ( .A(n_442), .Y(n_519) );
BUFx3_ASAP7_75t_L g588 ( .A(n_442), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g443 ( .A(n_444), .B(n_448), .C(n_451), .D(n_453), .Y(n_443) );
BUFx4f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g563 ( .A(n_447), .Y(n_563) );
BUFx3_ASAP7_75t_L g566 ( .A(n_452), .Y(n_566) );
INVx2_ASAP7_75t_L g479 ( .A(n_455), .Y(n_479) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_468), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .C(n_462), .D(n_464), .Y(n_458) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_460), .Y(n_587) );
BUFx3_ASAP7_75t_L g921 ( .A(n_463), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_467), .B(n_619), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .C(n_474), .D(n_476), .Y(n_468) );
BUFx2_ASAP7_75t_SL g569 ( .A(n_471), .Y(n_569) );
BUFx4f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
XNOR2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_557), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI22x1_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_538), .B2(n_556), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AO22x2_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_505), .B1(n_506), .B2(n_537), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g537 ( .A(n_489), .Y(n_537) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_491), .B(n_500), .Y(n_490) );
NAND4xp25_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .C(n_494), .D(n_495), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g526 ( .A(n_498), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_498), .B(n_635), .Y(n_634) );
INVx4_ASAP7_75t_L g891 ( .A(n_498), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_498), .B(n_919), .Y(n_918) );
INVx4_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g584 ( .A(n_499), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .C(n_503), .D(n_504), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
XNOR2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_527), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .C(n_520), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_510) );
INVxp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI21xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_524), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND2xp33_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
INVx1_ASAP7_75t_L g556 ( .A(n_538), .Y(n_556) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_548), .Y(n_541) );
NAND4xp25_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .C(n_545), .D(n_547), .Y(n_542) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .C(n_554), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_596), .B2(n_597), .Y(n_557) );
INVx4_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g594 ( .A(n_560), .Y(n_594) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_573), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .C(n_567), .D(n_570), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_586), .C(n_589), .Y(n_573) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B1(n_582), .B2(n_585), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx4_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI22x1_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_621), .B1(n_646), .B2(n_647), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g647 ( .A(n_600), .Y(n_647) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_611), .Y(n_603) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .C(n_608), .D(n_610), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .C(n_620), .Y(n_611) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_SL g641 ( .A(n_615), .Y(n_641) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g646 ( .A(n_621), .Y(n_646) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g643 ( .A(n_625), .B(n_626), .C(n_628), .D(n_638), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_627), .B(n_640), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_638), .C(n_640), .Y(n_629) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g644 ( .A(n_631), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
BUFx4_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .C(n_655), .Y(n_650) );
AND2x2_ASAP7_75t_L g906 ( .A(n_651), .B(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g911 ( .A(n_651), .B(n_908), .Y(n_911) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OA21x2_ASAP7_75t_L g938 ( .A1(n_652), .A2(n_691), .B(n_939), .Y(n_938) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g668 ( .A(n_653), .B(n_669), .Y(n_668) );
AND3x4_ASAP7_75t_L g690 ( .A(n_653), .B(n_670), .C(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g907 ( .A(n_654), .B(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_655), .Y(n_908) );
OAI221xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_877), .B1(n_879), .B2(n_904), .C(n_909), .Y(n_656) );
AND5x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_821), .C(n_838), .D(n_847), .E(n_867), .Y(n_657) );
AOI222xp33_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_744), .B1(n_758), .B2(n_767), .C1(n_800), .C2(n_820), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_738), .B1(n_744), .B2(n_749), .C(n_754), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_717), .C(n_730), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_684), .Y(n_661) );
AND2x2_ASAP7_75t_L g872 ( .A(n_662), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_663), .A2(n_718), .B1(n_723), .B2(n_727), .C(n_729), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_663), .B(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g817 ( .A(n_663), .Y(n_817) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g725 ( .A(n_664), .Y(n_725) );
AND2x2_ASAP7_75t_L g741 ( .A(n_664), .B(n_739), .Y(n_741) );
OR2x2_ASAP7_75t_L g775 ( .A(n_664), .B(n_733), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_664), .B(n_687), .Y(n_777) );
AND2x2_ASAP7_75t_L g789 ( .A(n_664), .B(n_733), .Y(n_789) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_676), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_672), .B1(n_673), .B2(n_675), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_666), .A2(n_673), .B1(n_746), .B2(n_747), .C(n_748), .Y(n_745) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
AND2x4_ASAP7_75t_L g679 ( .A(n_668), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g700 ( .A(n_668), .B(n_680), .Y(n_700) );
AND2x2_ASAP7_75t_L g713 ( .A(n_668), .B(n_680), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_670), .B(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g704 ( .A(n_670), .B(n_674), .Y(n_704) );
AND2x4_ASAP7_75t_L g716 ( .A(n_670), .B(n_674), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_673), .A2(n_689), .B1(n_692), .B2(n_693), .Y(n_688) );
AND2x4_ASAP7_75t_L g683 ( .A(n_674), .B(n_680), .Y(n_683) );
AND2x2_ASAP7_75t_L g697 ( .A(n_674), .B(n_680), .Y(n_697) );
AND2x2_ASAP7_75t_L g714 ( .A(n_674), .B(n_680), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_681), .B2(n_682), .Y(n_676) );
INVx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g939 ( .A(n_680), .Y(n_939) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx2_ASAP7_75t_L g878 ( .A(n_683), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_684), .B(n_783), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_701), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_685), .B(n_720), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_685), .B(n_783), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_685), .B(n_762), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_685), .B(n_719), .Y(n_876) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
CKINVDCx6p67_ASAP7_75t_R g726 ( .A(n_687), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_687), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g770 ( .A(n_687), .B(n_743), .Y(n_770) );
AND2x2_ASAP7_75t_L g780 ( .A(n_687), .B(n_725), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_687), .B(n_725), .Y(n_808) );
AND2x2_ASAP7_75t_L g827 ( .A(n_687), .B(n_793), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_687), .B(n_722), .Y(n_863) );
OR2x6_ASAP7_75t_SL g687 ( .A(n_688), .B(n_694), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_698), .B2(n_699), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g782 ( .A(n_701), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_701), .B(n_719), .Y(n_842) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_706), .Y(n_701) );
CKINVDCx6p67_ASAP7_75t_R g722 ( .A(n_702), .Y(n_722) );
INVx1_ASAP7_75t_L g753 ( .A(n_702), .Y(n_753) );
OR2x2_ASAP7_75t_L g757 ( .A(n_702), .B(n_707), .Y(n_757) );
OAI32xp33_ASAP7_75t_L g773 ( .A1(n_702), .A2(n_757), .A3(n_774), .B1(n_775), .B2(n_776), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_702), .B(n_707), .Y(n_791) );
AND2x2_ASAP7_75t_L g793 ( .A(n_702), .B(n_720), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_702), .B(n_721), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_702), .B(n_743), .Y(n_871) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
INVx2_ASAP7_75t_SL g766 ( .A(n_704), .Y(n_766) );
OR2x2_ASAP7_75t_L g774 ( .A(n_706), .B(n_720), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_706), .B(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g824 ( .A(n_706), .B(n_722), .Y(n_824) );
INVx1_ASAP7_75t_L g862 ( .A(n_706), .Y(n_862) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_707), .Y(n_721) );
AND2x2_ASAP7_75t_L g813 ( .A(n_707), .B(n_711), .Y(n_813) );
AND2x4_ASAP7_75t_SL g707 ( .A(n_708), .B(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g728 ( .A(n_710), .Y(n_728) );
AND2x2_ASAP7_75t_L g737 ( .A(n_710), .B(n_722), .Y(n_737) );
AND2x2_ASAP7_75t_L g743 ( .A(n_710), .B(n_721), .Y(n_743) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g720 ( .A(n_711), .B(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .Y(n_711) );
OAI211xp5_ASAP7_75t_SL g825 ( .A1(n_718), .A2(n_776), .B(n_826), .C(n_828), .Y(n_825) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_SL g719 ( .A(n_720), .B(n_722), .Y(n_719) );
AND2x2_ASAP7_75t_L g785 ( .A(n_720), .B(n_786), .Y(n_785) );
OAI21xp33_ASAP7_75t_L g815 ( .A1(n_720), .A2(n_724), .B(n_737), .Y(n_815) );
AND2x2_ASAP7_75t_L g854 ( .A(n_720), .B(n_830), .Y(n_854) );
OAI222xp33_ASAP7_75t_L g730 ( .A1(n_721), .A2(n_731), .B1(n_736), .B2(n_738), .C1(n_740), .C2(n_742), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_721), .B(n_752), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_721), .A2(n_789), .B1(n_802), .B2(n_803), .Y(n_801) );
AND2x2_ASAP7_75t_L g786 ( .A(n_722), .B(n_726), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_722), .B(n_743), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_722), .B(n_813), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_722), .B(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_722), .B(n_770), .Y(n_849) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_724), .B(n_759), .Y(n_790) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AND2x2_ASAP7_75t_L g732 ( .A(n_725), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g755 ( .A(n_725), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_725), .B(n_781), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_725), .B(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_725), .B(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_726), .B(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_726), .B(n_751), .Y(n_750) );
NOR2x1p5_ASAP7_75t_L g756 ( .A(n_726), .B(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_726), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g805 ( .A(n_726), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_726), .B(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g830 ( .A(n_726), .B(n_752), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_726), .B(n_741), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_726), .B(n_775), .Y(n_846) );
INVx1_ASAP7_75t_L g807 ( .A(n_727), .Y(n_807) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVxp67_ASAP7_75t_L g868 ( .A(n_731), .Y(n_868) );
INVx1_ASAP7_75t_L g814 ( .A(n_732), .Y(n_814) );
INVx2_ASAP7_75t_L g739 ( .A(n_733), .Y(n_739) );
AND2x2_ASAP7_75t_L g852 ( .A(n_733), .B(n_762), .Y(n_852) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_737), .A2(n_793), .B1(n_794), .B2(n_796), .C(n_797), .Y(n_792) );
AOI211xp5_ASAP7_75t_L g809 ( .A1(n_737), .A2(n_810), .B(n_811), .C(n_818), .Y(n_809) );
OAI211xp5_ASAP7_75t_SL g767 ( .A1(n_738), .A2(n_768), .B(n_771), .C(n_792), .Y(n_767) );
INVx3_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g781 ( .A(n_739), .B(n_762), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_739), .B(n_761), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_739), .B(n_762), .Y(n_874) );
OAI221xp5_ASAP7_75t_L g855 ( .A1(n_740), .A2(n_856), .B1(n_858), .B2(n_860), .C(n_864), .Y(n_855) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
BUFx3_ASAP7_75t_L g820 ( .A(n_745), .Y(n_820) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g769 ( .A(n_752), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx3_ASAP7_75t_L g772 ( .A(n_758), .Y(n_772) );
OAI311xp33_ASAP7_75t_L g811 ( .A1(n_758), .A2(n_812), .A3(n_814), .B1(n_815), .C1(n_816), .Y(n_811) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_760), .B(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_761), .B(n_785), .Y(n_784) );
INVx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g795 ( .A(n_762), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_762), .B(n_789), .Y(n_799) );
AND2x2_ASAP7_75t_L g836 ( .A(n_762), .B(n_837), .Y(n_836) );
AND2x4_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AOI211xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B(n_778), .C(n_787), .Y(n_771) );
INVx1_ASAP7_75t_L g837 ( .A(n_775), .Y(n_837) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OAI221xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_781), .B1(n_782), .B2(n_783), .C(n_784), .Y(n_778) );
INVx1_ASAP7_75t_L g803 ( .A(n_781), .Y(n_803) );
OAI221xp5_ASAP7_75t_SL g800 ( .A1(n_783), .A2(n_801), .B1(n_804), .B2(n_806), .C(n_809), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_786), .B(n_813), .Y(n_866) );
AOI21xp33_ASAP7_75t_SL g787 ( .A1(n_788), .A2(n_790), .B(n_791), .Y(n_787) );
AOI211xp5_ASAP7_75t_SL g847 ( .A1(n_789), .A2(n_848), .B(n_850), .C(n_855), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_791), .B(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g869 ( .A(n_791), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_793), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g819 ( .A(n_793), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_793), .B(n_857), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g802 ( .A(n_798), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g821 ( .A1(n_803), .A2(n_810), .B1(n_822), .B2(n_825), .C(n_831), .Y(n_821) );
CKINVDCx14_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
AND2x2_ASAP7_75t_L g829 ( .A(n_813), .B(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g834 ( .A(n_813), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_817), .B(n_827), .Y(n_826) );
AOI322xp5_ASAP7_75t_L g867 ( .A1(n_820), .A2(n_852), .A3(n_868), .B1(n_869), .B2(n_870), .C1(n_872), .C2(n_875), .Y(n_867) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_835), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_837), .B(n_859), .Y(n_858) );
OAI21xp33_ASAP7_75t_L g864 ( .A1(n_837), .A2(n_852), .B(n_865), .Y(n_864) );
AOI211xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_841), .B(n_843), .C(n_844), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVxp67_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_853), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_878), .Y(n_877) );
INVxp67_ASAP7_75t_SL g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_SL g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
XNOR2x1_ASAP7_75t_L g882 ( .A(n_883), .B(n_903), .Y(n_882) );
NAND4xp75_ASAP7_75t_L g883 ( .A(n_884), .B(n_892), .C(n_895), .D(n_899), .Y(n_883) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B(n_890), .Y(n_887) );
AND2x2_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
AND2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
AND2x2_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
HB1xp67_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
HB1xp67_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
HB1xp67_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
NOR2x1_ASAP7_75t_L g915 ( .A(n_916), .B(n_927), .Y(n_915) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_917), .B(n_920), .C(n_922), .Y(n_916) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_932), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_934), .B(n_935), .Y(n_933) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
endmodule