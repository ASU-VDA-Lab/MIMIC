module fake_jpeg_19021_n_101 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_24),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_0),
.C(n_3),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_20),
.B(n_10),
.Y(n_33)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_27),
.B1(n_12),
.B2(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_18),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_23),
.B1(n_27),
.B2(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_39),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_27),
.B1(n_15),
.B2(n_12),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_10),
.B1(n_20),
.B2(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_52),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_67),
.B(n_71),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_69),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_45),
.B1(n_43),
.B2(n_37),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_56),
.B(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_64),
.B(n_68),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.C(n_74),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_57),
.C(n_51),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_51),
.C(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_70),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_56),
.C(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_67),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_66),
.B(n_62),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_79),
.A2(n_75),
.B(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_61),
.B(n_63),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_32),
.B1(n_17),
.B2(n_6),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_4),
.Y(n_93)
);

OAI21x1_ASAP7_75t_SL g92 ( 
.A1(n_90),
.A2(n_81),
.B(n_16),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_94),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_7),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_8),
.C(n_9),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_97),
.B(n_16),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_96),
.A2(n_5),
.A3(n_6),
.B1(n_16),
.B2(n_25),
.C1(n_88),
.C2(n_90),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_25),
.C(n_5),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);


endmodule