module fake_jpeg_18694_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_52),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_58),
.B1(n_21),
.B2(n_34),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_16),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_24),
.B1(n_27),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_22),
.B1(n_30),
.B2(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_16),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_77),
.B1(n_102),
.B2(n_1),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_33),
.B1(n_30),
.B2(n_18),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_16),
.B(n_35),
.C(n_13),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_1),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_72),
.B(n_83),
.Y(n_124)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_84),
.Y(n_111)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_35),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_94),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_21),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_105),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_63),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_61),
.A2(n_34),
.B1(n_32),
.B2(n_26),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_32),
.B1(n_26),
.B2(n_19),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_108),
.B1(n_2),
.B2(n_3),
.Y(n_140)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_1),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_32),
.C(n_26),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_61),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_10),
.B(n_11),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_12),
.B(n_15),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_115),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_19),
.B1(n_29),
.B2(n_23),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_114),
.A2(n_122),
.B1(n_2),
.B2(n_4),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_29),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_102),
.B1(n_76),
.B2(n_105),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_15),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_70),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_14),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_81),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_152),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_97),
.B(n_103),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_170),
.B(n_138),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_90),
.B1(n_105),
.B2(n_97),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_151),
.B1(n_154),
.B2(n_172),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_120),
.B1(n_118),
.B2(n_117),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_150),
.B(n_159),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_110),
.B1(n_87),
.B2(n_82),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_143),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_87),
.B1(n_82),
.B2(n_80),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_89),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_156),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_139),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_126),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_75),
.B(n_85),
.C(n_9),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_164),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_80),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_130),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_4),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_73),
.B1(n_8),
.B2(n_9),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_171),
.B1(n_134),
.B2(n_119),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_2),
.B(n_4),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_11),
.B1(n_12),
.B2(n_5),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_174),
.B(n_190),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_115),
.C(n_125),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_169),
.C(n_154),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_182),
.B1(n_192),
.B2(n_162),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_138),
.B(n_139),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_208)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_167),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_170),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_145),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_118),
.B1(n_117),
.B2(n_121),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_201),
.B1(n_150),
.B2(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_147),
.A2(n_137),
.B1(n_119),
.B2(n_111),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_149),
.A2(n_128),
.B1(n_137),
.B2(n_131),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_155),
.A2(n_134),
.B1(n_5),
.B2(n_6),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_206),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_144),
.A2(n_5),
.B1(n_7),
.B2(n_12),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_171),
.B1(n_159),
.B2(n_168),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_7),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_223),
.B1(n_202),
.B2(n_216),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_160),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_210),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_217),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_215),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_220),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_152),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_231),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_197),
.C(n_196),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_165),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_153),
.B1(n_158),
.B2(n_148),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_222),
.A2(n_188),
.B(n_194),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_177),
.A2(n_7),
.B1(n_198),
.B2(n_176),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_7),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_225),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_175),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_226),
.B(n_194),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_232),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_179),
.B(n_206),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_189),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_199),
.B1(n_177),
.B2(n_198),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_183),
.B1(n_182),
.B2(n_178),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_242),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_237),
.A2(n_252),
.B1(n_224),
.B2(n_214),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_243),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_187),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_210),
.B(n_222),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_205),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_253),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_208),
.B1(n_220),
.B2(n_219),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_226),
.C(n_231),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_218),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_247),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_268),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_235),
.B(n_251),
.Y(n_286)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_246),
.B(n_212),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_262),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_274),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_208),
.B1(n_229),
.B2(n_230),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_272),
.B1(n_243),
.B2(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_270),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_275),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_224),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_250),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_253),
.C(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_288),
.C(n_289),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_255),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_245),
.B1(n_249),
.B2(n_237),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_286),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_239),
.C(n_251),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_239),
.C(n_254),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_262),
.C(n_267),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_288),
.C(n_280),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_263),
.B1(n_265),
.B2(n_264),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_296),
.A2(n_299),
.B1(n_301),
.B2(n_285),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_238),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_235),
.Y(n_298)
);

NOR2x1_ASAP7_75t_R g306 ( 
.A(n_298),
.B(n_273),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_265),
.B1(n_264),
.B2(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_284),
.B(n_258),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_286),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_310),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_287),
.B(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_306),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_309),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_279),
.C(n_280),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_276),
.B1(n_268),
.B2(n_254),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_296),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_293),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_314),
.B(n_315),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_295),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_310),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_319),
.B(n_320),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_305),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_308),
.Y(n_320)
);

OAI21x1_ASAP7_75t_SL g323 ( 
.A1(n_321),
.A2(n_306),
.B(n_304),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_303),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_322),
.C(n_313),
.Y(n_325)
);

OAI321xp33_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_313),
.A3(n_317),
.B1(n_311),
.B2(n_300),
.C(n_302),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_300),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_234),
.C(n_181),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_181),
.Y(n_329)
);


endmodule