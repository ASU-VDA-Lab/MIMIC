module fake_jpeg_23797_n_64 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_64);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_64;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_56;
wire n_31;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_9),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_26),
.B1(n_42),
.B2(n_50),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_49),
.B1(n_41),
.B2(n_53),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_43),
.B(n_31),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_20),
.C(n_23),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_44),
.B2(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_35),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_45),
.B1(n_47),
.B2(n_46),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_48),
.Y(n_64)
);


endmodule