module real_jpeg_33587_n_25 (n_17, n_8, n_0, n_21, n_2, n_188, n_185, n_180, n_10, n_186, n_9, n_12, n_24, n_189, n_187, n_6, n_190, n_183, n_179, n_23, n_11, n_14, n_7, n_22, n_18, n_3, n_5, n_4, n_181, n_1, n_182, n_20, n_19, n_184, n_16, n_15, n_13, n_25);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_188;
input n_185;
input n_180;
input n_10;
input n_186;
input n_9;
input n_12;
input n_24;
input n_189;
input n_187;
input n_6;
input n_190;
input n_183;
input n_179;
input n_23;
input n_11;
input n_14;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_181;
input n_1;
input n_182;
input n_20;
input n_19;
input n_184;
input n_16;
input n_15;
input n_13;

output n_25;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_174;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_0),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_1),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_2),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_2),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_3),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_4),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_5),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_79),
.Y(n_139)
);

AOI221xp5_ASAP7_75t_L g95 ( 
.A1(n_6),
.A2(n_23),
.B1(n_96),
.B2(n_101),
.C(n_105),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_6),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g140 ( 
.A1(n_8),
.A2(n_69),
.A3(n_71),
.B1(n_77),
.B2(n_141),
.C1(n_143),
.C2(n_189),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_9),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_11),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_11),
.B(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_12),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_13),
.B(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_14),
.B(n_52),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_15),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_16),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_16),
.B(n_130),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_17),
.B(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_18),
.Y(n_153)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_21),
.B(n_41),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_22),
.B(n_92),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_23),
.B(n_96),
.C(n_101),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_36),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_47),
.B(n_177),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_80),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_146),
.B(n_162),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_56),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI31xp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_85),
.A3(n_128),
.B(n_136),
.Y(n_58)
);

NOR3xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_76),
.C(n_82),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_60),
.A2(n_137),
.B(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_69),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_62),
.B(n_82),
.C(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_180),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OA21x2_ASAP7_75t_SL g137 ( 
.A1(n_76),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_120),
.C(n_121),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_109),
.B(n_119),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_95),
.B1(n_107),
.B2(n_108),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_185),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_154),
.C(n_157),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_172),
.C(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

OAI322xp33_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_158),
.A3(n_171),
.B1(n_174),
.B2(n_175),
.C1(n_176),
.C2(n_190),
.Y(n_170)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_163),
.B(n_169),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_179),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_181),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_182),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_183),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_184),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_186),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_187),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_188),
.Y(n_131)
);


endmodule