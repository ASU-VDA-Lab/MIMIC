module fake_netlist_5_768_n_1895 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1895);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1895;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_33),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_114),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_90),
.Y(n_198)
);

BUFx8_ASAP7_75t_SL g199 ( 
.A(n_115),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_106),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_181),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_57),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_64),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_77),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_54),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_50),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_96),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_160),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_57),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_18),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_8),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_60),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_76),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_130),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_66),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_176),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_128),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_101),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_42),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_97),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_59),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_119),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_146),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_149),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_110),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_103),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_151),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_112),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_63),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_50),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_182),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_22),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_7),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_129),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_24),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_82),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_183),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_131),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_161),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_166),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_107),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_165),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_134),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_51),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_118),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_55),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_102),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_139),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_167),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_172),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_95),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_180),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_87),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_144),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_111),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_62),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_170),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_138),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_93),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_173),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_7),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_63),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_157),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_147),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_116),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_40),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_58),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_44),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_155),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_22),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_14),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_123),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_88),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_41),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_45),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_125),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_4),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_16),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_41),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_46),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_71),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_25),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_13),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_137),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_156),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_113),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_40),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_175),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_25),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_53),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_190),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_35),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_45),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_158),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_67),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_43),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_98),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_86),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_135),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_28),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_143),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_89),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_30),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_68),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_14),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_47),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_186),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_124),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_174),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_104),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_48),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_99),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_2),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_163),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_8),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_21),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_185),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_44),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_70),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_35),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_75),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_27),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_1),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_132),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_80),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_78),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_184),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_164),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_5),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_79),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_24),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_117),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_56),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_187),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_189),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_11),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_122),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_54),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_121),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_12),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_141),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_56),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_177),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_28),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_9),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_67),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_12),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_37),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_34),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_9),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_4),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_32),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_0),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_53),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_3),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_74),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_49),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_68),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_148),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_29),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_27),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_19),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_65),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_52),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_6),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_60),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_5),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_48),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_178),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_73),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_168),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_72),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_284),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_284),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_203),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_203),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_199),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_284),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_315),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_284),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_193),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_284),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_209),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_217),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_217),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_196),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_198),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_224),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_219),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_232),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_201),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_224),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_297),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_297),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

INVxp33_ASAP7_75t_SL g412 ( 
.A(n_195),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_345),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_342),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_368),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_369),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_215),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_233),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_207),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_215),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_197),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_197),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_213),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_353),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_228),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_228),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_222),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_206),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_223),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_200),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_242),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_225),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_242),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_226),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_231),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_234),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_236),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_257),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_240),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_243),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_244),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_257),
.Y(n_445)
);

INVxp33_ASAP7_75t_SL g446 ( 
.A(n_212),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_274),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_247),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_274),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_287),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_216),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_287),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_292),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_292),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_249),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_294),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_304),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_250),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_200),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_252),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_255),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_304),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_253),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_256),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_306),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_306),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_258),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_317),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_202),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_263),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_194),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_317),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_265),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_266),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_337),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_218),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_267),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_337),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_354),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_354),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_268),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_397),
.B(n_194),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_399),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_420),
.B(n_315),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_396),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_433),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_402),
.B(n_227),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_433),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_405),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_463),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_459),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_451),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_459),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_R g501 ( 
.A(n_412),
.B(n_323),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_403),
.B(n_227),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_463),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_398),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_407),
.B(n_237),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_471),
.B(n_323),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_471),
.B(n_237),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_431),
.B(n_204),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_471),
.B(n_204),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_401),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_463),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_430),
.Y(n_514)
);

AND2x2_ASAP7_75t_SL g515 ( 
.A(n_476),
.B(n_260),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_463),
.B(n_253),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_469),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_390),
.B(n_307),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_469),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_401),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_421),
.B(n_261),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_446),
.B(n_261),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_391),
.B(n_307),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_427),
.A2(n_336),
.B1(n_230),
.B2(n_303),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_395),
.A2(n_296),
.B1(n_246),
.B2(n_382),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_423),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_392),
.B(n_221),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_409),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_432),
.B(n_272),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_424),
.Y(n_531)
);

CKINVDCx6p67_ASAP7_75t_R g532 ( 
.A(n_437),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_388),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_416),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_425),
.B(n_322),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_440),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_419),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_419),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_400),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_428),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_443),
.A2(n_291),
.B1(n_289),
.B2(n_288),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_429),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_429),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_400),
.Y(n_546)
);

AOI22x1_ASAP7_75t_SL g547 ( 
.A1(n_406),
.A2(n_205),
.B1(n_327),
.B2(n_245),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_435),
.B(n_322),
.Y(n_548)
);

OA22x2_ASAP7_75t_L g549 ( 
.A1(n_434),
.A2(n_361),
.B1(n_359),
.B2(n_381),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_434),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_438),
.B(n_221),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_393),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_439),
.B(n_214),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_436),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_404),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

AND2x2_ASAP7_75t_SL g558 ( 
.A(n_441),
.B(n_260),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_408),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_415),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_426),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_554),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_497),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_510),
.B(n_442),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_558),
.A2(n_309),
.B1(n_283),
.B2(n_356),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_515),
.B(n_444),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_486),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_527),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_522),
.B(n_455),
.C(n_448),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_508),
.B(n_283),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_521),
.B(n_458),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_497),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_515),
.B(n_460),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_535),
.B(n_464),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_482),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_484),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_509),
.B(n_202),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_508),
.B(n_473),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_508),
.B(n_408),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_543),
.B(n_474),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_490),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_530),
.B(n_477),
.Y(n_582)
);

NOR2x1p5_ASAP7_75t_L g583 ( 
.A(n_533),
.B(n_356),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_L g584 ( 
.A(n_501),
.B(n_454),
.C(n_239),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_503),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_486),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_503),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_511),
.B(n_410),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_483),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_506),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_558),
.B(n_276),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_520),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_552),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_514),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_548),
.B(n_481),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_526),
.B(n_461),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_486),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_506),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_518),
.A2(n_309),
.B1(n_366),
.B2(n_381),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_483),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_520),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_509),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_487),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_520),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_509),
.Y(n_605)
);

AND3x2_ASAP7_75t_L g606 ( 
.A(n_489),
.B(n_208),
.C(n_210),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_520),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_514),
.Y(n_608)
);

INVx8_ASAP7_75t_L g609 ( 
.A(n_511),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_520),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_524),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_531),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_486),
.Y(n_613)
);

CKINVDCx6p67_ASAP7_75t_R g614 ( 
.A(n_532),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_485),
.B(n_493),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_518),
.A2(n_366),
.B1(n_378),
.B2(n_376),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_524),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_504),
.B(n_467),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_545),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_523),
.B(n_359),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_550),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_499),
.B(n_470),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_524),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_524),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_487),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g627 ( 
.A1(n_491),
.A2(n_502),
.B(n_494),
.Y(n_627)
);

OAI22x1_ASAP7_75t_L g628 ( 
.A1(n_561),
.A2(n_211),
.B1(n_367),
.B2(n_301),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_507),
.A2(n_220),
.B(n_210),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_511),
.B(n_273),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_523),
.B(n_491),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_561),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_551),
.B(n_422),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_529),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g636 ( 
.A(n_528),
.B(n_332),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_536),
.B(n_221),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_538),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_486),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_538),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_529),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_549),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_539),
.B(n_441),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_549),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_536),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_539),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_532),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_529),
.B(n_277),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_541),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_529),
.B(n_286),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_549),
.A2(n_319),
.B1(n_318),
.B2(n_241),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_560),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_542),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_544),
.A2(n_361),
.B1(n_372),
.B2(n_380),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_544),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_557),
.B(n_238),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

BUFx8_ASAP7_75t_SL g660 ( 
.A(n_488),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_496),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_557),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_529),
.B(n_290),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_537),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_560),
.Y(n_665)
);

BUFx6f_ASAP7_75t_SL g666 ( 
.A(n_492),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_537),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_537),
.B(n_295),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_537),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_537),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_502),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_488),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_517),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_516),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_525),
.B(n_272),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_517),
.Y(n_676)
);

BUFx6f_ASAP7_75t_SL g677 ( 
.A(n_498),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_496),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_534),
.B(n_299),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_500),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_496),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_519),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_496),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_556),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_556),
.B(n_272),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_534),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_556),
.B(n_300),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_556),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_556),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_505),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_540),
.B(n_220),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_540),
.A2(n_344),
.B1(n_324),
.B2(n_321),
.Y(n_692)
);

OR2x6_ASAP7_75t_L g693 ( 
.A(n_546),
.B(n_372),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_546),
.A2(n_259),
.B1(n_269),
.B2(n_275),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_505),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_540),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_505),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_553),
.B(n_272),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_512),
.B(n_302),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_553),
.B(n_279),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_505),
.B(n_308),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_505),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_513),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_513),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_516),
.B(n_253),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_513),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_559),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_559),
.Y(n_708)
);

NOR2x1p5_ASAP7_75t_L g709 ( 
.A(n_547),
.B(n_280),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_513),
.B(n_281),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_513),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_516),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_516),
.Y(n_713)
);

INVx8_ASAP7_75t_L g714 ( 
.A(n_609),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_569),
.B(n_312),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_615),
.B(n_253),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_629),
.B(n_253),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_566),
.A2(n_335),
.B1(n_373),
.B2(n_355),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_584),
.B(n_313),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_642),
.A2(n_380),
.B1(n_378),
.B2(n_376),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_605),
.B(n_445),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_632),
.B(n_445),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_571),
.B(n_229),
.Y(n_723)
);

BUFx8_ASAP7_75t_L g724 ( 
.A(n_632),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_638),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_574),
.B(n_229),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_631),
.A2(n_248),
.B(n_235),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_602),
.B(n_235),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_620),
.B(n_447),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_633),
.B(n_564),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_602),
.B(n_248),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_696),
.B(n_251),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_609),
.B(n_591),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_643),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_640),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_696),
.B(n_251),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_583),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_620),
.Y(n_739)
);

AO221x1_ASAP7_75t_L g740 ( 
.A1(n_628),
.A2(n_298),
.B1(n_375),
.B2(n_254),
.C(n_264),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_605),
.B(n_254),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_572),
.Y(n_742)
);

AOI22x1_ASAP7_75t_L g743 ( 
.A1(n_642),
.A2(n_305),
.B1(n_383),
.B2(n_357),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_643),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_644),
.B(n_447),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_572),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_573),
.B(n_293),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_562),
.B(n_449),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_646),
.B(n_262),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_618),
.A2(n_339),
.B1(n_316),
.B2(n_326),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_649),
.B(n_652),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_609),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_644),
.B(n_298),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_578),
.B(n_298),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_L g755 ( 
.A1(n_620),
.A2(n_375),
.B1(n_371),
.B2(n_362),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_645),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_585),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_585),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_568),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_612),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_587),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_620),
.A2(n_282),
.B1(n_285),
.B2(n_305),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_654),
.Y(n_763)
);

BUFx5_ASAP7_75t_L g764 ( 
.A(n_712),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_593),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_562),
.B(n_298),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_672),
.B(n_449),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_570),
.B(n_450),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_655),
.B(n_262),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_691),
.A2(n_285),
.B1(n_282),
.B2(n_370),
.Y(n_770)
);

AND2x4_ASAP7_75t_SL g771 ( 
.A(n_645),
.B(n_495),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_562),
.B(n_298),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_657),
.B(n_264),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_662),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_579),
.B(n_270),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_577),
.B(n_328),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_580),
.B(n_310),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_609),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_579),
.B(n_270),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_587),
.Y(n_780)
);

AND2x4_ASAP7_75t_SL g781 ( 
.A(n_645),
.B(n_495),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_577),
.B(n_331),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_577),
.B(n_674),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_SL g784 ( 
.A1(n_653),
.A2(n_374),
.B1(n_314),
.B2(n_320),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_SL g785 ( 
.A(n_666),
.B(n_325),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_575),
.B(n_271),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_648),
.A2(n_357),
.B(n_271),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_588),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_588),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_SL g790 ( 
.A1(n_594),
.A2(n_350),
.B1(n_329),
.B2(n_330),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_680),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_680),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_674),
.B(n_338),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_595),
.B(n_334),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_674),
.B(n_346),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_712),
.B(n_516),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_575),
.B(n_340),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_576),
.B(n_340),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_619),
.B(n_343),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_576),
.B(n_341),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_622),
.B(n_347),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_682),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_636),
.A2(n_630),
.B1(n_596),
.B2(n_582),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_674),
.B(n_348),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_570),
.B(n_450),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_570),
.A2(n_370),
.B1(n_341),
.B2(n_383),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_713),
.B(n_516),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_682),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_636),
.A2(n_570),
.B1(n_635),
.B2(n_710),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_581),
.B(n_349),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_606),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_658),
.B(n_599),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_589),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_565),
.B(n_379),
.C(n_352),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_600),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_660),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_581),
.B(n_351),
.Y(n_817)
);

NOR3xp33_ASAP7_75t_SL g818 ( 
.A(n_675),
.B(n_364),
.C(n_365),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_623),
.B(n_452),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_653),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_616),
.A2(n_384),
.B1(n_386),
.B2(n_360),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_651),
.A2(n_453),
.B(n_480),
.C(n_479),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_600),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_SL g824 ( 
.A1(n_665),
.A2(n_358),
.B1(n_377),
.B2(n_547),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_660),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_603),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_603),
.B(n_626),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_699),
.B(n_278),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_626),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_674),
.B(n_278),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_709),
.B(n_452),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_590),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_691),
.A2(n_480),
.B1(n_479),
.B2(n_478),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_684),
.B(n_691),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_628),
.B(n_453),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_692),
.A2(n_700),
.B1(n_679),
.B2(n_685),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_598),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_693),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_656),
.A2(n_478),
.B1(n_475),
.B2(n_472),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_687),
.B(n_456),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_707),
.A2(n_465),
.B(n_472),
.C(n_468),
.Y(n_841)
);

OR2x2_ASAP7_75t_SL g842 ( 
.A(n_637),
.B(n_456),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_598),
.Y(n_843)
);

AND2x6_ASAP7_75t_L g844 ( 
.A(n_713),
.B(n_457),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_707),
.B(n_708),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_594),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_693),
.A2(n_694),
.B(n_705),
.C(n_698),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_693),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_671),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_708),
.B(n_457),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_693),
.A2(n_475),
.B1(n_468),
.B2(n_466),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_686),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_684),
.B(n_278),
.Y(n_853)
);

AND2x4_ASAP7_75t_SL g854 ( 
.A(n_614),
.B(n_278),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_665),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_671),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_695),
.A2(n_466),
.B(n_465),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_650),
.B(n_462),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_666),
.B(n_311),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_673),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_663),
.B(n_462),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_676),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_627),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_604),
.B(n_311),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_668),
.B(n_410),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_627),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_688),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_701),
.A2(n_418),
.B1(n_417),
.B2(n_414),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_688),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_689),
.B(n_411),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_604),
.B(n_311),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_666),
.B(n_311),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_607),
.B(n_333),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_607),
.B(n_333),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_705),
.A2(n_418),
.B(n_417),
.C(n_414),
.Y(n_875)
);

INVxp33_ASAP7_75t_L g876 ( 
.A(n_608),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_610),
.B(n_385),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_689),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_734),
.B(n_670),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_721),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_849),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_824),
.A2(n_608),
.B1(n_647),
.B2(n_614),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_SL g883 ( 
.A1(n_846),
.A2(n_647),
.B1(n_411),
.B2(n_413),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_734),
.B(n_723),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_726),
.B(n_670),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_856),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_721),
.Y(n_887)
);

BUFx12f_ASAP7_75t_L g888 ( 
.A(n_724),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_737),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_730),
.B(n_677),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_812),
.B(n_610),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_724),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_748),
.B(n_677),
.Y(n_893)
);

AO22x1_ASAP7_75t_L g894 ( 
.A1(n_777),
.A2(n_413),
.B1(n_677),
.B2(n_711),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_722),
.B(n_333),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_725),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_767),
.B(n_611),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_803),
.B(n_611),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_768),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_765),
.B(n_664),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_744),
.B(n_819),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_788),
.B(n_333),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_789),
.B(n_667),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_735),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_828),
.A2(n_669),
.B1(n_621),
.B2(n_634),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_840),
.B(n_617),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_813),
.B(n_617),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_778),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_815),
.B(n_621),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_823),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_778),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_778),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_745),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_826),
.B(n_624),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_778),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_829),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_805),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_858),
.B(n_624),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_861),
.B(n_634),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_852),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_794),
.B(n_729),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_771),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_844),
.Y(n_923)
);

BUFx2_ASAP7_75t_SL g924 ( 
.A(n_756),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_739),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_781),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_742),
.Y(n_927)
);

NOR2xp67_ASAP7_75t_L g928 ( 
.A(n_738),
.B(n_641),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_SL g929 ( 
.A1(n_717),
.A2(n_669),
.B(n_641),
.C(n_706),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_827),
.B(n_597),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_791),
.B(n_597),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_739),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_746),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_792),
.B(n_597),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_855),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_755),
.B(n_385),
.C(n_2),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_SL g937 ( 
.A(n_818),
.B(n_756),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_836),
.A2(n_809),
.B1(n_770),
.B2(n_747),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_714),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_757),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_820),
.B(n_697),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_764),
.B(n_697),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_764),
.B(n_702),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_845),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_802),
.B(n_639),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_835),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_844),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_808),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_763),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_717),
.A2(n_385),
.B1(n_704),
.B2(n_706),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_838),
.Y(n_951)
);

INVx5_ASAP7_75t_L g952 ( 
.A(n_844),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_816),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_794),
.B(n_592),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_811),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_828),
.A2(n_592),
.B1(n_601),
.B2(n_625),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_774),
.B(n_751),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_863),
.A2(n_703),
.B(n_690),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_747),
.B(n_592),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_L g960 ( 
.A(n_714),
.B(n_844),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_755),
.B(n_601),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_764),
.B(n_601),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_857),
.B(n_639),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_754),
.A2(n_625),
.B1(n_678),
.B2(n_681),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_714),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_752),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_865),
.B(n_639),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_SL g968 ( 
.A1(n_859),
.A2(n_872),
.B1(n_854),
.B2(n_790),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_775),
.B(n_703),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_779),
.B(n_759),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_876),
.B(n_625),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_764),
.B(n_567),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_760),
.B(n_683),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_799),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_867),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_869),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_878),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_764),
.B(n_567),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_862),
.B(n_659),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_859),
.B(n_678),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_716),
.B(n_703),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_799),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_716),
.A2(n_690),
.B1(n_659),
.B2(n_681),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_758),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_761),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_780),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_SL g987 ( 
.A(n_825),
.B(n_683),
.Y(n_987)
);

NAND2x1p5_ASAP7_75t_L g988 ( 
.A(n_752),
.B(n_683),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_844),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_870),
.Y(n_990)
);

AND2x4_ASAP7_75t_SL g991 ( 
.A(n_831),
.B(n_567),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_784),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_832),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_860),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_728),
.B(n_659),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_837),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_731),
.B(n_690),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_770),
.B(n_661),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_843),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_818),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_SL g1001 ( 
.A(n_831),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_764),
.B(n_661),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_741),
.B(n_661),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_842),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_831),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_866),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_720),
.A2(n_661),
.B1(n_613),
.B2(n_586),
.Y(n_1007)
);

NAND2x1p5_ASAP7_75t_L g1008 ( 
.A(n_783),
.B(n_834),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_850),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_732),
.B(n_661),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_866),
.Y(n_1011)
);

OR2x6_ASAP7_75t_L g1012 ( 
.A(n_848),
.B(n_613),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_766),
.B(n_613),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_736),
.B(n_613),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_SL g1015 ( 
.A1(n_787),
.A2(n_613),
.B(n_586),
.C(n_567),
.Y(n_1015)
);

BUFx4f_ASAP7_75t_SL g1016 ( 
.A(n_766),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_834),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_SL g1018 ( 
.A1(n_872),
.A2(n_586),
.B1(n_567),
.B2(n_6),
.Y(n_1018)
);

NOR2x2_ASAP7_75t_L g1019 ( 
.A(n_762),
.B(n_0),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_801),
.B(n_586),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_783),
.Y(n_1021)
);

NAND3xp33_ASAP7_75t_SL g1022 ( 
.A(n_750),
.B(n_3),
.C(n_10),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_749),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_SL g1024 ( 
.A1(n_814),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_1024)
);

BUFx8_ASAP7_75t_L g1025 ( 
.A(n_740),
.Y(n_1025)
);

NOR2x2_ASAP7_75t_L g1026 ( 
.A(n_762),
.B(n_15),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_786),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_801),
.B(n_15),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_753),
.B(n_16),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_769),
.Y(n_1030)
);

NAND2x1p5_ASAP7_75t_L g1031 ( 
.A(n_753),
.B(n_162),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_719),
.B(n_120),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_772),
.B(n_17),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_772),
.B(n_17),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_773),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_797),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_798),
.B(n_18),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_800),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_810),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_SL g1040 ( 
.A1(n_720),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_743),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_1041)
);

AND2x4_ASAP7_75t_SL g1042 ( 
.A(n_833),
.B(n_159),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_715),
.B(n_154),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_847),
.B(n_145),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_727),
.B(n_23),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_833),
.A2(n_142),
.B1(n_136),
.B2(n_133),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_822),
.A2(n_26),
.B(n_29),
.C(n_30),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_793),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_851),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_868),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_841),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_776),
.B(n_31),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_817),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_864),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_718),
.B(n_127),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_776),
.B(n_31),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_782),
.B(n_32),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_782),
.B(n_126),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_795),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_853),
.B(n_877),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_974),
.B(n_785),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_938),
.A2(n_795),
.B(n_804),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_R g1063 ( 
.A(n_1000),
.B(n_733),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_SL g1064 ( 
.A1(n_890),
.A2(n_796),
.B(n_807),
.C(n_875),
.Y(n_1064)
);

BUFx12f_ASAP7_75t_L g1065 ( 
.A(n_888),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_1057),
.A2(n_853),
.B(n_874),
.C(n_873),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_SL g1067 ( 
.A(n_953),
.B(n_806),
.Y(n_1067)
);

AOI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_974),
.A2(n_821),
.B(n_806),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_962),
.A2(n_804),
.B(n_830),
.Y(n_1069)
);

OR2x6_ASAP7_75t_L g1070 ( 
.A(n_924),
.B(n_830),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_884),
.B(n_877),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_1028),
.A2(n_874),
.B(n_873),
.C(n_871),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_897),
.B(n_871),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_942),
.A2(n_864),
.B(n_839),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_1044),
.A2(n_33),
.B(n_34),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_962),
.A2(n_839),
.B(n_108),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_1057),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_901),
.B(n_899),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1058),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_925),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_913),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_939),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_925),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_892),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_982),
.B(n_42),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1020),
.A2(n_978),
.B(n_972),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_895),
.A2(n_43),
.B(n_46),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_982),
.B(n_47),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_896),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1058),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_921),
.B(n_55),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_880),
.B(n_92),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1053),
.A2(n_100),
.B1(n_85),
.B2(n_84),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_SL g1094 ( 
.A1(n_1042),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1040),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_1095)
);

CKINVDCx6p67_ASAP7_75t_R g1096 ( 
.A(n_892),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_972),
.A2(n_69),
.B(n_81),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_944),
.B(n_65),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_882),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_1005),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_978),
.A2(n_66),
.B(n_1002),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_904),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_922),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1047),
.A2(n_891),
.B(n_1037),
.C(n_970),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1002),
.A2(n_954),
.B(n_959),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_893),
.B(n_957),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_939),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1009),
.B(n_1038),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_898),
.A2(n_1044),
.B(n_963),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1039),
.B(n_1027),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_939),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_908),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_968),
.B(n_1030),
.Y(n_1113)
);

OAI21xp33_ASAP7_75t_L g1114 ( 
.A1(n_902),
.A2(n_936),
.B(n_949),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1036),
.B(n_990),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1056),
.A2(n_1033),
.B1(n_1022),
.B2(n_1055),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_915),
.A2(n_1003),
.B(n_1007),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_922),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_961),
.A2(n_887),
.B1(n_1060),
.B2(n_980),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1036),
.B(n_1023),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_917),
.B(n_1004),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1047),
.A2(n_1050),
.B(n_1033),
.C(n_1055),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_889),
.Y(n_1123)
);

OR2x2_ASAP7_75t_L g1124 ( 
.A(n_941),
.B(n_946),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_915),
.A2(n_1007),
.B(n_958),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_955),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1023),
.B(n_910),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_916),
.B(n_948),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_932),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_879),
.B(n_920),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_971),
.B(n_987),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1035),
.B(n_1016),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1054),
.A2(n_961),
.B(n_1017),
.C(n_1052),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_926),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_992),
.B(n_1016),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_915),
.A2(n_969),
.B(n_1011),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1050),
.A2(n_1049),
.B(n_1034),
.C(n_1045),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_975),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_935),
.B(n_883),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_928),
.B(n_1005),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_926),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_976),
.B(n_977),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_900),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_915),
.A2(n_1006),
.B(n_1011),
.Y(n_1144)
);

NAND2xp33_ASAP7_75t_SL g1145 ( 
.A(n_939),
.B(n_965),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1006),
.A2(n_930),
.B(n_898),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_900),
.B(n_951),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_903),
.B(n_1049),
.Y(n_1148)
);

BUFx8_ASAP7_75t_L g1149 ( 
.A(n_1001),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_965),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_998),
.A2(n_1017),
.B(n_885),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1008),
.A2(n_1021),
.B1(n_973),
.B2(n_956),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1008),
.A2(n_1021),
.B1(n_973),
.B2(n_952),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_952),
.A2(n_1042),
.B1(n_1013),
.B2(n_1035),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_951),
.B(n_994),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_908),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_903),
.B(n_1035),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1018),
.A2(n_1025),
.B1(n_1059),
.B2(n_1048),
.Y(n_1158)
);

CKINVDCx16_ASAP7_75t_R g1159 ( 
.A(n_1001),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1025),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_SL g1161 ( 
.A(n_1024),
.B(n_936),
.C(n_1041),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_906),
.B(n_918),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_919),
.B(n_881),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_988),
.A2(n_942),
.B(n_943),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_988),
.A2(n_943),
.B(n_967),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1010),
.A2(n_1014),
.B(n_960),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_991),
.Y(n_1167)
);

NOR2x1_ASAP7_75t_L g1168 ( 
.A(n_966),
.B(n_965),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1029),
.A2(n_1051),
.B(n_909),
.C(n_914),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_995),
.A2(n_997),
.B(n_952),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_952),
.A2(n_1013),
.B(n_1015),
.Y(n_1171)
);

AOI33xp33_ASAP7_75t_L g1172 ( 
.A1(n_1041),
.A2(n_950),
.A3(n_991),
.B1(n_999),
.B2(n_996),
.B3(n_1032),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_886),
.A2(n_947),
.B(n_923),
.C(n_1043),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_907),
.A2(n_981),
.B(n_931),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_934),
.A2(n_945),
.B(n_979),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_923),
.A2(n_947),
.B1(n_983),
.B2(n_966),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1048),
.B(n_1059),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1015),
.A2(n_929),
.B(n_983),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_937),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_881),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1012),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_929),
.A2(n_964),
.B(n_908),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_933),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1043),
.B(n_1032),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1019),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1046),
.A2(n_984),
.B(n_986),
.C(n_985),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_965),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_908),
.A2(n_912),
.B(n_911),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_927),
.A2(n_940),
.B(n_950),
.C(n_986),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_911),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_993),
.B(n_985),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_905),
.A2(n_911),
.B1(n_912),
.B2(n_989),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_993),
.B(n_984),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_911),
.A2(n_912),
.B(n_1048),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_894),
.B(n_1012),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1012),
.A2(n_989),
.B(n_1031),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_989),
.B(n_1031),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_L g1198 ( 
.A(n_1026),
.B(n_938),
.C(n_623),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_884),
.B(n_615),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_938),
.A2(n_1040),
.B1(n_1057),
.B2(n_1022),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_941),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_938),
.A2(n_1044),
.B(n_891),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_974),
.B(n_982),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_938),
.A2(n_884),
.B(n_1028),
.C(n_629),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_924),
.B(n_922),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_938),
.A2(n_1057),
.B(n_982),
.C(n_974),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_962),
.A2(n_866),
.B(n_1020),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_896),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_938),
.A2(n_884),
.B(n_1028),
.C(n_629),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1204),
.A2(n_1209),
.B(n_1206),
.Y(n_1210)
);

AOI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1171),
.A2(n_1178),
.B(n_1182),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1089),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1146),
.A2(n_1164),
.B(n_1207),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_SL g1214 ( 
.A(n_1154),
.B(n_1190),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1106),
.B(n_1143),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1190),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1109),
.A2(n_1165),
.B(n_1105),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1166),
.A2(n_1174),
.B(n_1086),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1198),
.B(n_1185),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1202),
.A2(n_1162),
.B(n_1125),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_1062),
.A2(n_1151),
.B(n_1175),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1108),
.B(n_1115),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1152),
.A2(n_1209),
.B(n_1204),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1200),
.B(n_1198),
.C(n_1116),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1147),
.B(n_1201),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1200),
.B(n_1119),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1103),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1136),
.A2(n_1196),
.B(n_1170),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1143),
.B(n_1148),
.Y(n_1229)
);

AO22x1_ASAP7_75t_L g1230 ( 
.A1(n_1135),
.A2(n_1139),
.B1(n_1110),
.B2(n_1091),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1069),
.A2(n_1186),
.B(n_1144),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1078),
.B(n_1184),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1075),
.A2(n_1133),
.A3(n_1066),
.B(n_1189),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1130),
.A2(n_1113),
.B1(n_1120),
.B2(n_1157),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_1129),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_SL g1236 ( 
.A(n_1095),
.B(n_1122),
.C(n_1087),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1169),
.A2(n_1137),
.B(n_1153),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1122),
.A2(n_1161),
.B(n_1068),
.C(n_1085),
.Y(n_1238)
);

BUFx12f_ASAP7_75t_L g1239 ( 
.A(n_1065),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1129),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1186),
.A2(n_1192),
.B(n_1074),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1149),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1169),
.A2(n_1137),
.B(n_1104),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1117),
.A2(n_1194),
.B(n_1101),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1149),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1118),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1197),
.A2(n_1076),
.B(n_1176),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1071),
.B(n_1172),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1134),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1104),
.A2(n_1173),
.B(n_1163),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1127),
.A2(n_1128),
.B1(n_1142),
.B2(n_1073),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1188),
.A2(n_1177),
.B(n_1193),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1099),
.Y(n_1253)
);

NAND2xp33_ASAP7_75t_L g1254 ( 
.A(n_1082),
.B(n_1111),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1191),
.A2(n_1097),
.B(n_1180),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_SL g1256 ( 
.A1(n_1072),
.A2(n_1131),
.B(n_1092),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1203),
.B(n_1098),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1208),
.B(n_1102),
.Y(n_1258)
);

AOI221xp5_ASAP7_75t_L g1259 ( 
.A1(n_1161),
.A2(n_1095),
.B1(n_1088),
.B2(n_1090),
.C(n_1079),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1080),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1094),
.A2(n_1114),
.B1(n_1158),
.B2(n_1061),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1080),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1183),
.A2(n_1072),
.B(n_1168),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1138),
.B(n_1155),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1124),
.B(n_1132),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1126),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1112),
.A2(n_1156),
.B(n_1081),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1077),
.A2(n_1181),
.B(n_1064),
.C(n_1083),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1195),
.B(n_1092),
.Y(n_1269)
);

AOI211x1_ASAP7_75t_L g1270 ( 
.A1(n_1094),
.A2(n_1067),
.B(n_1083),
.C(n_1063),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_1190),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1084),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1190),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1107),
.Y(n_1274)
);

INVx3_ASAP7_75t_SL g1275 ( 
.A(n_1096),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1093),
.A2(n_1145),
.B(n_1121),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1107),
.A2(n_1150),
.B(n_1082),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1082),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1140),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_SL g1280 ( 
.A1(n_1070),
.A2(n_1179),
.B(n_1187),
.Y(n_1280)
);

O2A1O1Ixp33_ASAP7_75t_SL g1281 ( 
.A1(n_1070),
.A2(n_1160),
.B(n_1140),
.C(n_1167),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1111),
.A2(n_1150),
.B(n_1187),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1111),
.A2(n_1150),
.B(n_1187),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1111),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1141),
.B(n_1150),
.Y(n_1285)
);

AOI21x1_ASAP7_75t_SL g1286 ( 
.A1(n_1187),
.A2(n_1205),
.B(n_1100),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1205),
.Y(n_1287)
);

BUFx10_ASAP7_75t_L g1288 ( 
.A(n_1159),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1290)
);

INVx5_ASAP7_75t_L g1291 ( 
.A(n_1190),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1204),
.A2(n_938),
.B(n_1209),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1178),
.A2(n_938),
.A3(n_1075),
.B(n_1171),
.Y(n_1293)
);

CKINVDCx11_ASAP7_75t_R g1294 ( 
.A(n_1065),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1123),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_SL g1296 ( 
.A1(n_1152),
.A2(n_938),
.B(n_752),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1106),
.B(n_748),
.Y(n_1297)
);

AO22x2_ASAP7_75t_L g1298 ( 
.A1(n_1161),
.A2(n_938),
.B1(n_1198),
.B2(n_1113),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1106),
.B(n_748),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1204),
.A2(n_938),
.B(n_1209),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1301)
);

AOI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1171),
.A2(n_1178),
.B(n_1044),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1078),
.B(n_672),
.Y(n_1303)
);

NOR4xp25_ASAP7_75t_L g1304 ( 
.A(n_1095),
.B(n_1200),
.C(n_1161),
.D(n_1206),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1305)
);

AOI31xp67_ASAP7_75t_L g1306 ( 
.A1(n_1113),
.A2(n_1044),
.A3(n_716),
.B(n_898),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1140),
.B(n_1167),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1200),
.A2(n_1161),
.B1(n_1198),
.B2(n_938),
.Y(n_1308)
);

NOR4xp25_ASAP7_75t_L g1309 ( 
.A(n_1095),
.B(n_1200),
.C(n_1161),
.D(n_1206),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1080),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1178),
.A2(n_938),
.A3(n_1075),
.B(n_1171),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1106),
.B(n_748),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1089),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1129),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1089),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1146),
.A2(n_1164),
.B(n_1207),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1204),
.A2(n_938),
.B(n_1209),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1178),
.A2(n_938),
.A3(n_1075),
.B(n_1171),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_SL g1322 ( 
.A1(n_1075),
.A2(n_1196),
.B(n_1125),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1089),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1200),
.A2(n_1161),
.B1(n_1198),
.B2(n_938),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1146),
.A2(n_1164),
.B(n_1207),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1089),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1190),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1190),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1178),
.A2(n_938),
.A3(n_1075),
.B(n_1171),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1204),
.A2(n_1209),
.B(n_938),
.C(n_1122),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1178),
.A2(n_938),
.A3(n_1075),
.B(n_1171),
.Y(n_1333)
);

AO21x1_ASAP7_75t_L g1334 ( 
.A1(n_1204),
.A2(n_938),
.B(n_1209),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1107),
.Y(n_1336)
);

AOI211xp5_ASAP7_75t_L g1337 ( 
.A1(n_1198),
.A2(n_633),
.B(n_794),
.C(n_525),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1089),
.Y(n_1338)
);

INVx5_ASAP7_75t_L g1339 ( 
.A(n_1190),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1089),
.Y(n_1340)
);

AO21x2_ASAP7_75t_L g1341 ( 
.A1(n_1202),
.A2(n_1171),
.B(n_1178),
.Y(n_1341)
);

AO32x2_ASAP7_75t_L g1342 ( 
.A1(n_1152),
.A2(n_938),
.A3(n_1040),
.B1(n_1192),
.B2(n_1153),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1343)
);

AOI221x1_ASAP7_75t_L g1344 ( 
.A1(n_1198),
.A2(n_938),
.B1(n_1161),
.B2(n_1206),
.C(n_1202),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1129),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1146),
.A2(n_1164),
.B(n_1207),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1123),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1105),
.A2(n_1202),
.B(n_1162),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1103),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1089),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1204),
.A2(n_938),
.B(n_1209),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1089),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1204),
.A2(n_938),
.B(n_1209),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1129),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1103),
.Y(n_1356)
);

OA22x2_ASAP7_75t_L g1357 ( 
.A1(n_1185),
.A2(n_1040),
.B1(n_525),
.B2(n_675),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1103),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1204),
.A2(n_1209),
.B(n_938),
.C(n_1122),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1206),
.A2(n_938),
.B(n_1028),
.C(n_1113),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1199),
.B(n_1106),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_SL g1362 ( 
.A(n_1200),
.B(n_1198),
.C(n_726),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1258),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1231),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1295),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1291),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1269),
.B(n_1279),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1243),
.A2(n_1237),
.B(n_1223),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1298),
.B(n_1308),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1224),
.A2(n_1357),
.B1(n_1298),
.B2(n_1315),
.Y(n_1370)
);

NAND2x1p5_ASAP7_75t_L g1371 ( 
.A(n_1291),
.B(n_1339),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1308),
.A2(n_1324),
.B1(n_1328),
.B2(n_1361),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1235),
.B(n_1265),
.Y(n_1373)
);

AOI322xp5_ASAP7_75t_L g1374 ( 
.A1(n_1324),
.A2(n_1259),
.A3(n_1236),
.B1(n_1226),
.B2(n_1362),
.C1(n_1261),
.C2(n_1215),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1218),
.A2(n_1302),
.B(n_1217),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1213),
.A2(n_1325),
.B(n_1319),
.Y(n_1377)
);

INVx4_ASAP7_75t_L g1378 ( 
.A(n_1291),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1301),
.A2(n_1346),
.B1(n_1314),
.B2(n_1335),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1362),
.A2(n_1226),
.B1(n_1236),
.B2(n_1298),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1347),
.A2(n_1228),
.B(n_1244),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1247),
.A2(n_1255),
.B(n_1250),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1304),
.B(n_1309),
.Y(n_1383)
);

AO32x2_ASAP7_75t_L g1384 ( 
.A1(n_1234),
.A2(n_1251),
.A3(n_1334),
.B1(n_1354),
.B2(n_1352),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1295),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1305),
.B(n_1311),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1227),
.Y(n_1387)
);

AOI332xp33_ASAP7_75t_L g1388 ( 
.A1(n_1261),
.A2(n_1219),
.A3(n_1357),
.B1(n_1229),
.B2(n_1318),
.B3(n_1353),
.C1(n_1316),
.C2(n_1212),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1348),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1263),
.A2(n_1252),
.B(n_1220),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1313),
.A2(n_1332),
.B1(n_1343),
.B2(n_1337),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1238),
.B(n_1297),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1349),
.A2(n_1322),
.B(n_1267),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1210),
.A2(n_1320),
.B(n_1300),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1291),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1360),
.A2(n_1238),
.B(n_1344),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1360),
.A2(n_1248),
.B(n_1299),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1331),
.A2(n_1359),
.B(n_1256),
.Y(n_1398)
);

NAND2x1p5_ASAP7_75t_L g1399 ( 
.A(n_1339),
.B(n_1269),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1215),
.B(n_1222),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1331),
.A2(n_1359),
.B(n_1248),
.Y(n_1401)
);

AOI22x1_ASAP7_75t_L g1402 ( 
.A1(n_1280),
.A2(n_1326),
.B1(n_1340),
.B2(n_1338),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1257),
.A2(n_1268),
.B(n_1276),
.C(n_1264),
.Y(n_1403)
);

OAI222xp33_ASAP7_75t_L g1404 ( 
.A1(n_1317),
.A2(n_1355),
.B1(n_1345),
.B2(n_1240),
.C1(n_1262),
.C2(n_1303),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1221),
.A2(n_1286),
.B(n_1283),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1221),
.A2(n_1277),
.B(n_1282),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1341),
.A2(n_1214),
.B(n_1306),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1232),
.A2(n_1225),
.B(n_1281),
.Y(n_1408)
);

AO32x2_ASAP7_75t_L g1409 ( 
.A1(n_1342),
.A2(n_1321),
.A3(n_1293),
.B1(n_1330),
.B2(n_1333),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1230),
.B(n_1270),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1242),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1342),
.B(n_1323),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_SL g1413 ( 
.A1(n_1271),
.A2(n_1273),
.B(n_1284),
.C(n_1351),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1260),
.B(n_1310),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1341),
.A2(n_1254),
.B(n_1271),
.Y(n_1415)
);

OAI21xp33_ASAP7_75t_L g1416 ( 
.A1(n_1310),
.A2(n_1249),
.B(n_1246),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1281),
.A2(n_1266),
.B(n_1287),
.C(n_1285),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1307),
.A2(n_1274),
.B(n_1336),
.Y(n_1418)
);

AO31x2_ASAP7_75t_L g1419 ( 
.A1(n_1233),
.A2(n_1293),
.A3(n_1333),
.B(n_1330),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_SL g1420 ( 
.A1(n_1350),
.A2(n_1358),
.B(n_1356),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1275),
.A2(n_1307),
.B(n_1227),
.C(n_1249),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1312),
.Y(n_1422)
);

AO32x2_ASAP7_75t_L g1423 ( 
.A1(n_1312),
.A2(n_1333),
.A3(n_1330),
.B1(n_1321),
.B2(n_1233),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1233),
.A2(n_1333),
.B(n_1321),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1278),
.A2(n_1336),
.B(n_1274),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1312),
.A2(n_1321),
.B(n_1233),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1246),
.B(n_1216),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1272),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1312),
.A2(n_1339),
.B(n_1278),
.C(n_1216),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1339),
.A2(n_1216),
.B(n_1327),
.C(n_1329),
.Y(n_1430)
);

O2A1O1Ixp5_ASAP7_75t_L g1431 ( 
.A1(n_1288),
.A2(n_1216),
.B(n_1327),
.C(n_1329),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1327),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1329),
.A2(n_1288),
.B(n_1275),
.Y(n_1433)
);

OR2x6_ASAP7_75t_L g1434 ( 
.A(n_1239),
.B(n_1242),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1245),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1245),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1253),
.Y(n_1437)
);

NOR2xp67_ASAP7_75t_L g1438 ( 
.A(n_1239),
.B(n_1294),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1294),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1224),
.B(n_1289),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1231),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1235),
.B(n_1265),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1292),
.A2(n_1320),
.B(n_1300),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1291),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1243),
.A2(n_1237),
.B(n_1223),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1337),
.B(n_1200),
.C(n_1224),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1295),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1360),
.A2(n_938),
.B(n_1238),
.Y(n_1448)
);

OAI22x1_ASAP7_75t_L g1449 ( 
.A1(n_1224),
.A2(n_1226),
.B1(n_1113),
.B2(n_1215),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1231),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1227),
.Y(n_1451)
);

BUFx2_ASAP7_75t_R g1452 ( 
.A(n_1272),
.Y(n_1452)
);

BUFx4f_ASAP7_75t_L g1453 ( 
.A(n_1307),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1235),
.B(n_1265),
.Y(n_1454)
);

O2A1O1Ixp5_ASAP7_75t_L g1455 ( 
.A1(n_1292),
.A2(n_1300),
.B(n_1320),
.C(n_1352),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1258),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1292),
.A2(n_1320),
.B(n_1300),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1337),
.A2(n_636),
.B1(n_1198),
.B2(n_489),
.C(n_1200),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1308),
.A2(n_1200),
.B1(n_1324),
.B2(n_1290),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1231),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1292),
.A2(n_1320),
.B(n_1300),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1231),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1295),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1298),
.B(n_1308),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1224),
.A2(n_1198),
.B1(n_1324),
.B2(n_1308),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1292),
.A2(n_1320),
.B(n_1300),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1235),
.B(n_1265),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1295),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1231),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1295),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1295),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1272),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1296),
.B(n_1256),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1289),
.B(n_1361),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1291),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1289),
.B(n_1361),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1231),
.Y(n_1477)
);

AO21x2_ASAP7_75t_L g1478 ( 
.A1(n_1292),
.A2(n_1320),
.B(n_1300),
.Y(n_1478)
);

NAND2x1p5_ASAP7_75t_L g1479 ( 
.A(n_1291),
.B(n_1339),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1269),
.B(n_1279),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1295),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1224),
.B(n_1289),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1211),
.A2(n_1241),
.B(n_1231),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1227),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1295),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1360),
.A2(n_938),
.B(n_1238),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1243),
.A2(n_1237),
.B(n_1223),
.Y(n_1487)
);

NOR2xp67_ASAP7_75t_L g1488 ( 
.A(n_1266),
.B(n_765),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1258),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1224),
.A2(n_536),
.B1(n_514),
.B2(n_1198),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1291),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1295),
.Y(n_1492)
);

AO31x2_ASAP7_75t_L g1493 ( 
.A1(n_1334),
.A2(n_1331),
.A3(n_1359),
.B(n_1243),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1289),
.B(n_1361),
.Y(n_1494)
);

INVx6_ASAP7_75t_L g1495 ( 
.A(n_1291),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1291),
.Y(n_1496)
);

NAND2x1p5_ASAP7_75t_L g1497 ( 
.A(n_1291),
.B(n_1339),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1295),
.Y(n_1498)
);

AO31x2_ASAP7_75t_L g1499 ( 
.A1(n_1334),
.A2(n_1331),
.A3(n_1359),
.B(n_1243),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1387),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1414),
.B(n_1373),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1472),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1440),
.B(n_1482),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1440),
.B(n_1482),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1400),
.B(n_1392),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1400),
.B(n_1392),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1465),
.A2(n_1446),
.B1(n_1458),
.B2(n_1490),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1380),
.A2(n_1459),
.B1(n_1410),
.B2(n_1370),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1375),
.A2(n_1494),
.B1(n_1476),
.B2(n_1474),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1411),
.A2(n_1434),
.B1(n_1391),
.B2(n_1472),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1379),
.B(n_1386),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1372),
.A2(n_1383),
.B(n_1448),
.C(n_1486),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1383),
.A2(n_1398),
.B1(n_1416),
.B2(n_1396),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1364),
.A2(n_1450),
.B(n_1441),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1364),
.A2(n_1450),
.B(n_1441),
.Y(n_1515)
);

NAND2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1378),
.B(n_1402),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1408),
.A2(n_1453),
.B1(n_1473),
.B2(n_1363),
.Y(n_1517)
);

O2A1O1Ixp5_ASAP7_75t_L g1518 ( 
.A1(n_1455),
.A2(n_1403),
.B(n_1415),
.C(n_1397),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1453),
.A2(n_1473),
.B1(n_1456),
.B2(n_1489),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1442),
.B(n_1454),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1374),
.B(n_1467),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1449),
.B(n_1369),
.Y(n_1522)
);

O2A1O1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1403),
.A2(n_1404),
.B(n_1417),
.C(n_1421),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1395),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1430),
.A2(n_1473),
.B(n_1497),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1367),
.B(n_1480),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1449),
.B(n_1464),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1388),
.A2(n_1453),
.B(n_1431),
.C(n_1430),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1427),
.B(n_1418),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1428),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1443),
.B(n_1457),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1443),
.B(n_1457),
.Y(n_1532)
);

INVx5_ASAP7_75t_L g1533 ( 
.A(n_1395),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1411),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1427),
.B(n_1412),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1461),
.B(n_1478),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1461),
.B(n_1478),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1466),
.A2(n_1394),
.B(n_1445),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1427),
.B(n_1412),
.Y(n_1539)
);

OAI211xp5_ASAP7_75t_L g1540 ( 
.A1(n_1394),
.A2(n_1401),
.B(n_1488),
.C(n_1368),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1466),
.A2(n_1394),
.B(n_1413),
.C(n_1429),
.Y(n_1541)
);

O2A1O1Ixp5_ASAP7_75t_L g1542 ( 
.A1(n_1422),
.A2(n_1429),
.B(n_1471),
.C(n_1470),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1466),
.A2(n_1413),
.B(n_1399),
.C(n_1420),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1451),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1399),
.A2(n_1451),
.B1(n_1484),
.B2(n_1435),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1401),
.B(n_1365),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1460),
.A2(n_1483),
.B(n_1477),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1401),
.B(n_1385),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1368),
.A2(n_1487),
.B(n_1445),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1452),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1435),
.B(n_1437),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1484),
.A2(n_1434),
.B1(n_1495),
.B2(n_1436),
.Y(n_1552)
);

O2A1O1Ixp5_ASAP7_75t_L g1553 ( 
.A1(n_1422),
.A2(n_1481),
.B(n_1447),
.C(n_1498),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1389),
.B(n_1468),
.Y(n_1554)
);

AOI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1384),
.A2(n_1439),
.B1(n_1426),
.B2(n_1436),
.C(n_1470),
.Y(n_1555)
);

INVxp33_ASAP7_75t_L g1556 ( 
.A(n_1438),
.Y(n_1556)
);

OA22x2_ASAP7_75t_L g1557 ( 
.A1(n_1434),
.A2(n_1475),
.B1(n_1432),
.B2(n_1378),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1463),
.B(n_1471),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1485),
.B(n_1492),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1432),
.B(n_1433),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1434),
.A2(n_1495),
.B1(n_1371),
.B2(n_1479),
.Y(n_1561)
);

OA22x2_ASAP7_75t_L g1562 ( 
.A1(n_1366),
.A2(n_1496),
.B1(n_1425),
.B2(n_1405),
.Y(n_1562)
);

O2A1O1Ixp5_ASAP7_75t_L g1563 ( 
.A1(n_1384),
.A2(n_1366),
.B(n_1496),
.C(n_1487),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1460),
.A2(n_1483),
.B(n_1469),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1495),
.A2(n_1496),
.B1(n_1491),
.B2(n_1444),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1493),
.B(n_1499),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1493),
.B(n_1499),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1499),
.B(n_1426),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1491),
.A2(n_1444),
.B1(n_1424),
.B2(n_1409),
.Y(n_1569)
);

AOI21x1_ASAP7_75t_SL g1570 ( 
.A1(n_1423),
.A2(n_1409),
.B(n_1407),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1426),
.B(n_1419),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1393),
.B(n_1406),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1419),
.B(n_1423),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1419),
.B(n_1424),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1381),
.A2(n_1377),
.B(n_1382),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1423),
.Y(n_1576)
);

AOI21x1_ASAP7_75t_SL g1577 ( 
.A1(n_1409),
.A2(n_1393),
.B(n_1382),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1390),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1462),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1377),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1376),
.A2(n_1308),
.B1(n_1324),
.B2(n_1465),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1376),
.A2(n_1308),
.B1(n_1324),
.B2(n_1465),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1381),
.A2(n_1458),
.B(n_1238),
.C(n_1362),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1414),
.B(n_1373),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1465),
.A2(n_1308),
.B1(n_1324),
.B2(n_1200),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_R g1586 ( 
.A(n_1472),
.B(n_846),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1387),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1448),
.A2(n_938),
.B(n_1106),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1367),
.B(n_1480),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1503),
.B(n_1504),
.Y(n_1590)
);

OR2x6_ASAP7_75t_L g1591 ( 
.A(n_1541),
.B(n_1525),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1568),
.B(n_1567),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1532),
.B(n_1537),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

INVxp67_ASAP7_75t_SL g1595 ( 
.A(n_1541),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1553),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1557),
.Y(n_1597)
);

AOI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1575),
.A2(n_1549),
.B(n_1538),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1546),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1535),
.B(n_1539),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1548),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1557),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1511),
.B(n_1509),
.Y(n_1603)
);

AOI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1585),
.A2(n_1512),
.B1(n_1507),
.B2(n_1588),
.C(n_1508),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1549),
.A2(n_1518),
.B(n_1538),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1505),
.B(n_1506),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1574),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1566),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_SL g1609 ( 
.A(n_1540),
.B(n_1513),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1573),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1512),
.B(n_1522),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1569),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1542),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1526),
.B(n_1589),
.Y(n_1615)
);

OR2x6_ASAP7_75t_L g1616 ( 
.A(n_1572),
.B(n_1543),
.Y(n_1616)
);

AOI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1580),
.A2(n_1531),
.B(n_1536),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1562),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1527),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1583),
.A2(n_1523),
.B(n_1581),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1576),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1514),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1501),
.B(n_1584),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1560),
.B(n_1529),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1528),
.A2(n_1523),
.B(n_1517),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1572),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1572),
.B(n_1579),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1516),
.Y(n_1628)
);

INVx5_ASAP7_75t_L g1629 ( 
.A(n_1533),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1515),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1555),
.B(n_1582),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1554),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1563),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1530),
.B(n_1520),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1555),
.B(n_1559),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_SL g1636 ( 
.A1(n_1510),
.A2(n_1521),
.B1(n_1519),
.B2(n_1552),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1613),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1593),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1601),
.B(n_1558),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1597),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1599),
.B(n_1603),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1603),
.B(n_1545),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1618),
.B(n_1564),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1622),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1597),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1605),
.A2(n_1516),
.B(n_1564),
.Y(n_1647)
);

OAI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1598),
.A2(n_1577),
.B(n_1570),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1627),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1618),
.B(n_1551),
.Y(n_1650)
);

INVx4_ASAP7_75t_L g1651 ( 
.A(n_1629),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1634),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1611),
.B(n_1561),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1610),
.B(n_1630),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1604),
.A2(n_1534),
.B1(n_1565),
.B2(n_1556),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1593),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1626),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1638),
.B(n_1612),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1651),
.B(n_1657),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1642),
.B(n_1619),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1653),
.A2(n_1604),
.B1(n_1620),
.B2(n_1625),
.C(n_1611),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1653),
.A2(n_1620),
.B1(n_1625),
.B2(n_1631),
.C(n_1590),
.Y(n_1662)
);

AOI211xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1643),
.A2(n_1631),
.B(n_1595),
.C(n_1612),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1600),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1651),
.B(n_1597),
.Y(n_1665)
);

NOR4xp25_ASAP7_75t_SL g1666 ( 
.A(n_1652),
.B(n_1595),
.C(n_1550),
.D(n_1502),
.Y(n_1666)
);

AOI222xp33_ASAP7_75t_L g1667 ( 
.A1(n_1643),
.A2(n_1609),
.B1(n_1652),
.B2(n_1623),
.C1(n_1635),
.C2(n_1642),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1641),
.A2(n_1636),
.B1(n_1591),
.B2(n_1602),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1638),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1641),
.A2(n_1636),
.B1(n_1591),
.B2(n_1602),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1641),
.A2(n_1591),
.B1(n_1602),
.B2(n_1646),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1638),
.A2(n_1633),
.B1(n_1623),
.B2(n_1635),
.C(n_1606),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_R g1673 ( 
.A(n_1650),
.B(n_1500),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1654),
.B(n_1600),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1654),
.B(n_1649),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1637),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1655),
.A2(n_1591),
.B1(n_1628),
.B2(n_1629),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1651),
.Y(n_1679)
);

INVx4_ASAP7_75t_L g1680 ( 
.A(n_1651),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1637),
.Y(n_1681)
);

AOI31xp33_ASAP7_75t_L g1682 ( 
.A1(n_1655),
.A2(n_1609),
.A3(n_1614),
.B(n_1615),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_SL g1683 ( 
.A(n_1651),
.B(n_1586),
.Y(n_1683)
);

OA222x2_ASAP7_75t_L g1684 ( 
.A1(n_1646),
.A2(n_1616),
.B1(n_1614),
.B2(n_1621),
.C1(n_1608),
.C2(n_1607),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1646),
.A2(n_1655),
.B1(n_1650),
.B2(n_1624),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1654),
.B(n_1649),
.Y(n_1686)
);

NOR3xp33_ASAP7_75t_L g1687 ( 
.A(n_1647),
.B(n_1617),
.C(n_1587),
.Y(n_1687)
);

NAND4xp25_ASAP7_75t_L g1688 ( 
.A(n_1647),
.B(n_1614),
.C(n_1544),
.D(n_1632),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1648),
.A2(n_1596),
.B(n_1594),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1656),
.B(n_1621),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1644),
.A2(n_1632),
.B(n_1627),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1646),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1667),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1674),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1674),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1677),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1676),
.B(n_1639),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_L g1699 ( 
.A(n_1661),
.B(n_1524),
.C(n_1651),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1639),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1677),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1681),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1692),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1667),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1659),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1689),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1686),
.B(n_1639),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1680),
.Y(n_1708)
);

INVx3_ASAP7_75t_L g1709 ( 
.A(n_1679),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1669),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1687),
.A2(n_1691),
.B(n_1645),
.Y(n_1712)
);

BUFx8_ASAP7_75t_L g1713 ( 
.A(n_1679),
.Y(n_1713)
);

INVx4_ASAP7_75t_SL g1714 ( 
.A(n_1679),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1690),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1714),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1695),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1706),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1714),
.B(n_1664),
.Y(n_1719)
);

NAND3xp33_ASAP7_75t_L g1720 ( 
.A(n_1694),
.B(n_1662),
.C(n_1663),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1714),
.B(n_1664),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1714),
.B(n_1705),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1694),
.B(n_1672),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1699),
.B(n_1683),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1713),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1695),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1704),
.B(n_1660),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1706),
.Y(n_1728)
);

INVxp67_ASAP7_75t_L g1729 ( 
.A(n_1711),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1670),
.C(n_1668),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1715),
.B(n_1658),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1699),
.B(n_1682),
.Y(n_1733)
);

NAND2x1p5_ASAP7_75t_L g1734 ( 
.A(n_1712),
.B(n_1651),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1698),
.B(n_1684),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1706),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1711),
.B(n_1693),
.Y(n_1737)
);

NAND4xp25_ASAP7_75t_L g1738 ( 
.A(n_1708),
.B(n_1678),
.C(n_1685),
.D(n_1688),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1695),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1714),
.B(n_1686),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1709),
.B(n_1682),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1703),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1696),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1705),
.B(n_1665),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1703),
.B(n_1690),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1698),
.B(n_1684),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1697),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1713),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1713),
.B(n_1673),
.Y(n_1750)
);

NAND2xp33_ASAP7_75t_R g1751 ( 
.A(n_1725),
.B(n_1666),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1723),
.B(n_1701),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1743),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1719),
.B(n_1709),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1720),
.A2(n_1688),
.B1(n_1712),
.B2(n_1671),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1744),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1744),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1700),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1719),
.B(n_1709),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1748),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1748),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1721),
.B(n_1709),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1721),
.B(n_1708),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1746),
.B(n_1712),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1723),
.B(n_1701),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1746),
.B(n_1712),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1727),
.B(n_1702),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1727),
.B(n_1708),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1730),
.B(n_1710),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1717),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1730),
.B(n_1710),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1740),
.B(n_1710),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1718),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1717),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1733),
.B(n_1713),
.Y(n_1775)
);

NAND2x1_ASAP7_75t_L g1776 ( 
.A(n_1716),
.B(n_1712),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1731),
.B(n_1700),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1740),
.B(n_1707),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1718),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1726),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1729),
.B(n_1702),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1726),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1741),
.B(n_1707),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1731),
.B(n_1707),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1718),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1728),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1729),
.B(n_1702),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1783),
.B(n_1716),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1773),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1776),
.A2(n_1734),
.B(n_1722),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1775),
.A2(n_1724),
.B1(n_1738),
.B2(n_1742),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1776),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1777),
.A2(n_1738),
.B1(n_1712),
.B2(n_1749),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1753),
.B(n_1743),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1773),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1763),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1783),
.B(n_1716),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1756),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1756),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1763),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1757),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1778),
.B(n_1716),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1757),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1760),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1760),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1761),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1761),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1758),
.B(n_1739),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1778),
.B(n_1722),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1773),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1784),
.A2(n_1755),
.B(n_1752),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1752),
.B(n_1737),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1765),
.B(n_1737),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1779),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1798),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1793),
.A2(n_1755),
.B1(n_1751),
.B2(n_1768),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1791),
.A2(n_1765),
.B1(n_1767),
.B2(n_1747),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1793),
.B(n_1725),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1798),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1811),
.A2(n_1767),
.B(n_1734),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1794),
.Y(n_1821)
);

OAI32xp33_ASAP7_75t_L g1822 ( 
.A1(n_1796),
.A2(n_1800),
.A3(n_1794),
.B1(n_1812),
.B2(n_1813),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1788),
.B(n_1749),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1788),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1811),
.A2(n_1747),
.B1(n_1735),
.B2(n_1769),
.Y(n_1825)
);

NAND4xp25_ASAP7_75t_L g1826 ( 
.A(n_1796),
.B(n_1769),
.C(n_1771),
.D(n_1772),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1800),
.B(n_1732),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1809),
.B(n_1771),
.Y(n_1828)
);

NOR3xp33_ASAP7_75t_L g1829 ( 
.A(n_1812),
.B(n_1813),
.C(n_1801),
.Y(n_1829)
);

AOI21xp33_ASAP7_75t_L g1830 ( 
.A1(n_1808),
.A2(n_1772),
.B(n_1781),
.Y(n_1830)
);

AOI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1808),
.A2(n_1787),
.B(n_1781),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_SL g1832 ( 
.A1(n_1788),
.A2(n_1802),
.B1(n_1797),
.B2(n_1809),
.Y(n_1832)
);

OAI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1808),
.A2(n_1734),
.B1(n_1764),
.B2(n_1766),
.C(n_1750),
.Y(n_1833)
);

OAI222xp33_ASAP7_75t_L g1834 ( 
.A1(n_1797),
.A2(n_1734),
.B1(n_1766),
.B2(n_1764),
.C1(n_1747),
.C2(n_1735),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1809),
.B(n_1754),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1799),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1824),
.B(n_1797),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1828),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1815),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1819),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1827),
.Y(n_1841)
);

NOR2x1_ASAP7_75t_L g1842 ( 
.A(n_1818),
.B(n_1792),
.Y(n_1842)
);

INVxp67_ASAP7_75t_L g1843 ( 
.A(n_1823),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1828),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1835),
.B(n_1802),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1836),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1821),
.B(n_1799),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1835),
.B(n_1802),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1816),
.A2(n_1741),
.B1(n_1666),
.B2(n_1735),
.Y(n_1849)
);

NOR3xp33_ASAP7_75t_L g1850 ( 
.A(n_1843),
.B(n_1818),
.C(n_1822),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1842),
.A2(n_1820),
.B(n_1829),
.C(n_1830),
.Y(n_1851)
);

OAI211xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1841),
.A2(n_1817),
.B(n_1825),
.C(n_1831),
.Y(n_1852)
);

O2A1O1Ixp33_ASAP7_75t_L g1853 ( 
.A1(n_1847),
.A2(n_1826),
.B(n_1817),
.C(n_1833),
.Y(n_1853)
);

NOR3xp33_ASAP7_75t_L g1854 ( 
.A(n_1837),
.B(n_1832),
.C(n_1803),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1844),
.A2(n_1825),
.B(n_1834),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1845),
.B(n_1801),
.Y(n_1856)
);

AOI211xp5_ASAP7_75t_L g1857 ( 
.A1(n_1849),
.A2(n_1805),
.B(n_1803),
.C(n_1804),
.Y(n_1857)
);

AOI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1845),
.A2(n_1754),
.B1(n_1762),
.B2(n_1759),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_SL g1859 ( 
.A(n_1838),
.B(n_1759),
.Y(n_1859)
);

AOI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1847),
.A2(n_1848),
.B(n_1839),
.C(n_1840),
.Y(n_1860)
);

AOI31xp33_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1846),
.A3(n_1848),
.B(n_1804),
.Y(n_1861)
);

OAI21xp33_ASAP7_75t_L g1862 ( 
.A1(n_1859),
.A2(n_1806),
.B(n_1805),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1854),
.B(n_1806),
.Y(n_1863)
);

AOI221x1_ASAP7_75t_SL g1864 ( 
.A1(n_1857),
.A2(n_1807),
.B1(n_1810),
.B2(n_1814),
.C(n_1795),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1856),
.Y(n_1865)
);

AOI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1850),
.A2(n_1807),
.B1(n_1762),
.B2(n_1792),
.Y(n_1866)
);

OAI311xp33_ASAP7_75t_L g1867 ( 
.A1(n_1855),
.A2(n_1792),
.A3(n_1787),
.B1(n_1782),
.C1(n_1774),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1866),
.B(n_1858),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1862),
.Y(n_1869)
);

NOR2x1_ASAP7_75t_L g1870 ( 
.A(n_1863),
.B(n_1861),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1863),
.B(n_1853),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1865),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1864),
.Y(n_1873)
);

AOI211xp5_ASAP7_75t_L g1874 ( 
.A1(n_1871),
.A2(n_1867),
.B(n_1851),
.C(n_1852),
.Y(n_1874)
);

OAI21xp33_ASAP7_75t_L g1875 ( 
.A1(n_1871),
.A2(n_1792),
.B(n_1789),
.Y(n_1875)
);

NOR2x1_ASAP7_75t_L g1876 ( 
.A(n_1870),
.B(n_1789),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1868),
.B(n_1789),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1869),
.B(n_1745),
.Y(n_1878)
);

XOR2xp5_ASAP7_75t_L g1879 ( 
.A(n_1878),
.B(n_1873),
.Y(n_1879)
);

NAND2xp33_ASAP7_75t_SL g1880 ( 
.A(n_1877),
.B(n_1872),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1876),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1879),
.B(n_1874),
.Y(n_1882)
);

OAI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1882),
.A2(n_1880),
.B1(n_1875),
.B2(n_1881),
.C(n_1810),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1883),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1883),
.A2(n_1814),
.B1(n_1810),
.B2(n_1795),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1885),
.A2(n_1884),
.B1(n_1814),
.B2(n_1795),
.C(n_1779),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1884),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_SL g1888 ( 
.A1(n_1887),
.A2(n_1782),
.B1(n_1780),
.B2(n_1774),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1886),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1889),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1890),
.B(n_1888),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_SL g1892 ( 
.A1(n_1891),
.A2(n_1780),
.B(n_1770),
.Y(n_1892)
);

AOI22xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1892),
.A2(n_1770),
.B1(n_1785),
.B2(n_1779),
.Y(n_1893)
);

AOI221xp5_ASAP7_75t_L g1894 ( 
.A1(n_1893),
.A2(n_1785),
.B1(n_1786),
.B2(n_1728),
.C(n_1736),
.Y(n_1894)
);

AOI211xp5_ASAP7_75t_L g1895 ( 
.A1(n_1894),
.A2(n_1790),
.B(n_1786),
.C(n_1785),
.Y(n_1895)
);


endmodule