module fake_jpeg_542_n_672 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_672);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_672;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_59),
.B(n_62),
.Y(n_148)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_17),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_64),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_65),
.B(n_70),
.Y(n_156)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

INVx11_ASAP7_75t_SL g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_16),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_20),
.B(n_0),
.CON(n_71),
.SN(n_71)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_71),
.B(n_119),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_81),
.Y(n_158)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_76),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_84),
.B(n_93),
.Y(n_179)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_86),
.Y(n_166)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_0),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_90),
.Y(n_203)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_94),
.B(n_99),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_98),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_96),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_97),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_37),
.B(n_1),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_100),
.Y(n_186)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_105),
.B(n_117),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_106),
.B(n_110),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_45),
.B(n_15),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_107),
.B(n_122),
.C(n_53),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_108),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_49),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_49),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_112),
.B(n_116),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_113),
.Y(n_229)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_51),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_51),
.B(n_34),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

BUFx12f_ASAP7_75t_SL g119 ( 
.A(n_34),
.Y(n_119)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_51),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_121),
.B(n_125),
.Y(n_220)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_24),
.B(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_43),
.B(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_123),
.B(n_124),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_43),
.B(n_27),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_25),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_38),
.Y(n_126)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_38),
.Y(n_127)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_41),
.Y(n_128)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_128),
.Y(n_215)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_41),
.B(n_27),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_30),
.Y(n_145)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_41),
.Y(n_131)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_30),
.B1(n_53),
.B2(n_44),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_132),
.B(n_109),
.Y(n_276)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_133),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_33),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_134),
.B(n_216),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_80),
.B1(n_119),
.B2(n_126),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_142),
.A2(n_147),
.B1(n_226),
.B2(n_71),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_88),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_144),
.B(n_170),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_145),
.B(n_120),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_25),
.B1(n_32),
.B2(n_39),
.Y(n_147)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_67),
.Y(n_170)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_107),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_178),
.B(n_180),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_107),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_113),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_184),
.B(n_190),
.Y(n_303)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_61),
.Y(n_187)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_122),
.B(n_40),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_228),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_129),
.Y(n_190)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

OR2x2_ASAP7_75t_SL g261 ( 
.A(n_195),
.B(n_196),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_117),
.A2(n_39),
.B(n_32),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_78),
.B(n_40),
.C(n_44),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_199),
.B(n_10),
.Y(n_313)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_83),
.Y(n_204)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_73),
.Y(n_207)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_208),
.Y(n_260)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_74),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_77),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_104),
.Y(n_213)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_115),
.B(n_36),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_69),
.Y(n_217)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_76),
.Y(n_218)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_79),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_221),
.B(n_5),
.Y(n_304)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_64),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_111),
.Y(n_225)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_103),
.A2(n_38),
.B1(n_36),
.B2(n_33),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_87),
.Y(n_227)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_66),
.B(n_4),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_135),
.Y(n_233)
);

INVx11_ASAP7_75t_L g377 ( 
.A(n_233),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_168),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_234),
.B(n_247),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_236),
.Y(n_332)
);

CKINVDCx12_ASAP7_75t_R g237 ( 
.A(n_164),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_237),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_181),
.A2(n_97),
.B1(n_89),
.B2(n_90),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_242),
.A2(n_309),
.B1(n_173),
.B2(n_159),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_142),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_243),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_168),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_136),
.Y(n_248)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_248),
.Y(n_362)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_136),
.Y(n_253)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_253),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_148),
.B(n_128),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_255),
.B(n_267),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_259),
.Y(n_351)
);

XNOR2x1_ASAP7_75t_SL g341 ( 
.A(n_262),
.B(n_313),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_141),
.Y(n_263)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_263),
.Y(n_364)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_160),
.Y(n_266)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_151),
.B(n_118),
.Y(n_267)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_164),
.Y(n_270)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_270),
.Y(n_334)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_164),
.Y(n_271)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_143),
.Y(n_272)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_272),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_153),
.B(n_4),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_273),
.B(n_275),
.Y(n_373)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_143),
.Y(n_274)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_220),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_276),
.B(n_289),
.Y(n_360)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_223),
.A2(n_100),
.B(n_63),
.C(n_57),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_315),
.Y(n_322)
);

AOI32xp33_ASAP7_75t_L g278 ( 
.A1(n_156),
.A2(n_194),
.A3(n_179),
.B1(n_206),
.B2(n_162),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_278),
.B(n_294),
.Y(n_348)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_158),
.Y(n_279)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_209),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_287),
.Y(n_320)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_152),
.Y(n_283)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_283),
.Y(n_358)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_171),
.Y(n_285)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_285),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_201),
.Y(n_286)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_286),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_137),
.B(n_5),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_139),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_292),
.Y(n_333)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_152),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_146),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_291),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_229),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_167),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_295),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_197),
.A2(n_96),
.B1(n_57),
.B2(n_56),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_177),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_192),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_298),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_166),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_297),
.A2(n_300),
.B1(n_312),
.B2(n_314),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_154),
.B(n_163),
.Y(n_298)
);

CKINVDCx9p33_ASAP7_75t_R g299 ( 
.A(n_166),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_299),
.Y(n_346)
);

INVx11_ASAP7_75t_L g300 ( 
.A(n_138),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_169),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_301),
.B(n_304),
.Y(n_349)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_191),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_302),
.B(n_307),
.Y(n_378)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_192),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_305),
.B(n_306),
.Y(n_376)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_157),
.B(n_161),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_193),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_308),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_165),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_226),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_310),
.A2(n_207),
.B1(n_224),
.B2(n_219),
.Y(n_339)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_191),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_311),
.Y(n_365)
);

INVx11_ASAP7_75t_L g312 ( 
.A(n_138),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_186),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_198),
.B(n_11),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_212),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_316),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_140),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_319),
.B(n_328),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_264),
.B(n_215),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_321),
.B(n_345),
.C(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_174),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_324),
.B(n_343),
.Y(n_398)
);

AND2x4_ASAP7_75t_SL g325 ( 
.A(n_262),
.B(n_261),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_325),
.B(n_274),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_326),
.A2(n_338),
.B1(n_350),
.B2(n_356),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_243),
.A2(n_140),
.B1(n_202),
.B2(n_147),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_254),
.A2(n_176),
.B1(n_224),
.B2(n_219),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_330),
.A2(n_331),
.B1(n_339),
.B2(n_353),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_236),
.A2(n_210),
.B1(n_211),
.B2(n_133),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_276),
.A2(n_183),
.B1(n_182),
.B2(n_174),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_149),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_239),
.B(n_183),
.C(n_182),
.Y(n_345)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_231),
.B(n_149),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_302),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_251),
.A2(n_155),
.B1(n_203),
.B2(n_189),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_277),
.A2(n_155),
.B1(n_203),
.B2(n_189),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_249),
.A2(n_150),
.B1(n_176),
.B2(n_172),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_355),
.A2(n_312),
.B1(n_300),
.B2(n_291),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_303),
.A2(n_146),
.B1(n_172),
.B2(n_150),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_250),
.B(n_229),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_366),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_314),
.A2(n_200),
.B1(n_13),
.B2(n_14),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_245),
.B1(n_235),
.B2(n_285),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_265),
.B(n_12),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_260),
.B(n_12),
.C(n_13),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_258),
.B(n_12),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_369),
.A2(n_297),
.B(n_245),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_238),
.B(n_13),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_370),
.B(n_372),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_240),
.B(n_14),
.Y(n_372)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_380),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_364),
.Y(n_381)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_376),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_382),
.B(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_383),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_373),
.B(n_290),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_335),
.B(n_257),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_388),
.B(n_407),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_325),
.B(n_269),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_390),
.B(n_399),
.C(n_421),
.Y(n_441)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_317),
.Y(n_391)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_391),
.Y(n_436)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_392),
.Y(n_438)
);

OAI21xp33_ASAP7_75t_SL g460 ( 
.A1(n_393),
.A2(n_409),
.B(n_411),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_394),
.A2(n_417),
.B(n_369),
.Y(n_452)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_395),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_332),
.A2(n_246),
.B1(n_232),
.B2(n_252),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_396),
.A2(n_400),
.B1(n_329),
.B2(n_356),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_397),
.B(n_408),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_324),
.C(n_321),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_332),
.A2(n_246),
.B1(n_232),
.B2(n_252),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_322),
.A2(n_280),
.B1(n_244),
.B2(n_311),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_402),
.A2(n_339),
.B1(n_365),
.B2(n_345),
.Y(n_457)
);

OAI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_403),
.A2(n_328),
.B1(n_368),
.B2(n_346),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_404),
.Y(n_443)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_323),
.B(n_268),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_406),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_378),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_323),
.B(n_320),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_325),
.B(n_282),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_419),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_349),
.B(n_268),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_318),
.Y(n_412)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_342),
.A2(n_295),
.B1(n_263),
.B2(n_259),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_414),
.A2(n_415),
.B1(n_423),
.B2(n_425),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_342),
.A2(n_256),
.B1(n_284),
.B2(n_233),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_360),
.A2(n_235),
.B(n_284),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_416),
.A2(n_360),
.B(n_346),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_341),
.A2(n_233),
.B(n_241),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_344),
.Y(n_418)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_418),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_335),
.B(n_244),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_366),
.B(n_256),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_426),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_325),
.B(n_280),
.C(n_241),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_352),
.B(n_248),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_422),
.B(n_424),
.C(n_358),
.Y(n_467)
);

INVx13_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_319),
.B(n_347),
.C(n_322),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_344),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_347),
.B(n_253),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_427),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_428),
.B(n_446),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_431),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_360),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_437),
.B(n_456),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_386),
.A2(n_353),
.B1(n_348),
.B2(n_319),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_439),
.A2(n_457),
.B1(n_466),
.B2(n_390),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_389),
.A2(n_331),
.B1(n_326),
.B2(n_329),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_445),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_343),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_448),
.B(n_387),
.C(n_424),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_452),
.A2(n_453),
.B(n_374),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_409),
.A2(n_348),
.B(n_369),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_398),
.B(n_338),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_397),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_458),
.B(n_357),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_386),
.A2(n_350),
.B1(n_363),
.B2(n_365),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_459),
.A2(n_463),
.B1(n_469),
.B2(n_418),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_413),
.B(n_370),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_462),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_413),
.B(n_372),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_380),
.A2(n_369),
.B1(n_327),
.B2(n_362),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_351),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_465),
.B(n_412),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_379),
.A2(n_402),
.B1(n_401),
.B2(n_410),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_422),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_401),
.B(n_357),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_383),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_379),
.A2(n_383),
.B1(n_409),
.B2(n_420),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_432),
.Y(n_470)
);

NOR3xp33_ASAP7_75t_L g516 ( 
.A(n_470),
.B(n_486),
.C(n_491),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_471),
.B(n_480),
.C(n_448),
.Y(n_540)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_472),
.Y(n_514)
);

BUFx5_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_473),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_395),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_474),
.B(n_478),
.Y(n_518)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_476),
.Y(n_524)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_477),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_405),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_479),
.B(n_488),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_392),
.Y(n_481)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_481),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_456),
.A2(n_421),
.B1(n_379),
.B2(n_387),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_483),
.A2(n_441),
.B1(n_480),
.B2(n_485),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_391),
.Y(n_484)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_484),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_485),
.A2(n_499),
.B1(n_507),
.B2(n_463),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_455),
.Y(n_486)
);

O2A1O1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_435),
.A2(n_394),
.B(n_409),
.C(n_393),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_462),
.Y(n_489)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_489),
.Y(n_542)
);

OAI21xp33_ASAP7_75t_L g492 ( 
.A1(n_452),
.A2(n_416),
.B(n_396),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_L g544 ( 
.A1(n_492),
.A2(n_436),
.B(n_433),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_334),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_494),
.B(n_503),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_495),
.A2(n_500),
.B1(n_506),
.B2(n_438),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_434),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_496),
.B(n_498),
.Y(n_530)
);

AND2x4_ASAP7_75t_SL g510 ( 
.A(n_497),
.B(n_469),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_429),
.B(n_426),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_439),
.A2(n_400),
.B1(n_385),
.B2(n_381),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_456),
.A2(n_351),
.B1(n_375),
.B2(n_364),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_465),
.A2(n_359),
.B(n_423),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_501),
.A2(n_508),
.B(n_453),
.Y(n_536)
);

CKINVDCx12_ASAP7_75t_R g502 ( 
.A(n_443),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_502),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_447),
.B(n_334),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_454),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_504),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_460),
.B(n_375),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_444),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_459),
.A2(n_358),
.B1(n_371),
.B2(n_359),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_457),
.A2(n_371),
.B1(n_337),
.B2(n_374),
.Y(n_507)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_509),
.Y(n_548)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_510),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_470),
.B(n_447),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_512),
.B(n_523),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_513),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_515),
.B(n_488),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_517),
.A2(n_525),
.B1(n_543),
.B2(n_500),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_471),
.B(n_441),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_519),
.B(n_508),
.Y(n_556)
);

OA21x2_ASAP7_75t_SL g523 ( 
.A1(n_475),
.A2(n_435),
.B(n_429),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_482),
.A2(n_465),
.B1(n_437),
.B2(n_428),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_497),
.A2(n_493),
.B(n_505),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_526),
.A2(n_529),
.B(n_535),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_493),
.A2(n_437),
.B(n_444),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_481),
.B(n_454),
.Y(n_531)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_531),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_496),
.B(n_430),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_532),
.B(n_489),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_484),
.B(n_443),
.Y(n_533)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_533),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_491),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_534),
.B(n_487),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_493),
.A2(n_466),
.B(n_446),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_536),
.A2(n_544),
.B(n_337),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_486),
.B(n_438),
.Y(n_537)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_537),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_540),
.B(n_541),
.C(n_502),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_483),
.B(n_467),
.C(n_440),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_482),
.A2(n_440),
.B1(n_464),
.B2(n_436),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_475),
.B(n_433),
.Y(n_545)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_545),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_518),
.B(n_477),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_547),
.B(n_564),
.Y(n_593)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_527),
.Y(n_549)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_549),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_527),
.Y(n_551)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_551),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_528),
.A2(n_487),
.B1(n_499),
.B2(n_490),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_552),
.A2(n_562),
.B1(n_563),
.B2(n_510),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_553),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_554),
.A2(n_560),
.B1(n_509),
.B2(n_525),
.Y(n_576)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_555),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_556),
.B(n_541),
.C(n_515),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_558),
.B(n_561),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_517),
.A2(n_495),
.B1(n_490),
.B2(n_505),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_540),
.B(n_479),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_528),
.A2(n_501),
.B1(n_507),
.B2(n_498),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_538),
.A2(n_472),
.B1(n_504),
.B2(n_476),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_518),
.B(n_451),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_534),
.B(n_506),
.Y(n_565)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_565),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_567),
.B(n_574),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_539),
.B(n_367),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_568),
.B(n_571),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_539),
.B(n_473),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_573),
.A2(n_536),
.B(n_513),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_SL g574 ( 
.A(n_519),
.B(n_377),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_531),
.B(n_15),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_575),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_576),
.A2(n_579),
.B1(n_589),
.B2(n_598),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_550),
.B(n_521),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_577),
.B(n_587),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_554),
.A2(n_538),
.B1(n_542),
.B2(n_511),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_561),
.B(n_567),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_583),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_586),
.B(n_559),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_568),
.B(n_521),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_548),
.A2(n_542),
.B1(n_511),
.B2(n_535),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_590),
.A2(n_594),
.B1(n_569),
.B2(n_559),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_558),
.B(n_529),
.C(n_526),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_591),
.B(n_596),
.C(n_600),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_592),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_548),
.A2(n_543),
.B1(n_537),
.B2(n_510),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_556),
.B(n_513),
.C(n_523),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g598 ( 
.A1(n_560),
.A2(n_570),
.B1(n_557),
.B2(n_572),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_566),
.B(n_522),
.Y(n_599)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_599),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_574),
.B(n_545),
.C(n_522),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_584),
.B(n_553),
.Y(n_601)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_601),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_602),
.B(n_605),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_603),
.B(n_611),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_573),
.Y(n_605)
);

A2O1A1O1Ixp25_ASAP7_75t_L g609 ( 
.A1(n_591),
.A2(n_516),
.B(n_570),
.C(n_557),
.D(n_566),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_609),
.A2(n_592),
.B(n_590),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_585),
.B(n_530),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_613),
.Y(n_623)
);

OAI21x1_ASAP7_75t_SL g611 ( 
.A1(n_595),
.A2(n_530),
.B(n_565),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_580),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_612),
.B(n_571),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_593),
.B(n_549),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_595),
.B(n_520),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_614),
.B(n_618),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_579),
.B(n_533),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_615),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_581),
.B(n_546),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_616),
.B(n_588),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_583),
.B(n_546),
.C(n_562),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_598),
.B(n_578),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_620),
.B(n_589),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_619),
.A2(n_609),
.B(n_601),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_621),
.A2(n_630),
.B(n_635),
.Y(n_645)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_625),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_607),
.B(n_586),
.C(n_582),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_627),
.B(n_629),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_604),
.B(n_563),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_619),
.A2(n_617),
.B(n_594),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g648 ( 
.A1(n_631),
.A2(n_510),
.B(n_514),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_602),
.B(n_582),
.C(n_600),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_633),
.B(n_637),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_634),
.B(n_575),
.Y(n_641)
);

NOR2xp67_ASAP7_75t_SL g635 ( 
.A(n_608),
.B(n_596),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_636),
.B(n_616),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_608),
.B(n_552),
.C(n_578),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_621),
.A2(n_617),
.B1(n_615),
.B2(n_603),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_638),
.B(n_642),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_641),
.B(n_643),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_627),
.B(n_618),
.C(n_605),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_637),
.B(n_633),
.C(n_626),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_644),
.B(n_646),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_626),
.B(n_606),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_631),
.B(n_597),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g652 ( 
.A(n_647),
.B(n_628),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_648),
.A2(n_630),
.B(n_629),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_650),
.B(n_652),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_645),
.A2(n_624),
.B(n_623),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_654),
.B(n_656),
.Y(n_658)
);

XNOR2x1_ASAP7_75t_SL g656 ( 
.A(n_646),
.B(n_628),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_644),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_657),
.B(n_643),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_651),
.B(n_649),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_660),
.B(n_662),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_655),
.B(n_639),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_661),
.B(n_653),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_658),
.A2(n_645),
.B(n_640),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_664),
.A2(n_659),
.B(n_638),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_665),
.B(n_632),
.Y(n_667)
);

AO21x2_ASAP7_75t_L g668 ( 
.A1(n_666),
.A2(n_667),
.B(n_663),
.Y(n_668)
);

AOI322xp5_ASAP7_75t_L g669 ( 
.A1(n_668),
.A2(n_622),
.A3(n_648),
.B1(n_524),
.B2(n_514),
.C1(n_642),
.C2(n_636),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_669),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_670),
.A2(n_524),
.B(n_597),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_L g672 ( 
.A(n_671),
.B(n_377),
.Y(n_672)
);


endmodule