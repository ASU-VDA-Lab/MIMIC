module fake_jpeg_24273_n_231 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_32),
.Y(n_45)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_13),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_51),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_46),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_44),
.B1(n_20),
.B2(n_14),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_26),
.B1(n_16),
.B2(n_21),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_50),
.B1(n_31),
.B2(n_35),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_17),
.B1(n_24),
.B2(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_26),
.B1(n_16),
.B2(n_21),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_22),
.C(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_54),
.Y(n_78)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_59),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_35),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_65),
.B(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_64),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_27),
.B1(n_28),
.B2(n_14),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_34),
.B1(n_29),
.B2(n_32),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_34),
.B1(n_51),
.B2(n_13),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_31),
.B1(n_34),
.B2(n_29),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_50),
.B1(n_40),
.B2(n_31),
.Y(n_84)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_68),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_57),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_19),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_33),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_59),
.B1(n_48),
.B2(n_28),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_55),
.B1(n_71),
.B2(n_47),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_58),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_60),
.C(n_61),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_107),
.C(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_103),
.B1(n_108),
.B2(n_111),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_100),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_60),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_80),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_69),
.B(n_66),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_89),
.B(n_85),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_49),
.C(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_75),
.B(n_30),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_23),
.Y(n_111)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_116),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_79),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_128),
.C(n_130),
.Y(n_133)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_77),
.B1(n_73),
.B2(n_72),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_R g122 ( 
.A1(n_102),
.A2(n_73),
.B(n_77),
.C(n_81),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_123),
.B(n_43),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_85),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_84),
.B1(n_47),
.B2(n_48),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_47),
.B1(n_41),
.B2(n_31),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_107),
.C(n_104),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_31),
.B1(n_28),
.B2(n_63),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_130),
.C(n_115),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_143),
.C(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_148),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_141),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_86),
.C(n_88),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_108),
.B1(n_91),
.B2(n_68),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_144),
.A2(n_27),
.B1(n_38),
.B2(n_26),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_108),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_151),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_33),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_162),
.C(n_133),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_120),
.B1(n_38),
.B2(n_28),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_143),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_137),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_27),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_33),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_179),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_146),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_162),
.C(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_140),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_132),
.B1(n_150),
.B2(n_134),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_182),
.B1(n_161),
.B2(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_166),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_133),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_191),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_193),
.B(n_173),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_146),
.C(n_152),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_161),
.B1(n_158),
.B2(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_174),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_168),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_181),
.B(n_157),
.C(n_173),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_196),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_176),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_199),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_200),
.C(n_201),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_168),
.C(n_171),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_160),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_151),
.C(n_4),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_194),
.C(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_210),
.C(n_211),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_202),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_185),
.C(n_169),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_215),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_203),
.B(n_196),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_8),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_5),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_8),
.B(n_4),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_5),
.B(n_7),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_8),
.B(n_4),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_222),
.C(n_218),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_5),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_225),
.B(n_7),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_9),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.C(n_9),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_9),
.B1(n_11),
.B2(n_1),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_11),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_33),
.B(n_226),
.Y(n_231)
);


endmodule