module fake_jpeg_22154_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_38),
.Y(n_46)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_25),
.B1(n_15),
.B2(n_28),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_2),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp67_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_23),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_19),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_57),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_23),
.B(n_29),
.C(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_54),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_30),
.B(n_23),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_56),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_29),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_37),
.B(n_33),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_28),
.B1(n_21),
.B2(n_29),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_32),
.A2(n_25),
.B1(n_26),
.B2(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_26),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_17),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_71),
.Y(n_98)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_62),
.B1(n_57),
.B2(n_45),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_21),
.B1(n_44),
.B2(n_16),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_45),
.B1(n_68),
.B2(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_4),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_4),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_5),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_46),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_89),
.B1(n_83),
.B2(n_91),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_75),
.B1(n_71),
.B2(n_45),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_51),
.C(n_46),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_101),
.C(n_100),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_119),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_116),
.B1(n_80),
.B2(n_97),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_118),
.C(n_120),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_84),
.B(n_70),
.C(n_80),
.D(n_48),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_84),
.C(n_73),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_84),
.C(n_73),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_124),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_80),
.B(n_72),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_110),
.B(n_106),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_50),
.C(n_72),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_48),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_132),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_134),
.B(n_135),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_93),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_115),
.C(n_126),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_111),
.B(n_94),
.Y(n_134)
);

AOI222xp33_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_111),
.B1(n_94),
.B2(n_96),
.C1(n_95),
.C2(n_90),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_124),
.B1(n_122),
.B2(n_120),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_133),
.B1(n_137),
.B2(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_145),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.C(n_144),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_97),
.C(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_129),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_50),
.C(n_68),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_150),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_146),
.Y(n_150)
);

AOI31xp67_ASAP7_75t_SL g155 ( 
.A1(n_151),
.A2(n_85),
.A3(n_16),
.B(n_55),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_95),
.B1(n_104),
.B2(n_77),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_102),
.B1(n_119),
.B2(n_5),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_140),
.A3(n_141),
.B1(n_144),
.B2(n_119),
.C1(n_55),
.C2(n_85),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_157),
.C(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_11),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_147),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.C(n_157),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.C(n_6),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_12),
.C(n_5),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_6),
.Y(n_164)
);


endmodule