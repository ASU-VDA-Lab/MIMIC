module fake_jpeg_20803_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_62),
.Y(n_85)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_17),
.B1(n_16),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_28),
.B1(n_42),
.B2(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_23),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_73),
.A2(n_94),
.B1(n_87),
.B2(n_99),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_79),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_39),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_50),
.C(n_48),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_28),
.B1(n_31),
.B2(n_16),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_21),
.A3(n_29),
.B1(n_22),
.B2(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_99),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_31),
.B1(n_28),
.B2(n_37),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_92),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_139)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_46),
.B1(n_44),
.B2(n_41),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_95),
.B(n_96),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_106),
.Y(n_149)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_59),
.A2(n_42),
.B1(n_37),
.B2(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_20),
.B1(n_26),
.B2(n_34),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_60),
.A2(n_20),
.B1(n_26),
.B2(n_34),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_67),
.A2(n_49),
.B(n_15),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_19),
.C(n_33),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_111),
.A2(n_113),
.B1(n_49),
.B2(n_20),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_32),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_94),
.B1(n_80),
.B2(n_75),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_146),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_123),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_73),
.A2(n_22),
.B(n_23),
.C(n_36),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_132),
.B(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_85),
.B(n_35),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_141),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_48),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_131),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_43),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_84),
.A2(n_25),
.B1(n_29),
.B2(n_22),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_43),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_27),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_93),
.A2(n_25),
.B1(n_19),
.B2(n_33),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_88),
.B(n_33),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_95),
.B(n_96),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_88),
.B(n_105),
.C(n_101),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_19),
.B1(n_33),
.B2(n_27),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_150),
.A2(n_154),
.B1(n_168),
.B2(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_75),
.B1(n_77),
.B2(n_82),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_162),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_157),
.B(n_180),
.Y(n_204)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_77),
.A3(n_89),
.B1(n_81),
.B2(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_179),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_100),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_4),
.B(n_5),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_119),
.C(n_128),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_169),
.C(n_144),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_97),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_173),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_103),
.B1(n_90),
.B2(n_100),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_170),
.B1(n_177),
.B2(n_178),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_112),
.B1(n_113),
.B2(n_98),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_86),
.C(n_32),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_122),
.A2(n_27),
.B1(n_24),
.B2(n_76),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_5),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_122),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_32),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_78),
.B1(n_27),
.B2(n_24),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_129),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_175),
.A2(n_124),
.B1(n_137),
.B2(n_121),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_125),
.A2(n_24),
.B1(n_86),
.B2(n_2),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_116),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_134),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_145),
.B(n_132),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_184),
.A2(n_187),
.B(n_189),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_116),
.B(n_144),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_196),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_136),
.B(n_134),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_120),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_212),
.C(n_10),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_120),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_197),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_121),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_124),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_206),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_142),
.B1(n_137),
.B2(n_143),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_205),
.B1(n_178),
.B2(n_203),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_181),
.A2(n_129),
.B(n_127),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_201),
.A2(n_203),
.B(n_208),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_137),
.B1(n_142),
.B2(n_127),
.Y(n_202)
);

OAI22x1_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_209),
.B1(n_179),
.B2(n_174),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_150),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_3),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_7),
.B(n_8),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_163),
.A2(n_4),
.B(n_5),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_153),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_7),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_154),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_11),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_217),
.B(n_236),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_223),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_224),
.B1(n_214),
.B2(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_199),
.B1(n_195),
.B2(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_203),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_194),
.A2(n_182),
.B1(n_161),
.B2(n_172),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_226),
.B1(n_240),
.B2(n_185),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_182),
.B1(n_174),
.B2(n_171),
.Y(n_226)
);

NAND2xp33_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_182),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_226),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_182),
.B(n_170),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_234),
.B(n_207),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_173),
.B(n_8),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_206),
.B(n_198),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_241),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_8),
.B(n_10),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_204),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_191),
.Y(n_244)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_242),
.A2(n_257),
.B(n_260),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_261),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_188),
.C(n_196),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_215),
.C(n_212),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_204),
.B(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_220),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_258),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_255),
.B1(n_256),
.B2(n_224),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_238),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_198),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_221),
.A2(n_197),
.B1(n_185),
.B2(n_205),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_259),
.A2(n_258),
.B1(n_219),
.B2(n_229),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_267),
.A2(n_270),
.B1(n_275),
.B2(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_269),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_259),
.A2(n_229),
.B1(n_232),
.B2(n_223),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_243),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_235),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_273),
.A2(n_278),
.B(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_277),
.C(n_280),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_255),
.A2(n_240),
.B1(n_227),
.B2(n_222),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_261),
.C(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_235),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_250),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_222),
.C(n_228),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_257),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_286),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_228),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_249),
.C(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_289),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_242),
.B1(n_234),
.B2(n_260),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_252),
.C(n_248),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_242),
.C(n_231),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_237),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_272),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_269),
.B1(n_270),
.B2(n_265),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_290),
.B1(n_289),
.B2(n_287),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_R g299 ( 
.A(n_288),
.B(n_271),
.C(n_279),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_299),
.A2(n_233),
.B(n_285),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_305),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_267),
.B1(n_275),
.B2(n_265),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_301),
.A2(n_302),
.B1(n_292),
.B2(n_216),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_218),
.B1(n_268),
.B2(n_266),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_282),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_266),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_308),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_311),
.B(n_312),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_216),
.B1(n_291),
.B2(n_286),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_310),
.A2(n_304),
.B1(n_298),
.B2(n_297),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_285),
.C(n_237),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_300),
.B(n_305),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_313),
.A2(n_298),
.B(n_296),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_317),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_312),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_321),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_309),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_313),
.B(n_307),
.C(n_314),
.D(n_321),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_314),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_323),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_297),
.B(n_13),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_12),
.B(n_14),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_12),
.B(n_14),
.Y(n_329)
);


endmodule