module fake_jpeg_31102_n_46 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_21),
.B(n_0),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_26),
.C(n_0),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_18),
.B1(n_20),
.B2(n_11),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_22),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_36),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_32),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_40),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_5),
.C(n_8),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_39),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OAI311xp33_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_41),
.A3(n_13),
.B1(n_14),
.C1(n_15),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_12),
.C(n_16),
.Y(n_46)
);


endmodule