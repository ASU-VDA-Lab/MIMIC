module fake_jpeg_23224_n_249 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_5),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_15),
.Y(n_46)
);

CKINVDCx12_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_24),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_20),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_30),
.A2(n_14),
.B1(n_24),
.B2(n_25),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_25),
.B1(n_23),
.B2(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_30),
.B1(n_14),
.B2(n_24),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_73),
.B1(n_59),
.B2(n_21),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_64),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_22),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_50),
.B1(n_45),
.B2(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_25),
.B1(n_23),
.B2(n_16),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_90),
.B(n_93),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_34),
.C(n_39),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_82),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_85),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_45),
.B1(n_48),
.B2(n_52),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_58),
.B1(n_62),
.B2(n_73),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_56),
.B1(n_35),
.B2(n_21),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_46),
.B1(n_19),
.B2(n_21),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_84),
.B1(n_57),
.B2(n_61),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_39),
.C(n_38),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_35),
.B1(n_33),
.B2(n_39),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_92),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_96),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_103),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_60),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_87),
.B(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_74),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_41),
.B1(n_44),
.B2(n_33),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_109),
.B1(n_88),
.B2(n_83),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_61),
.B1(n_57),
.B2(n_55),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_121),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_76),
.C(n_93),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_129),
.C(n_95),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_120),
.B(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_122),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_91),
.B(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_132),
.B1(n_107),
.B2(n_96),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_74),
.Y(n_126)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_93),
.C(n_83),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_44),
.B1(n_41),
.B2(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_121),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_146),
.B(n_59),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_148),
.B(n_94),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_150),
.Y(n_155)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_105),
.B(n_99),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_108),
.B1(n_107),
.B2(n_105),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_124),
.B1(n_59),
.B2(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_109),
.B1(n_103),
.B2(n_113),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_122),
.B1(n_127),
.B2(n_131),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_116),
.C(n_129),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_139),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_116),
.B(n_129),
.C(n_126),
.D(n_121),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_162),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_125),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_170),
.A2(n_115),
.B1(n_104),
.B2(n_69),
.Y(n_190)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_69),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_173),
.B1(n_135),
.B2(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_172),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_174),
.A2(n_153),
.B1(n_140),
.B2(n_147),
.Y(n_180)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_177),
.B(n_174),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_183),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_144),
.B1(n_152),
.B2(n_143),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_191),
.B1(n_156),
.B2(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_188),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_115),
.B1(n_128),
.B2(n_104),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_190),
.B1(n_155),
.B2(n_166),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_115),
.B1(n_70),
.B2(n_44),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_160),
.C(n_157),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_202),
.C(n_203),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_197),
.B(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_155),
.B(n_163),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_170),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_200),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_201),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_180),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_172),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_161),
.C(n_41),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_51),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_51),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_207),
.A2(n_212),
.B(n_217),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_178),
.B1(n_189),
.B2(n_182),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_209),
.A2(n_201),
.B1(n_202),
.B2(n_199),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_182),
.B(n_41),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_7),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_5),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_0),
.C(n_1),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_216),
.C(n_208),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_0),
.C(n_1),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_7),
.B(n_12),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_223),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_5),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_224),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_19),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_215),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_8),
.Y(n_223)
);

AOI21x1_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_0),
.B(n_1),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_226),
.B(n_11),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_8),
.B(n_12),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_4),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_227),
.B(n_216),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_231),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_4),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_235),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_19),
.A3(n_4),
.B1(n_9),
.B2(n_11),
.C1(n_1),
.C2(n_2),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_224),
.B(n_225),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_218),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_240),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_0),
.B(n_2),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_2),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_243),
.B(n_237),
.Y(n_245)
);

AOI31xp33_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_246),
.A3(n_236),
.B(n_244),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_237),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_233),
.B(n_3),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_3),
.Y(n_249)
);


endmodule