module fake_jpeg_14704_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_53),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_22),
.B1(n_18),
.B2(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_42),
.B1(n_31),
.B2(n_28),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_57),
.Y(n_82)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_42),
.B1(n_46),
.B2(n_22),
.Y(n_73)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_41),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_45),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_76),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_72),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_31),
.B1(n_28),
.B2(n_24),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_28),
.B(n_31),
.Y(n_103)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_46),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_93),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_92),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_89),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_36),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_44),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_44),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_52),
.C(n_49),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_105),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_64),
.B1(n_65),
.B2(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_106),
.B1(n_123),
.B2(n_90),
.Y(n_141)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_112),
.B(n_116),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_49),
.C(n_41),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_115),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_58),
.B1(n_38),
.B2(n_66),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_88),
.B1(n_89),
.B2(n_116),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_53),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_102),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_86),
.B(n_73),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_19),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_58),
.B1(n_38),
.B2(n_48),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_116),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_141),
.B1(n_117),
.B2(n_108),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_129),
.A2(n_135),
.B1(n_25),
.B2(n_20),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_72),
.B1(n_92),
.B2(n_83),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_131),
.A2(n_143),
.B1(n_144),
.B2(n_138),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_88),
.B1(n_77),
.B2(n_87),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_82),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_116),
.A2(n_76),
.B1(n_24),
.B2(n_80),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_150),
.B(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_90),
.B1(n_80),
.B2(n_82),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_119),
.B1(n_111),
.B2(n_96),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_66),
.B1(n_50),
.B2(n_45),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_50),
.B1(n_45),
.B2(n_44),
.Y(n_144)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_151),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_146),
.B(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_44),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_69),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_99),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_114),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_156),
.B(n_164),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_112),
.B(n_103),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_96),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_105),
.B1(n_119),
.B2(n_106),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_173),
.B1(n_174),
.B2(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_181),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_136),
.B1(n_140),
.B2(n_145),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_127),
.A2(n_97),
.B1(n_107),
.B2(n_44),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_107),
.B1(n_97),
.B2(n_45),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_121),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_132),
.B(n_30),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_133),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_129),
.B1(n_139),
.B2(n_147),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_95),
.B(n_101),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_182),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_29),
.B(n_26),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_131),
.B(n_30),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_145),
.B1(n_172),
.B2(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_208),
.B1(n_209),
.B2(n_174),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_163),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_196),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_128),
.Y(n_200)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_207),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_158),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_210),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_144),
.B1(n_140),
.B2(n_143),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_25),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_25),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_213),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_155),
.B(n_101),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_157),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_184),
.A2(n_211),
.B1(n_197),
.B2(n_201),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_217),
.A2(n_225),
.B1(n_226),
.B2(n_230),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_164),
.C(n_182),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_154),
.C(n_166),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_185),
.C(n_194),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_227),
.C(n_228),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_188),
.B1(n_190),
.B2(n_210),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_161),
.B1(n_160),
.B2(n_156),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_180),
.B1(n_173),
.B2(n_181),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_101),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_95),
.C(n_69),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_35),
.B1(n_26),
.B2(n_29),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_193),
.A2(n_35),
.B1(n_29),
.B2(n_95),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_235),
.B1(n_237),
.B2(n_188),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_17),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_238),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_193),
.A2(n_25),
.B1(n_32),
.B2(n_23),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_186),
.A2(n_34),
.B1(n_32),
.B2(n_23),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_17),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_17),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_34),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_207),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_189),
.B(n_186),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_226),
.B(n_231),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_242),
.A2(n_251),
.B1(n_253),
.B2(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_190),
.B(n_196),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_1),
.B(n_2),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_236),
.B(n_206),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_252),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_203),
.B1(n_195),
.B2(n_205),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_206),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_203),
.B1(n_205),
.B2(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_258),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_204),
.B1(n_191),
.B2(n_208),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_34),
.Y(n_274)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_238),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_10),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_265),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_216),
.C(n_219),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_245),
.C(n_259),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_220),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_241),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_255),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_239),
.C(n_235),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_274),
.Y(n_279)
);

AO21x1_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_278),
.B(n_11),
.Y(n_291)
);

OAI321xp33_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_34),
.A3(n_32),
.B1(n_23),
.B2(n_5),
.C(n_6),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_286),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_276),
.A2(n_251),
.B1(n_242),
.B2(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_282),
.B(n_283),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_240),
.B1(n_256),
.B2(n_253),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_268),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_292),
.C(n_267),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_245),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_287),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_11),
.B(n_16),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_291),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_32),
.C(n_23),
.Y(n_292)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_266),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_306),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_302),
.C(n_305),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_272),
.B1(n_274),
.B2(n_4),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_7),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_2),
.C(n_3),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_3),
.C(n_4),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_3),
.C(n_6),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_283),
.B1(n_282),
.B2(n_279),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_291),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_279),
.B(n_8),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_314),
.B(n_316),
.Y(n_321)
);

NAND2x1_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_7),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_10),
.B(n_12),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_10),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_319),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_308),
.B(n_305),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_322),
.B(n_13),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_299),
.B(n_306),
.Y(n_322)
);

A2O1A1O1Ixp25_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_315),
.B(n_310),
.C(n_307),
.D(n_313),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_326),
.B(n_13),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_309),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_321),
.C(n_14),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_329),
.C(n_327),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_15),
.B(n_16),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_16),
.Y(n_333)
);


endmodule