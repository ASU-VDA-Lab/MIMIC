module real_aes_6733_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g172 ( .A1(n_0), .A2(n_173), .B(n_176), .C(n_180), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_1), .B(n_164), .Y(n_183) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_2), .B(n_88), .C(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g119 ( .A(n_2), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_3), .B(n_174), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_4), .A2(n_133), .B(n_486), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_5), .A2(n_138), .B(n_141), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_6), .A2(n_133), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_7), .B(n_164), .Y(n_492) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_8), .A2(n_166), .B(n_241), .Y(n_240) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_10), .A2(n_138), .B(n_141), .C(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g526 ( .A(n_11), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_12), .B(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_12), .B(n_41), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_13), .B(n_179), .Y(n_515) );
INVx1_ASAP7_75t_L g159 ( .A(n_14), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_15), .B(n_174), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_16), .A2(n_175), .B(n_546), .C(n_548), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_17), .B(n_164), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_18), .B(n_153), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_19), .A2(n_141), .B(n_144), .C(n_152), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_20), .A2(n_178), .B(n_234), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_21), .B(n_179), .Y(n_464) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_22), .A2(n_23), .B1(n_443), .B2(n_710), .C1(n_715), .C2(n_716), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_22), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_24), .B(n_179), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_25), .Y(n_460) );
INVx1_ASAP7_75t_L g499 ( .A(n_26), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_27), .A2(n_141), .B(n_152), .C(n_244), .Y(n_243) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_28), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_29), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_30), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g477 ( .A(n_31), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_32), .A2(n_133), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g136 ( .A(n_33), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_34), .A2(n_192), .B(n_193), .C(n_197), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_35), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_36), .A2(n_178), .B(n_489), .C(n_491), .Y(n_488) );
INVxp67_ASAP7_75t_L g478 ( .A(n_37), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_38), .B(n_246), .Y(n_245) );
CKINVDCx14_ASAP7_75t_R g487 ( .A(n_39), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_40), .A2(n_141), .B(n_152), .C(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g103 ( .A(n_41), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_42), .A2(n_180), .B(n_524), .C(n_525), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_43), .B(n_132), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_44), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_45), .B(n_174), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_46), .B(n_133), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_47), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_48), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_49), .A2(n_192), .B(n_197), .C(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g177 ( .A(n_50), .Y(n_177) );
INVx1_ASAP7_75t_L g220 ( .A(n_51), .Y(n_220) );
INVx1_ASAP7_75t_L g532 ( .A(n_52), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_53), .B(n_133), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_54), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_55), .A2(n_100), .B1(n_108), .B2(n_721), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g522 ( .A(n_56), .Y(n_522) );
INVx1_ASAP7_75t_L g139 ( .A(n_57), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_58), .B(n_133), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_59), .B(n_164), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_60), .A2(n_151), .B(n_207), .C(n_209), .Y(n_206) );
INVx1_ASAP7_75t_L g158 ( .A(n_61), .Y(n_158) );
INVx1_ASAP7_75t_SL g490 ( .A(n_62), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_63), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_64), .B(n_174), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_65), .B(n_164), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_66), .B(n_175), .Y(n_231) );
INVx1_ASAP7_75t_L g463 ( .A(n_67), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_68), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_69), .B(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_70), .A2(n_141), .B(n_197), .C(n_260), .Y(n_259) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_71), .Y(n_205) );
INVx1_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_73), .A2(n_133), .B(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_74), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_75), .A2(n_133), .B(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_76), .A2(n_122), .B1(n_123), .B2(n_437), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_76), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_77), .A2(n_132), .B(n_473), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_78), .Y(n_496) );
INVx1_ASAP7_75t_L g544 ( .A(n_79), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_80), .B(n_149), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_81), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_82), .A2(n_133), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g547 ( .A(n_83), .Y(n_547) );
INVx2_ASAP7_75t_L g156 ( .A(n_84), .Y(n_156) );
INVx1_ASAP7_75t_L g514 ( .A(n_85), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_86), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_87), .B(n_179), .Y(n_232) );
OR2x2_ASAP7_75t_L g116 ( .A(n_88), .B(n_117), .Y(n_116) );
OR2x2_ASAP7_75t_L g446 ( .A(n_88), .B(n_118), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_88), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_89), .A2(n_141), .B(n_197), .C(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_90), .B(n_133), .Y(n_190) );
INVx1_ASAP7_75t_L g194 ( .A(n_91), .Y(n_194) );
INVxp67_ASAP7_75t_L g210 ( .A(n_92), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_93), .B(n_166), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_94), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g227 ( .A(n_95), .Y(n_227) );
INVx1_ASAP7_75t_L g261 ( .A(n_96), .Y(n_261) );
INVx2_ASAP7_75t_L g535 ( .A(n_97), .Y(n_535) );
AND2x2_ASAP7_75t_L g222 ( .A(n_98), .B(n_155), .Y(n_222) );
INVx1_ASAP7_75t_SL g721 ( .A(n_100), .Y(n_721) );
CKINVDCx6p67_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OA21x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_114), .B(n_441), .Y(n_108) );
BUFx2_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_SL g720 ( .A(n_112), .Y(n_720) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_121), .B(n_438), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_116), .Y(n_440) );
NOR2x2_ASAP7_75t_L g718 ( .A(n_117), .B(n_448), .Y(n_718) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g447 ( .A(n_118), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_123), .A2(n_444), .B1(n_447), .B2(n_449), .Y(n_443) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g710 ( .A1(n_124), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_710) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_373), .Y(n_124) );
NOR5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_304), .C(n_333), .D(n_353), .E(n_360), .Y(n_125) );
OAI211xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_184), .B(n_248), .C(n_291), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_128), .A2(n_376), .B1(n_378), .B2(n_379), .Y(n_375) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_129), .Y(n_251) );
AND2x4_ASAP7_75t_L g284 ( .A(n_129), .B(n_285), .Y(n_284) );
INVx5_ASAP7_75t_L g302 ( .A(n_129), .Y(n_302) );
AND2x2_ASAP7_75t_L g311 ( .A(n_129), .B(n_303), .Y(n_311) );
AND2x2_ASAP7_75t_L g323 ( .A(n_129), .B(n_188), .Y(n_323) );
AND2x2_ASAP7_75t_L g419 ( .A(n_129), .B(n_287), .Y(n_419) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_160), .Y(n_129) );
AOI21xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_140), .B(n_153), .Y(n_130) );
BUFx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_134), .B(n_138), .Y(n_228) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g151 ( .A(n_135), .Y(n_151) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g235 ( .A(n_136), .Y(n_235) );
INVx1_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_137), .Y(n_147) );
INVx3_ASAP7_75t_L g175 ( .A(n_137), .Y(n_175) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
INVx1_ASAP7_75t_L g246 ( .A(n_137), .Y(n_246) );
BUFx3_ASAP7_75t_L g152 ( .A(n_138), .Y(n_152) );
INVx4_ASAP7_75t_SL g182 ( .A(n_138), .Y(n_182) );
INVx5_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_142), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B(n_150), .Y(n_144) );
INVx2_ASAP7_75t_L g149 ( .A(n_146), .Y(n_149) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_149), .A2(n_194), .B(n_195), .C(n_196), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_149), .A2(n_196), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_149), .A2(n_463), .B(n_464), .C(n_465), .Y(n_462) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_149), .A2(n_465), .B(n_514), .C(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_150), .A2(n_174), .B(n_499), .C(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_151), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_154), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g162 ( .A(n_155), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_155), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_155), .A2(n_217), .B(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_155), .A2(n_228), .B(n_496), .C(n_497), .Y(n_495) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_155), .A2(n_520), .B(n_527), .Y(n_519) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_156), .B(n_157), .Y(n_155) );
AND2x2_ASAP7_75t_L g167 ( .A(n_156), .B(n_157), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_162), .A2(n_510), .B(n_516), .Y(n_509) );
INVx2_ASAP7_75t_L g285 ( .A(n_163), .Y(n_285) );
AND2x2_ASAP7_75t_L g303 ( .A(n_163), .B(n_257), .Y(n_303) );
AND2x2_ASAP7_75t_L g322 ( .A(n_163), .B(n_256), .Y(n_322) );
AND2x2_ASAP7_75t_L g362 ( .A(n_163), .B(n_302), .Y(n_362) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_168), .B(n_183), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_165), .B(n_199), .Y(n_198) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_165), .A2(n_226), .B(n_236), .Y(n_225) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_165), .A2(n_258), .B(n_266), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_165), .B(n_267), .Y(n_266) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_165), .A2(n_459), .B(n_466), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_165), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_165), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_166), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_166), .A2(n_242), .B(n_243), .Y(n_241) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g238 ( .A(n_167), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g169 ( .A1(n_170), .A2(n_171), .B(n_172), .C(n_182), .Y(n_169) );
INVx2_ASAP7_75t_L g192 ( .A(n_171), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_171), .A2(n_182), .B(n_205), .C(n_206), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_SL g473 ( .A1(n_171), .A2(n_182), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_171), .A2(n_182), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_171), .A2(n_182), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_171), .A2(n_182), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g543 ( .A1(n_171), .A2(n_182), .B(n_544), .C(n_545), .Y(n_543) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_174), .B(n_210), .Y(n_209) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_174), .A2(n_208), .B1(n_477), .B2(n_478), .Y(n_476) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_175), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_178), .B(n_490), .Y(n_489) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g524 ( .A(n_179), .Y(n_524) );
INVx2_ASAP7_75t_L g465 ( .A(n_180), .Y(n_465) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_181), .Y(n_196) );
INVx1_ASAP7_75t_L g548 ( .A(n_181), .Y(n_548) );
INVx1_ASAP7_75t_L g197 ( .A(n_182), .Y(n_197) );
INVxp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_212), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_187), .A2(n_223), .A3(n_276), .B1(n_284), .B2(n_338), .C1(n_422), .C2(n_425), .Y(n_421) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_200), .Y(n_187) );
INVx5_ASAP7_75t_L g253 ( .A(n_188), .Y(n_253) );
AND2x2_ASAP7_75t_L g270 ( .A(n_188), .B(n_255), .Y(n_270) );
BUFx2_ASAP7_75t_L g348 ( .A(n_188), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_188), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g425 ( .A(n_188), .B(n_332), .Y(n_425) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_198), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_200), .B(n_214), .Y(n_279) );
INVx1_ASAP7_75t_L g306 ( .A(n_200), .Y(n_306) );
AND2x2_ASAP7_75t_L g319 ( .A(n_200), .B(n_239), .Y(n_319) );
AND2x2_ASAP7_75t_L g420 ( .A(n_200), .B(n_338), .Y(n_420) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g274 ( .A(n_201), .B(n_214), .Y(n_274) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_201), .Y(n_282) );
OR2x2_ASAP7_75t_L g289 ( .A(n_201), .B(n_239), .Y(n_289) );
AND2x2_ASAP7_75t_L g299 ( .A(n_201), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_201), .B(n_225), .Y(n_328) );
INVxp67_ASAP7_75t_L g352 ( .A(n_201), .Y(n_352) );
AND2x2_ASAP7_75t_L g359 ( .A(n_201), .B(n_223), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_201), .B(n_239), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_201), .B(n_224), .Y(n_385) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_201) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_202), .A2(n_485), .B(n_492), .Y(n_484) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_202), .A2(n_530), .B(n_536), .Y(n_529) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_202), .A2(n_542), .B(n_549), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_207), .A2(n_261), .B(n_262), .C(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_208), .B(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_208), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_223), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_214), .B(n_240), .Y(n_329) );
OR2x2_ASAP7_75t_L g351 ( .A(n_214), .B(n_224), .Y(n_351) );
AND2x2_ASAP7_75t_L g364 ( .A(n_214), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_214), .B(n_319), .Y(n_370) );
OAI211xp5_ASAP7_75t_SL g374 ( .A1(n_214), .A2(n_375), .B(n_380), .C(n_389), .Y(n_374) );
AND2x2_ASAP7_75t_L g435 ( .A(n_214), .B(n_239), .Y(n_435) );
INVx5_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g288 ( .A(n_215), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_215), .B(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_215), .B(n_283), .Y(n_295) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_215), .Y(n_297) );
OR2x2_ASAP7_75t_L g308 ( .A(n_215), .B(n_224), .Y(n_308) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_215), .B(n_299), .Y(n_313) );
AND2x2_ASAP7_75t_L g338 ( .A(n_215), .B(n_224), .Y(n_338) );
AND2x2_ASAP7_75t_L g358 ( .A(n_215), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g396 ( .A(n_215), .B(n_223), .Y(n_396) );
OR2x2_ASAP7_75t_L g399 ( .A(n_215), .B(n_385), .Y(n_399) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_239), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_224), .A2(n_343), .B(n_346), .C(n_352), .Y(n_342) );
INVx5_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_225), .B(n_239), .Y(n_273) );
AND2x2_ASAP7_75t_L g277 ( .A(n_225), .B(n_240), .Y(n_277) );
OR2x2_ASAP7_75t_L g283 ( .A(n_225), .B(n_239), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_229), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_228), .A2(n_460), .B(n_461), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_228), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_233), .A2(n_245), .B(n_247), .Y(n_244) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g470 ( .A(n_238), .Y(n_470) );
INVx1_ASAP7_75t_SL g300 ( .A(n_239), .Y(n_300) );
OR2x2_ASAP7_75t_L g428 ( .A(n_239), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_268), .B(n_271), .C(n_280), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AOI31xp33_ASAP7_75t_L g353 ( .A1(n_250), .A2(n_354), .A3(n_356), .B(n_357), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_251), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_252), .B(n_284), .Y(n_290) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_253), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g310 ( .A(n_253), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g315 ( .A(n_253), .B(n_285), .Y(n_315) );
AND2x2_ASAP7_75t_L g325 ( .A(n_253), .B(n_284), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_253), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g345 ( .A(n_253), .B(n_302), .Y(n_345) );
AND2x2_ASAP7_75t_L g350 ( .A(n_253), .B(n_322), .Y(n_350) );
OR2x2_ASAP7_75t_L g369 ( .A(n_253), .B(n_255), .Y(n_369) );
OR2x2_ASAP7_75t_L g371 ( .A(n_253), .B(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_253), .Y(n_418) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g318 ( .A(n_255), .B(n_285), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_255), .B(n_302), .Y(n_341) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx2_ASAP7_75t_L g287 ( .A(n_257), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_265), .Y(n_258) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx3_ASAP7_75t_L g491 ( .A(n_264), .Y(n_491) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g378 ( .A(n_270), .B(n_302), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g380 ( .A1(n_270), .A2(n_284), .A3(n_322), .B1(n_381), .B2(n_382), .C1(n_383), .C2(n_386), .Y(n_380) );
INVx1_ASAP7_75t_L g388 ( .A(n_270), .Y(n_388) );
NAND2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
INVx1_ASAP7_75t_SL g382 ( .A(n_272), .Y(n_382) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
OR2x2_ASAP7_75t_L g334 ( .A(n_273), .B(n_279), .Y(n_334) );
INVx1_ASAP7_75t_L g365 ( .A(n_273), .Y(n_365) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI32xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .A3(n_286), .B1(n_288), .B2(n_290), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AOI21xp33_ASAP7_75t_SL g320 ( .A1(n_283), .A2(n_298), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g335 ( .A(n_284), .Y(n_335) );
AND2x4_ASAP7_75t_L g332 ( .A(n_285), .B(n_302), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_285), .B(n_368), .Y(n_367) );
AOI322xp5_ASAP7_75t_L g397 ( .A1(n_286), .A2(n_313), .A3(n_332), .B1(n_365), .B2(n_398), .C1(n_400), .C2(n_401), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_286), .A2(n_363), .B1(n_427), .B2(n_428), .C(n_430), .Y(n_426) );
AND2x2_ASAP7_75t_L g314 ( .A(n_287), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_SL g294 ( .A(n_289), .Y(n_294) );
OR2x2_ASAP7_75t_L g366 ( .A(n_289), .B(n_351), .Y(n_366) );
OAI31xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .A3(n_296), .B(n_301), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_292), .A2(n_325), .B1(n_326), .B2(n_330), .Y(n_324) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g337 ( .A(n_294), .B(n_338), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_296), .A2(n_337), .B1(n_390), .B2(n_393), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g379 ( .A(n_299), .B(n_348), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_299), .B(n_338), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_300), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g413 ( .A(n_300), .B(n_351), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_301), .A2(n_396), .B1(n_409), .B2(n_412), .Y(n_408) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g317 ( .A(n_302), .Y(n_317) );
AND2x2_ASAP7_75t_L g400 ( .A(n_302), .B(n_322), .Y(n_400) );
OR2x2_ASAP7_75t_L g402 ( .A(n_302), .B(n_369), .Y(n_402) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_302), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_303), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_303), .B(n_348), .Y(n_356) );
OAI211xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_309), .B(n_312), .C(n_324), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_316), .B2(n_319), .C(n_320), .Y(n_312) );
INVxp67_ASAP7_75t_L g424 ( .A(n_315), .Y(n_424) );
INVx1_ASAP7_75t_L g391 ( .A(n_316), .Y(n_391) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g355 ( .A(n_317), .B(n_322), .Y(n_355) );
INVx1_ASAP7_75t_L g372 ( .A(n_318), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_318), .B(n_345), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g387 ( .A(n_322), .Y(n_387) );
AND2x2_ASAP7_75t_L g393 ( .A(n_322), .B(n_348), .Y(n_393) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_SL g381 ( .A(n_329), .Y(n_381) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_332), .B(n_368), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B1(n_336), .B2(n_339), .C(n_342), .Y(n_333) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g429 ( .A(n_338), .Y(n_429) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g347 ( .A(n_341), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_345), .B(n_404), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B(n_351), .Y(n_346) );
OAI211xp5_ASAP7_75t_SL g394 ( .A1(n_349), .A2(n_395), .B(n_397), .C(n_403), .Y(n_394) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g406 ( .A(n_351), .Y(n_406) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI222xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B1(n_366), .B2(n_367), .C1(n_370), .C2(n_371), .Y(n_360) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g436 ( .A(n_367), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_368), .B(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_368), .A2(n_415), .B1(n_417), .B2(n_420), .Y(n_414) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NOR4xp25_ASAP7_75t_L g373 ( .A(n_374), .B(n_394), .C(n_407), .D(n_426), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_376), .B(n_406), .Y(n_416) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g383 ( .A(n_381), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_384), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_414), .C(n_421), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx2_ASAP7_75t_L g423 ( .A(n_419), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_433), .B(n_436), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_438), .B(n_442), .C(n_719), .Y(n_441) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g711 ( .A(n_445), .Y(n_711) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g714 ( .A(n_447), .Y(n_714) );
INVx2_ASAP7_75t_L g712 ( .A(n_449), .Y(n_712) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_644), .Y(n_449) );
NAND5xp2_ASAP7_75t_L g450 ( .A(n_451), .B(n_573), .C(n_603), .D(n_624), .E(n_630), .Y(n_450) );
AOI221xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_506), .B1(n_537), .B2(n_539), .C(n_550), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_503), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_481), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_SL g624 ( .A1(n_456), .A2(n_493), .B(n_625), .C(n_628), .Y(n_624) );
AND2x2_ASAP7_75t_L g694 ( .A(n_456), .B(n_494), .Y(n_694) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_468), .Y(n_456) );
AND2x2_ASAP7_75t_L g552 ( .A(n_457), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g556 ( .A(n_457), .B(n_553), .Y(n_556) );
OR2x2_ASAP7_75t_L g582 ( .A(n_457), .B(n_494), .Y(n_582) );
AND2x2_ASAP7_75t_L g584 ( .A(n_457), .B(n_484), .Y(n_584) );
AND2x2_ASAP7_75t_L g602 ( .A(n_457), .B(n_483), .Y(n_602) );
INVx1_ASAP7_75t_L g635 ( .A(n_457), .Y(n_635) );
INVx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g505 ( .A(n_458), .Y(n_505) );
AND2x2_ASAP7_75t_L g538 ( .A(n_458), .B(n_484), .Y(n_538) );
AND2x2_ASAP7_75t_L g691 ( .A(n_458), .B(n_494), .Y(n_691) );
AND2x2_ASAP7_75t_L g572 ( .A(n_468), .B(n_482), .Y(n_572) );
OR2x2_ASAP7_75t_L g576 ( .A(n_468), .B(n_494), .Y(n_576) );
AND2x2_ASAP7_75t_L g601 ( .A(n_468), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g648 ( .A(n_468), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_468), .B(n_610), .Y(n_696) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B(n_479), .Y(n_468) );
INVx1_ASAP7_75t_L g554 ( .A(n_469), .Y(n_554) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_472), .A2(n_480), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI322xp33_ASAP7_75t_L g697 ( .A1(n_481), .A2(n_633), .A3(n_656), .B1(n_677), .B2(n_698), .C1(n_700), .C2(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_482), .B(n_553), .Y(n_700) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
AND2x2_ASAP7_75t_L g504 ( .A(n_483), .B(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_L g569 ( .A(n_483), .B(n_494), .Y(n_569) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g610 ( .A(n_484), .B(n_494), .Y(n_610) );
AND2x2_ASAP7_75t_L g654 ( .A(n_484), .B(n_493), .Y(n_654) );
AND2x2_ASAP7_75t_L g537 ( .A(n_493), .B(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g555 ( .A(n_493), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_493), .B(n_584), .Y(n_708) );
INVx3_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g503 ( .A(n_494), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_494), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g622 ( .A(n_494), .B(n_553), .Y(n_622) );
AND2x2_ASAP7_75t_L g649 ( .A(n_494), .B(n_584), .Y(n_649) );
OR2x2_ASAP7_75t_L g705 ( .A(n_494), .B(n_556), .Y(n_705) );
OR2x6_ASAP7_75t_L g494 ( .A(n_495), .B(n_501), .Y(n_494) );
INVx1_ASAP7_75t_SL g591 ( .A(n_503), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_504), .B(n_622), .Y(n_623) );
AND2x2_ASAP7_75t_L g657 ( .A(n_504), .B(n_647), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_504), .B(n_580), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_504), .B(n_702), .Y(n_701) );
OAI31xp33_ASAP7_75t_L g675 ( .A1(n_506), .A2(n_537), .A3(n_676), .B(n_678), .Y(n_675) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_507), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g658 ( .A(n_507), .B(n_593), .Y(n_658) );
OR2x2_ASAP7_75t_L g665 ( .A(n_507), .B(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g677 ( .A(n_507), .B(n_566), .Y(n_677) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g611 ( .A(n_508), .B(n_612), .Y(n_611) );
BUFx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g539 ( .A(n_509), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g560 ( .A(n_509), .Y(n_560) );
AND2x2_ASAP7_75t_L g597 ( .A(n_509), .B(n_541), .Y(n_597) );
AND2x2_ASAP7_75t_L g596 ( .A(n_518), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_SL g666 ( .A(n_518), .Y(n_666) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_519), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g566 ( .A(n_519), .B(n_529), .Y(n_566) );
INVx2_ASAP7_75t_L g586 ( .A(n_519), .Y(n_586) );
AND2x2_ASAP7_75t_L g600 ( .A(n_519), .B(n_529), .Y(n_600) );
AND2x2_ASAP7_75t_L g607 ( .A(n_519), .B(n_563), .Y(n_607) );
BUFx3_ASAP7_75t_L g617 ( .A(n_519), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_519), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g562 ( .A(n_528), .Y(n_562) );
AND2x2_ASAP7_75t_L g570 ( .A(n_528), .B(n_560), .Y(n_570) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g540 ( .A(n_529), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_529), .Y(n_594) );
INVx2_ASAP7_75t_SL g577 ( .A(n_538), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_538), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_538), .B(n_647), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_539), .B(n_617), .Y(n_670) );
INVx1_ASAP7_75t_SL g704 ( .A(n_539), .Y(n_704) );
INVx1_ASAP7_75t_SL g612 ( .A(n_540), .Y(n_612) );
INVx1_ASAP7_75t_SL g563 ( .A(n_541), .Y(n_563) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_541), .Y(n_574) );
OR2x2_ASAP7_75t_L g585 ( .A(n_541), .B(n_560), .Y(n_585) );
AND2x2_ASAP7_75t_L g599 ( .A(n_541), .B(n_560), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_541), .B(n_589), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_555), .B(n_557), .C(n_568), .Y(n_550) );
AOI31xp33_ASAP7_75t_L g667 ( .A1(n_551), .A2(n_668), .A3(n_669), .B(n_670), .Y(n_667) );
AND2x2_ASAP7_75t_L g640 ( .A(n_552), .B(n_569), .Y(n_640) );
BUFx3_ASAP7_75t_L g580 ( .A(n_553), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_553), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g616 ( .A(n_553), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_553), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g571 ( .A(n_556), .Y(n_571) );
OAI222xp33_ASAP7_75t_L g680 ( .A1(n_556), .A2(n_681), .B1(n_684), .B2(n_685), .C1(n_686), .C2(n_687), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_564), .Y(n_557) );
INVx1_ASAP7_75t_L g686 ( .A(n_558), .Y(n_686) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_560), .B(n_563), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_560), .B(n_586), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_560), .B(n_561), .Y(n_656) );
INVx1_ASAP7_75t_L g707 ( .A(n_560), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_561), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g709 ( .A(n_561), .Y(n_709) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx2_ASAP7_75t_L g589 ( .A(n_562), .Y(n_589) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_563), .Y(n_632) );
AOI32xp33_ASAP7_75t_L g568 ( .A1(n_564), .A2(n_569), .A3(n_570), .B1(n_571), .B2(n_572), .Y(n_568) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_566), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g643 ( .A(n_566), .Y(n_643) );
OR2x2_ASAP7_75t_L g684 ( .A(n_566), .B(n_585), .Y(n_684) );
INVx1_ASAP7_75t_L g620 ( .A(n_567), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_569), .B(n_580), .Y(n_605) );
INVx3_ASAP7_75t_L g614 ( .A(n_569), .Y(n_614) );
AOI322xp5_ASAP7_75t_L g630 ( .A1(n_569), .A2(n_614), .A3(n_631), .B1(n_633), .B2(n_636), .C1(n_640), .C2(n_641), .Y(n_630) );
AND2x2_ASAP7_75t_L g606 ( .A(n_570), .B(n_607), .Y(n_606) );
INVxp67_ASAP7_75t_L g683 ( .A(n_570), .Y(n_683) );
A2O1A1O1Ixp25_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B(n_578), .C(n_586), .D(n_587), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_574), .B(n_617), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_576), .A2(n_588), .B1(n_591), .B2(n_592), .C(n_595), .Y(n_587) );
INVx1_ASAP7_75t_SL g702 ( .A(n_576), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .B(n_585), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_580), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI221xp5_ASAP7_75t_SL g672 ( .A1(n_582), .A2(n_666), .B1(n_673), .B2(n_674), .C(n_675), .Y(n_672) );
OAI222xp33_ASAP7_75t_L g703 ( .A1(n_583), .A2(n_704), .B1(n_705), .B2(n_706), .C1(n_708), .C2(n_709), .Y(n_703) );
AND2x2_ASAP7_75t_L g661 ( .A(n_584), .B(n_647), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_584), .A2(n_599), .B(n_646), .Y(n_673) );
INVx1_ASAP7_75t_L g687 ( .A(n_584), .Y(n_687) );
INVx2_ASAP7_75t_SL g590 ( .A(n_585), .Y(n_590) );
AND2x2_ASAP7_75t_L g593 ( .A(n_586), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_SL g627 ( .A(n_589), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_589), .B(n_599), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_590), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_590), .B(n_600), .Y(n_629) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_598), .B(n_601), .Y(n_595) );
INVx1_ASAP7_75t_SL g613 ( .A(n_597), .Y(n_613) );
AND2x2_ASAP7_75t_L g660 ( .A(n_597), .B(n_643), .Y(n_660) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g699 ( .A(n_599), .B(n_617), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_600), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g685 ( .A(n_601), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B1(n_608), .B2(n_615), .C(n_618), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_612), .A2(n_619), .B1(n_621), .B2(n_623), .Y(n_618) );
OR2x2_ASAP7_75t_L g689 ( .A(n_613), .B(n_617), .Y(n_689) );
OR2x2_ASAP7_75t_L g692 ( .A(n_613), .B(n_627), .Y(n_692) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_634), .A2(n_689), .B1(n_690), .B2(n_692), .C(n_693), .Y(n_688) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND3xp33_ASAP7_75t_SL g644 ( .A(n_645), .B(n_659), .C(n_671), .Y(n_644) );
AOI222xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_650), .B1(n_652), .B2(n_655), .C1(n_657), .C2(n_658), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_647), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g669 ( .A(n_649), .Y(n_669) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_664), .C(n_667), .Y(n_659) );
INVx1_ASAP7_75t_L g674 ( .A(n_660), .Y(n_674) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI21xp33_ASAP7_75t_L g693 ( .A1(n_664), .A2(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NOR5xp2_ASAP7_75t_L g671 ( .A(n_672), .B(n_680), .C(n_688), .D(n_697), .E(n_703), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
endmodule