module fake_jpeg_11469_n_179 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_1),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_36),
.B(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g84 ( 
.A(n_39),
.Y(n_84)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_2),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_12),
.B(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_49),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_22),
.A2(n_5),
.B(n_6),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_53),
.Y(n_87)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_22),
.B(n_6),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_8),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_82),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_10),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_9),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_71),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_35),
.A2(n_17),
.B1(n_15),
.B2(n_21),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_76),
.B1(n_79),
.B2(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_26),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_34),
.A2(n_15),
.B1(n_21),
.B2(n_17),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_74),
.B1(n_54),
.B2(n_53),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_17),
.B1(n_18),
.B2(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_38),
.A2(n_18),
.B1(n_32),
.B2(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_30),
.B(n_31),
.C(n_26),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_39),
.B(n_46),
.C(n_42),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_87),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_91),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_99),
.Y(n_115)
);

AO22x2_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_52),
.B1(n_43),
.B2(n_54),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_110),
.B1(n_114),
.B2(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_37),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_11),
.B1(n_46),
.B2(n_73),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_75),
.B(n_66),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_46),
.C(n_11),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_11),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_60),
.B(n_81),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_86),
.B1(n_72),
.B2(n_62),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_88),
.B(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_75),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_68),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_72),
.B1(n_62),
.B2(n_89),
.Y(n_114)
);

NOR4xp25_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_84),
.C(n_85),
.D(n_66),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_129),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_84),
.B(n_61),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_108),
.B(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_94),
.B1(n_99),
.B2(n_93),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_98),
.B1(n_94),
.B2(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_92),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_122),
.C(n_132),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_96),
.B(n_106),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_136),
.B(n_121),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_144),
.B1(n_122),
.B2(n_123),
.Y(n_150)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_140),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_94),
.B1(n_110),
.B2(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_117),
.B1(n_124),
.B2(n_120),
.Y(n_152)
);

OAI22x1_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_119),
.B1(n_133),
.B2(n_129),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_124),
.B1(n_128),
.B2(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_115),
.B1(n_123),
.B2(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_131),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_151),
.B(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_142),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_154),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_128),
.B(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_128),
.C(n_130),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_156),
.C(n_137),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_125),
.C(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_143),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_161),
.C(n_159),
.Y(n_167)
);

AO221x1_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_136),
.B1(n_146),
.B2(n_140),
.C(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_160),
.A2(n_156),
.B(n_150),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_157),
.B(n_161),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_172),
.B(n_134),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_158),
.C(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_157),
.C(n_139),
.Y(n_173)
);

OR2x6_ASAP7_75t_SL g172 ( 
.A(n_165),
.B(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_174),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_155),
.C(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_141),
.C(n_140),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_176),
.Y(n_179)
);


endmodule