module fake_netlist_5_1559_n_1167 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1167);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1167;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_843;
wire n_855;
wire n_389;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_1055;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_155;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_1157;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_443;
wire n_293;
wire n_372;
wire n_244;
wire n_677;
wire n_173;
wire n_859;
wire n_864;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_753;
wire n_621;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_212;
wire n_498;
wire n_516;
wire n_385;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_1024;
wire n_556;
wire n_1063;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_1163;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1100;
wire n_862;
wire n_900;
wire n_1016;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_731;
wire n_390;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_167;
wire n_607;
wire n_976;
wire n_1096;
wire n_234;
wire n_343;
wire n_1095;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_156;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_157;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_750;
wire n_669;
wire n_742;
wire n_995;
wire n_454;
wire n_961;
wire n_472;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_1149;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1073;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_1020;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_196;
wire n_211;
wire n_218;
wire n_400;
wire n_962;
wire n_181;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_1071;
wire n_485;
wire n_1043;
wire n_1165;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_974;
wire n_395;
wire n_164;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_432;
wire n_311;
wire n_813;
wire n_1159;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_685;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_928;
wire n_749;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_866;
wire n_573;
wire n_796;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_151;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_1031;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_834;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1000;
wire n_239;
wire n_466;
wire n_1164;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_170;
wire n_332;
wire n_1053;
wire n_1101;
wire n_161;
wire n_273;
wire n_1106;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_774;
wire n_365;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_176;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_832;
wire n_795;
wire n_695;
wire n_857;
wire n_180;
wire n_1072;
wire n_656;
wire n_560;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_160;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_154;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_200;
wire n_1056;
wire n_162;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_1029;
wire n_166;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_82),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_149),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_54),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_13),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_55),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_113),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_62),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_20),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_9),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_7),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_87),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_106),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_39),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_1),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_63),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_93),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_66),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_96),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_38),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_150),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_53),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_4),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_103),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_15),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_27),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_101),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_49),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_18),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_31),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_8),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_35),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_11),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_99),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_47),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_3),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_147),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_136),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_116),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_188),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_161),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_163),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_168),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_170),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_173),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_157),
.B(n_0),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_176),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_180),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_192),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_182),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_191),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_158),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_227),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

BUFx8_ASAP7_75t_SL g234 ( 
.A(n_221),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_202),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_221),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_205),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_218),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_226),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_174),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_229),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_210),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_212),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_217),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_216),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_220),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_222),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_223),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_225),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_221),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_203),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_227),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_227),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_214),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_239),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_230),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_242),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

INVxp33_ASAP7_75t_SL g296 ( 
.A(n_269),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

BUFx6f_ASAP7_75t_SL g299 ( 
.A(n_238),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_239),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_269),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_250),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_267),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_238),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_271),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_267),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_254),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_276),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_285),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_280),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_285),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_287),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_308),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_277),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_264),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_277),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_286),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_309),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_300),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_310),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_310),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_296),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_313),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_261),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_296),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_275),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_314),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_312),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_271),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_312),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_311),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_311),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_354),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_318),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_252),
.Y(n_358)
);

OAI21x1_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_315),
.B(n_307),
.Y(n_359)
);

BUFx8_ASAP7_75t_SL g360 ( 
.A(n_325),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_318),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_235),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_345),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_291),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_317),
.Y(n_366)
);

AOI22x1_ASAP7_75t_SL g367 ( 
.A1(n_325),
.A2(n_247),
.B1(n_255),
.B2(n_254),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_342),
.Y(n_370)
);

OAI21x1_ASAP7_75t_L g371 ( 
.A1(n_320),
.A2(n_329),
.B(n_326),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_321),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_259),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_261),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_305),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_355),
.A2(n_260),
.B1(n_231),
.B2(n_268),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_293),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_294),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

NAND3xp33_ASAP7_75t_L g394 ( 
.A(n_335),
.B(n_241),
.C(n_240),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_328),
.A2(n_297),
.B(n_295),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_331),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_332),
.B(n_155),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_334),
.B(n_305),
.Y(n_402)
);

CKINVDCx6p67_ASAP7_75t_R g403 ( 
.A(n_330),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_317),
.B(n_255),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_345),
.A2(n_256),
.B1(n_243),
.B2(n_253),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_339),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_343),
.B(n_263),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_343),
.B(n_263),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_345),
.A2(n_299),
.B1(n_305),
.B2(n_155),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_345),
.A2(n_299),
.B1(n_302),
.B2(n_274),
.Y(n_415)
);

OAI22x1_ASAP7_75t_L g416 ( 
.A1(n_317),
.A2(n_236),
.B1(n_234),
.B2(n_158),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_345),
.A2(n_299),
.B1(n_302),
.B2(n_292),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_339),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_347),
.B(n_247),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_347),
.B(n_159),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_317),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_367),
.B(n_234),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_418),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_360),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_375),
.B(n_292),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_360),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_424),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_366),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_424),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_368),
.B(n_378),
.Y(n_437)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_179),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_R g439 ( 
.A(n_373),
.B(n_152),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_425),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_403),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_379),
.B(n_162),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_392),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_392),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_392),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_357),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_392),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_393),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_393),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_376),
.B(n_189),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_393),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_421),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_393),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_410),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_411),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_377),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_377),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_376),
.B(n_187),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_414),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_377),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_359),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_420),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_368),
.B(n_151),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_372),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_371),
.B(n_188),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_377),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_383),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_369),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_435),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g479 ( 
.A(n_440),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_449),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_435),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_441),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_447),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_444),
.B(n_374),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_426),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_447),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_456),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_441),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_463),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_447),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_431),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

BUFx10_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_374),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_443),
.B(n_407),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_445),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_446),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_427),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_446),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_431),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_430),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_450),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_450),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_434),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_447),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_451),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_433),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_469),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_433),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_451),
.B(n_404),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_452),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_453),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_453),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_481),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_509),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_477),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_498),
.B(n_407),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_409),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_480),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_481),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_515),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_512),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_487),
.B(n_409),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_485),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_490),
.A2(n_400),
.B1(n_415),
.B2(n_388),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_483),
.A2(n_400),
.B1(n_405),
.B2(n_422),
.Y(n_532)
);

BUFx4f_ASAP7_75t_L g533 ( 
.A(n_509),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_514),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_509),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_485),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_479),
.B(n_396),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_488),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_486),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_506),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_495),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_499),
.B(n_402),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_496),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_507),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_508),
.B(n_437),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_517),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_484),
.B(n_398),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_500),
.B(n_402),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_495),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_483),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_504),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_496),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_504),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_486),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_486),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_489),
.B(n_443),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_489),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_496),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_502),
.B(n_381),
.Y(n_562)
);

BUFx8_ASAP7_75t_SL g563 ( 
.A(n_494),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_491),
.B(n_401),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_493),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_505),
.B(n_358),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_517),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_493),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_493),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_510),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_516),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_492),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_492),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_478),
.B(n_468),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_503),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_503),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_494),
.A2(n_401),
.B1(n_399),
.B2(n_397),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_513),
.B(n_455),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_513),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_511),
.B(n_382),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_511),
.B(n_468),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_509),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_508),
.B(n_464),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_498),
.B(n_381),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_498),
.B(n_397),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_481),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_517),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_509),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_514),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_481),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_477),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_498),
.B(n_395),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_498),
.B(n_358),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g595 ( 
.A(n_514),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_498),
.B(n_417),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_481),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_509),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_477),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_498),
.B(n_385),
.Y(n_600)
);

BUFx4f_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_585),
.B(n_397),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_546),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_561),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_521),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_524),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_527),
.Y(n_608)
);

INVx6_ASAP7_75t_L g609 ( 
.A(n_552),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_549),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_592),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_520),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_523),
.B(n_380),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_529),
.A2(n_399),
.B1(n_198),
.B2(n_195),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_520),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_522),
.B(n_594),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_538),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_599),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_561),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_600),
.B(n_572),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_561),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_542),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_572),
.B(n_457),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_558),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_558),
.B(n_473),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_545),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_528),
.Y(n_628)
);

AO22x2_ASAP7_75t_L g629 ( 
.A1(n_531),
.A2(n_473),
.B1(n_428),
.B2(n_460),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_519),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_532),
.B(n_399),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_544),
.B(n_467),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_573),
.B(n_395),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_573),
.B(n_395),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_552),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_564),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_518),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_584),
.B(n_399),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_518),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_581),
.B(n_575),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_581),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_526),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_580),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_563),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_581),
.B(n_387),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_526),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_530),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_593),
.B(n_459),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_530),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_519),
.Y(n_650)
);

INVx5_ASAP7_75t_L g651 ( 
.A(n_574),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_533),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_581),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_L g654 ( 
.A(n_554),
.B(n_467),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_536),
.Y(n_655)
);

BUFx10_ASAP7_75t_L g656 ( 
.A(n_579),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_570),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_536),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_541),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_540),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_584),
.B(n_471),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_583),
.B(n_447),
.Y(n_662)
);

CKINVDCx8_ASAP7_75t_R g663 ( 
.A(n_534),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_520),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_552),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_593),
.B(n_465),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_541),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_551),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_551),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_583),
.B(n_553),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_575),
.B(n_387),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_553),
.B(n_466),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_562),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_559),
.B(n_476),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_555),
.B(n_586),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_562),
.B(n_543),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_555),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_547),
.Y(n_678)
);

BUFx6f_ASAP7_75t_SL g679 ( 
.A(n_567),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_576),
.B(n_391),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_567),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_582),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_550),
.B(n_356),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_544),
.B(n_554),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_586),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_582),
.Y(n_686)
);

INVx4_ASAP7_75t_SL g687 ( 
.A(n_574),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_SL g688 ( 
.A(n_644),
.B(n_455),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_616),
.B(n_537),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_616),
.B(n_596),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_635),
.B(n_570),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_620),
.B(n_596),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_618),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_676),
.B(n_554),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_676),
.B(n_547),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_603),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_673),
.B(n_577),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_617),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_673),
.B(n_633),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_629),
.A2(n_631),
.B1(n_613),
.B2(n_661),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_634),
.B(n_574),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_610),
.B(n_570),
.Y(n_702)
);

OAI221xp5_ASAP7_75t_L g703 ( 
.A1(n_614),
.A2(n_438),
.B1(n_566),
.B2(n_428),
.C(n_590),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_638),
.B(n_661),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_617),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_605),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_610),
.B(n_571),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_678),
.B(n_574),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_643),
.B(n_571),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_643),
.B(n_571),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_640),
.B(n_576),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_606),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_609),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_614),
.B(n_578),
.C(n_413),
.Y(n_714)
);

NOR3xp33_ASAP7_75t_L g715 ( 
.A(n_645),
.B(n_454),
.C(n_578),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_678),
.B(n_574),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_624),
.B(n_548),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_608),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_660),
.B(n_574),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_611),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_622),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_665),
.B(n_458),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_660),
.B(n_588),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_670),
.B(n_624),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_651),
.A2(n_595),
.B(n_458),
.C(n_474),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_629),
.A2(n_198),
.B1(n_188),
.B2(n_595),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_670),
.B(n_588),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_626),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_628),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_602),
.B(n_641),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_629),
.B(n_380),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_641),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_648),
.B(n_591),
.Y(n_733)
);

NAND2x1_ASAP7_75t_L g734 ( 
.A(n_684),
.B(n_556),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_648),
.B(n_391),
.C(n_461),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_679),
.A2(n_680),
.B1(n_671),
.B2(n_681),
.Y(n_736)
);

NOR2x1p5_ASAP7_75t_L g737 ( 
.A(n_657),
.B(n_461),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_651),
.B(n_656),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_666),
.B(n_591),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_666),
.B(n_597),
.Y(n_740)
);

INVxp33_ASAP7_75t_L g741 ( 
.A(n_683),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_609),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_651),
.B(n_656),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_636),
.B(n_474),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_623),
.B(n_597),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_675),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_653),
.B(n_587),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_630),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_650),
.B(n_559),
.Y(n_749)
);

BUFx8_ASAP7_75t_L g750 ( 
.A(n_679),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_639),
.B(n_642),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_646),
.B(n_560),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_653),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_684),
.B(n_525),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_604),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_637),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_647),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_636),
.B(n_557),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_649),
.B(n_560),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_658),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_655),
.B(n_565),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_755),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_690),
.B(n_667),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_689),
.B(n_663),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_726),
.A2(n_625),
.B1(n_356),
.B2(n_416),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_706),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_711),
.B(n_604),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_718),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_712),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_691),
.B(n_604),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_720),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_750),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_755),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_721),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_729),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_695),
.B(n_668),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_726),
.A2(n_714),
.B(n_731),
.C(n_700),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_728),
.Y(n_778)
);

AO22x2_ASAP7_75t_L g779 ( 
.A1(n_753),
.A2(n_698),
.B1(n_705),
.B2(n_694),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_704),
.B(n_625),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_747),
.B(n_607),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_693),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_728),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_746),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_741),
.B(n_385),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_696),
.Y(n_786)
);

NAND2x1p5_ASAP7_75t_L g787 ( 
.A(n_738),
.B(n_651),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_746),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_704),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_751),
.Y(n_790)
);

AO22x2_ASAP7_75t_L g791 ( 
.A1(n_694),
.A2(n_687),
.B1(n_632),
.B2(n_615),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_692),
.B(n_625),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_732),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_732),
.B(n_687),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_756),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_757),
.Y(n_796)
);

AO22x2_ASAP7_75t_L g797 ( 
.A1(n_735),
.A2(n_687),
.B1(n_632),
.B2(n_615),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_760),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_724),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_748),
.B(n_607),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_730),
.B(n_625),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_730),
.B(n_659),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_717),
.B(n_607),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_752),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_738),
.B(n_654),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_723),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_749),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_702),
.B(n_707),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_703),
.B(n_563),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_759),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_755),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_761),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_750),
.Y(n_813)
);

AO22x2_ASAP7_75t_L g814 ( 
.A1(n_719),
.A2(n_627),
.B1(n_664),
.B2(n_612),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_699),
.B(n_619),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_733),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_739),
.Y(n_817)
);

INVxp33_ASAP7_75t_SL g818 ( 
.A(n_688),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_740),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_727),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_715),
.A2(n_736),
.B1(n_710),
.B2(n_709),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_745),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_744),
.B(n_619),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_708),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_716),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_734),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_754),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_715),
.B(n_439),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_754),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_758),
.B(n_669),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_755),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_758),
.B(n_677),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_713),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_743),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_697),
.B(n_685),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_701),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_743),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_742),
.Y(n_838)
);

AO22x2_ASAP7_75t_L g839 ( 
.A1(n_722),
.A2(n_627),
.B1(n_664),
.B2(n_612),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_737),
.B(n_619),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_826),
.B(n_621),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_784),
.Y(n_842)
);

INVx5_ASAP7_75t_L g843 ( 
.A(n_772),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_814),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_777),
.A2(n_725),
.B(n_654),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_814),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_769),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_762),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_769),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_797),
.B(n_805),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_827),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_828),
.A2(n_780),
.B1(n_808),
.B2(n_809),
.Y(n_852)
);

AND2x6_ASAP7_75t_L g853 ( 
.A(n_821),
.B(n_621),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_824),
.B(n_621),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_825),
.B(n_672),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_778),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_783),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_762),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_833),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_803),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_813),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_837),
.B(n_682),
.Y(n_862)
);

AO22x1_ASAP7_75t_L g863 ( 
.A1(n_818),
.A2(n_662),
.B1(n_442),
.B2(n_674),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_825),
.B(n_662),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_800),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_789),
.B(n_380),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_829),
.B(n_682),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_840),
.B(n_792),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_762),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_793),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_785),
.B(n_380),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_794),
.B(n_834),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_794),
.B(n_686),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_771),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_816),
.B(n_817),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_784),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_819),
.B(n_820),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_773),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_838),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_806),
.B(n_662),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_793),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_788),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_774),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_779),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_781),
.Y(n_885)
);

OR2x6_ASAP7_75t_L g886 ( 
.A(n_797),
.B(n_652),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_770),
.A2(n_672),
.B(n_568),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_766),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_807),
.B(n_662),
.Y(n_889)
);

BUFx8_ASAP7_75t_L g890 ( 
.A(n_840),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_765),
.A2(n_652),
.B1(n_533),
.B2(n_601),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_SL g892 ( 
.A(n_764),
.B(n_390),
.C(n_442),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_773),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_768),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_822),
.B(n_674),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_775),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_799),
.B(n_674),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_847),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_843),
.B(n_801),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_845),
.A2(n_791),
.B(n_839),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_863),
.A2(n_791),
.B(n_839),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_861),
.B(n_386),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_859),
.B(n_823),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_886),
.A2(n_805),
.B(n_779),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_886),
.A2(n_787),
.B(n_834),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_843),
.A2(n_852),
.B1(n_850),
.B2(n_891),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_892),
.A2(n_835),
.B(n_763),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_843),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_848),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_849),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_884),
.A2(n_832),
.B(n_830),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_850),
.A2(n_836),
.B1(n_799),
.B2(n_790),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_848),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_875),
.B(n_815),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_853),
.A2(n_776),
.B(n_804),
.Y(n_915)
);

BUFx8_ASAP7_75t_L g916 ( 
.A(n_853),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_868),
.A2(n_802),
.B(n_804),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_872),
.B(n_844),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_862),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_877),
.A2(n_810),
.B(n_812),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_872),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_862),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_846),
.A2(n_866),
.B(n_871),
.C(n_879),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_853),
.A2(n_800),
.B1(n_767),
.B2(n_810),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_870),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_864),
.A2(n_831),
.B1(n_773),
.B2(n_811),
.Y(n_926)
);

INVx3_ASAP7_75t_SL g927 ( 
.A(n_859),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_856),
.B(n_782),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_841),
.B(n_831),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_897),
.A2(n_786),
.B(n_795),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_895),
.A2(n_798),
.B(n_796),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_881),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_853),
.A2(n_422),
.B(n_384),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_L g934 ( 
.A(n_880),
.B(n_811),
.C(n_167),
.Y(n_934)
);

XOR2xp5_ASAP7_75t_L g935 ( 
.A(n_878),
.B(n_412),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_890),
.B(n_386),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_889),
.A2(n_183),
.B(n_165),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_848),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_854),
.A2(n_601),
.B(n_533),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_857),
.A2(n_601),
.B(n_811),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_855),
.A2(n_569),
.B(n_565),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_851),
.A2(n_686),
.B1(n_535),
.B2(n_598),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_890),
.B(n_386),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_882),
.A2(n_569),
.B(n_535),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_883),
.B(n_674),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_887),
.A2(n_539),
.B(n_535),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_865),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_882),
.A2(n_598),
.B(n_525),
.Y(n_948)
);

BUFx4f_ASAP7_75t_L g949 ( 
.A(n_858),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_894),
.A2(n_190),
.B(n_184),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_L g951 ( 
.A(n_842),
.B(n_686),
.C(n_389),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_858),
.B(n_386),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_883),
.B(n_539),
.Y(n_953)
);

NOR2xp67_ASAP7_75t_L g954 ( 
.A(n_842),
.B(n_389),
.Y(n_954)
);

CKINVDCx10_ASAP7_75t_R g955 ( 
.A(n_858),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_869),
.B(n_389),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_865),
.A2(n_389),
.B(n_153),
.C(n_156),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_874),
.A2(n_598),
.B(n_525),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_841),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_869),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_908),
.B(n_873),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_916),
.B(n_906),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_916),
.B(n_873),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_907),
.B(n_860),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_915),
.B(n_869),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_911),
.B(n_885),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_900),
.B(n_893),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_927),
.B(n_867),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_901),
.B(n_888),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_917),
.B(n_876),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_918),
.B(n_896),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_920),
.B(n_0),
.Y(n_972)
);

NAND2xp33_ASAP7_75t_SL g973 ( 
.A(n_902),
.B(n_470),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_903),
.B(n_582),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_SL g975 ( 
.A(n_943),
.B(n_582),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_923),
.B(n_589),
.Y(n_976)
);

AND2x2_ASAP7_75t_SL g977 ( 
.A(n_936),
.B(n_362),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_SL g978 ( 
.A(n_924),
.B(n_589),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_962),
.A2(n_904),
.B(n_950),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_977),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_965),
.A2(n_967),
.B1(n_976),
.B2(n_978),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_972),
.A2(n_905),
.B(n_957),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_969),
.A2(n_912),
.B(n_899),
.C(n_937),
.Y(n_983)
);

AOI21xp33_ASAP7_75t_L g984 ( 
.A1(n_970),
.A2(n_934),
.B(n_951),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_963),
.B(n_955),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_964),
.B(n_932),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_966),
.A2(n_973),
.B(n_961),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_971),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_971),
.B(n_918),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_968),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_974),
.B(n_898),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_975),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_973),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_962),
.A2(n_952),
.B(n_956),
.C(n_933),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_972),
.A2(n_925),
.B1(n_949),
.B2(n_954),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_971),
.B(n_921),
.Y(n_996)
);

AO22x1_ASAP7_75t_L g997 ( 
.A1(n_972),
.A2(n_947),
.B1(n_960),
.B2(n_913),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_971),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_962),
.A2(n_930),
.B(n_931),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_SL g1000 ( 
.A1(n_972),
.A2(n_958),
.B(n_939),
.C(n_940),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_962),
.A2(n_948),
.B(n_944),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_962),
.A2(n_945),
.B(n_926),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_964),
.B(n_914),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_977),
.Y(n_1004)
);

O2A1O1Ixp5_ASAP7_75t_L g1005 ( 
.A1(n_997),
.A2(n_953),
.B(n_942),
.C(n_919),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_979),
.A2(n_935),
.B(n_941),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_983),
.A2(n_946),
.B(n_928),
.Y(n_1007)
);

OAI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_999),
.A2(n_959),
.B1(n_922),
.B2(n_913),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_985),
.B(n_913),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_993),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_990),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_982),
.B(n_910),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_1011),
.Y(n_1013)
);

NAND2x1p5_ASAP7_75t_L g1014 ( 
.A(n_1010),
.B(n_980),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1013),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_1013),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_1015),
.A2(n_1014),
.B(n_1005),
.Y(n_1017)
);

AOI22x1_ASAP7_75t_L g1018 ( 
.A1(n_1016),
.A2(n_987),
.B1(n_992),
.B2(n_1006),
.Y(n_1018)
);

BUFx5_ASAP7_75t_L g1019 ( 
.A(n_1018),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1017),
.B(n_1011),
.Y(n_1020)
);

BUFx8_ASAP7_75t_SL g1021 ( 
.A(n_1020),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_1019),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1022),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_SL g1024 ( 
.A1(n_1021),
.A2(n_1017),
.B1(n_1016),
.B2(n_1012),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1024),
.B(n_1016),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_1023),
.B(n_1009),
.C(n_1016),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1023),
.B(n_989),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1027),
.B(n_1026),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1025),
.Y(n_1029)
);

CKINVDCx11_ASAP7_75t_R g1030 ( 
.A(n_1026),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1029),
.Y(n_1031)
);

NOR2x1_ASAP7_75t_L g1032 ( 
.A(n_1028),
.B(n_1030),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1031),
.B(n_988),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1032),
.B(n_998),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1034),
.Y(n_1035)
);

AO21x2_ASAP7_75t_L g1036 ( 
.A1(n_1033),
.A2(n_1008),
.B(n_986),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1036),
.B(n_986),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_1035),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_L g1039 ( 
.A(n_1038),
.B(n_362),
.C(n_981),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1037),
.Y(n_1040)
);

NAND4xp75_ASAP7_75t_L g1041 ( 
.A(n_1040),
.B(n_1001),
.C(n_984),
.D(n_1007),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1039),
.B(n_995),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1042),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1041),
.B(n_996),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_1042),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_1044),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1045),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_1043),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1046),
.B(n_995),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1047),
.B(n_1003),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_1049),
.B(n_1048),
.Y(n_1051)
);

AO221x2_ASAP7_75t_L g1052 ( 
.A1(n_1050),
.A2(n_991),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1052),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1051),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_1054),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_1053),
.B(n_1),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1055),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1056),
.B(n_1004),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1057),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_1058),
.Y(n_1060)
);

AOI31xp33_ASAP7_75t_L g1061 ( 
.A1(n_1060),
.A2(n_153),
.A3(n_156),
.B(n_151),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1059),
.B(n_2),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1059),
.B(n_5),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1061),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1062),
.B(n_1002),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1063),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1066),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1065),
.B(n_980),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1068),
.B(n_1064),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1067),
.A2(n_160),
.B1(n_201),
.B2(n_196),
.Y(n_1070)
);

NOR2x1_ASAP7_75t_L g1071 ( 
.A(n_1069),
.B(n_160),
.Y(n_1071)
);

OAI32xp33_ASAP7_75t_L g1072 ( 
.A1(n_1070),
.A2(n_196),
.A3(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_1071),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1072),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1073),
.Y(n_1075)
);

OAI32xp33_ASAP7_75t_L g1076 ( 
.A1(n_1074),
.A2(n_199),
.A3(n_200),
.B1(n_984),
.B2(n_9),
.Y(n_1076)
);

NOR3x1_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_6),
.C(n_7),
.Y(n_1077)
);

NOR3x1_ASAP7_75t_L g1078 ( 
.A(n_1076),
.B(n_6),
.C(n_8),
.Y(n_1078)
);

NOR2x1p5_ASAP7_75t_L g1079 ( 
.A(n_1078),
.B(n_10),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1077),
.Y(n_1080)
);

AOI211xp5_ASAP7_75t_L g1081 ( 
.A1(n_1078),
.A2(n_185),
.B(n_12),
.C(n_13),
.Y(n_1081)
);

AO22x2_ASAP7_75t_L g1082 ( 
.A1(n_1080),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1079),
.A2(n_423),
.B1(n_464),
.B2(n_17),
.Y(n_1083)
);

NAND4xp25_ASAP7_75t_L g1084 ( 
.A(n_1081),
.B(n_14),
.C(n_16),
.D(n_17),
.Y(n_1084)
);

AOI211xp5_ASAP7_75t_L g1085 ( 
.A1(n_1084),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1082),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.C(n_22),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1085),
.B(n_1083),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1086),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_1088),
.B(n_1087),
.C(n_21),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_1088),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_1090),
.B(n_22),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1089),
.B(n_23),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1092),
.Y(n_1093)
);

NAND5xp2_ASAP7_75t_L g1094 ( 
.A(n_1091),
.B(n_23),
.C(n_24),
.D(n_25),
.E(n_26),
.Y(n_1094)
);

NAND2xp33_ASAP7_75t_SL g1095 ( 
.A(n_1093),
.B(n_24),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1094),
.B(n_25),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_1096),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_1095),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1096),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1097),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1098),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1101),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1100),
.Y(n_1104)
);

AO22x2_ASAP7_75t_L g1105 ( 
.A1(n_1103),
.A2(n_1102),
.B1(n_29),
.B2(n_30),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1104),
.B(n_28),
.Y(n_1106)
);

XNOR2xp5_ASAP7_75t_L g1107 ( 
.A(n_1105),
.B(n_30),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_1106),
.Y(n_1108)
);

OAI211xp5_ASAP7_75t_L g1109 ( 
.A1(n_1108),
.A2(n_994),
.B(n_33),
.C(n_34),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1107),
.A2(n_960),
.B1(n_938),
.B2(n_909),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1110),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1109),
.Y(n_1112)
);

OAI22x1_ASAP7_75t_L g1113 ( 
.A1(n_1111),
.A2(n_365),
.B1(n_36),
.B2(n_37),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_1112),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1114),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1113),
.B(n_32),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1114),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1115),
.A2(n_423),
.B1(n_960),
.B2(n_365),
.Y(n_1118)
);

AOI31xp33_ASAP7_75t_L g1119 ( 
.A1(n_1117),
.A2(n_40),
.A3(n_41),
.B(n_42),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1116),
.A2(n_423),
.B1(n_909),
.B2(n_938),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1120),
.A2(n_43),
.B(n_44),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_45),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1118),
.A2(n_423),
.B1(n_589),
.B2(n_472),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_423),
.B1(n_589),
.B2(n_432),
.Y(n_1124)
);

XOR2xp5_ASAP7_75t_L g1125 ( 
.A(n_1121),
.B(n_46),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_SL g1126 ( 
.A1(n_1123),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_1126)
);

NAND4xp25_ASAP7_75t_SL g1127 ( 
.A(n_1125),
.B(n_1124),
.C(n_1126),
.D(n_57),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1125),
.B(n_52),
.Y(n_1128)
);

XNOR2xp5_ASAP7_75t_L g1129 ( 
.A(n_1125),
.B(n_56),
.Y(n_1129)
);

XNOR2xp5_ASAP7_75t_L g1130 ( 
.A(n_1127),
.B(n_58),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1129),
.A2(n_1128),
.B1(n_432),
.B2(n_929),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1127),
.B(n_59),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1127),
.B(n_60),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_SL g1134 ( 
.A1(n_1127),
.A2(n_61),
.B(n_65),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1127),
.B(n_67),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1127),
.B(n_68),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1127),
.A2(n_69),
.B(n_70),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1127),
.B(n_71),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1127),
.B(n_72),
.Y(n_1139)
);

XOR2xp5_ASAP7_75t_L g1140 ( 
.A(n_1127),
.B(n_73),
.Y(n_1140)
);

AOI21xp33_ASAP7_75t_L g1141 ( 
.A1(n_1127),
.A2(n_74),
.B(n_75),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1127),
.B(n_76),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_SL g1143 ( 
.A1(n_1133),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_1143)
);

AOI222xp33_ASAP7_75t_L g1144 ( 
.A1(n_1130),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.C1(n_84),
.C2(n_85),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_R g1145 ( 
.A1(n_1140),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_1145)
);

XNOR2xp5_ASAP7_75t_L g1146 ( 
.A(n_1138),
.B(n_90),
.Y(n_1146)
);

AOI222xp33_ASAP7_75t_L g1147 ( 
.A1(n_1132),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.C1(n_95),
.C2(n_97),
.Y(n_1147)
);

OAI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_1135),
.A2(n_100),
.B1(n_102),
.B2(n_104),
.C(n_105),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1136),
.A2(n_108),
.B(n_109),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1139),
.A2(n_432),
.B1(n_929),
.B2(n_462),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1142),
.B(n_462),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1151),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1151),
.A2(n_1131),
.B1(n_1137),
.B2(n_1134),
.Y(n_1153)
);

NAND2xp33_ASAP7_75t_L g1154 ( 
.A(n_1146),
.B(n_1141),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1149),
.A2(n_1000),
.B(n_112),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1150),
.B(n_111),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_SL g1157 ( 
.A1(n_1153),
.A2(n_1145),
.B1(n_1148),
.B2(n_1143),
.Y(n_1157)
);

AOI322xp5_ASAP7_75t_L g1158 ( 
.A1(n_1154),
.A2(n_1144),
.A3(n_1147),
.B1(n_991),
.B2(n_118),
.C1(n_119),
.C2(n_120),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_SL g1159 ( 
.A1(n_1152),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1156),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1157),
.A2(n_1155),
.B1(n_125),
.B2(n_126),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1161),
.B(n_1158),
.Y(n_1162)
);

OAI221xp5_ASAP7_75t_R g1163 ( 
.A1(n_1162),
.A2(n_1160),
.B1(n_1159),
.B2(n_130),
.C(n_131),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1163),
.A2(n_124),
.B1(n_129),
.B2(n_132),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_SL g1165 ( 
.A1(n_1164),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_1165)
);

AOI211xp5_ASAP7_75t_L g1166 ( 
.A1(n_1165),
.A2(n_137),
.B(n_138),
.C(n_139),
.Y(n_1166)
);

AOI211xp5_ASAP7_75t_L g1167 ( 
.A1(n_1166),
.A2(n_140),
.B(n_141),
.C(n_142),
.Y(n_1167)
);


endmodule