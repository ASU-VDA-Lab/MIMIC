module real_jpeg_2047_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_249;
wire n_78;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_197;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_2),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_5),
.A2(n_19),
.B1(n_24),
.B2(n_34),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_5),
.A2(n_34),
.B1(n_64),
.B2(n_65),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_5),
.A2(n_34),
.B1(n_52),
.B2(n_54),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_19),
.B1(n_24),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_31),
.B1(n_52),
.B2(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_6),
.A2(n_31),
.B1(n_64),
.B2(n_65),
.Y(n_120)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_19),
.B1(n_24),
.B2(n_44),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_8),
.B(n_19),
.C(n_23),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_8),
.A2(n_44),
.B1(n_64),
.B2(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_8),
.A2(n_44),
.B1(n_52),
.B2(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_8),
.B(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_49),
.C(n_52),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_8),
.B(n_62),
.C(n_65),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_8),
.B(n_94),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_8),
.B(n_63),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_11),
.A2(n_14),
.B(n_262),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_11),
.B(n_263),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_36),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_35),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_32),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_32),
.Y(n_35)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B(n_30),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_18),
.A2(n_25),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

AO21x2_ASAP7_75t_SL g42 ( 
.A1(n_18),
.A2(n_25),
.B(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_18),
.A2(n_25),
.B1(n_33),
.B2(n_43),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_18),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_18)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_19),
.A2(n_24),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_19),
.B(n_148),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_28),
.B(n_89),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_32),
.B(n_38),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_72),
.B(n_261),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_70),
.C(n_71),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_39),
.A2(n_40),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.C(n_56),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_42),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

AOI211xp5_ASAP7_75t_SL g107 ( 
.A1(n_41),
.A2(n_103),
.B(n_108),
.C(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_41),
.B(n_83),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_41),
.A2(n_42),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_41),
.A2(n_42),
.B1(n_199),
.B2(n_204),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_41),
.A2(n_42),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_41),
.A2(n_204),
.B(n_215),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_41),
.A2(n_42),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_41),
.A2(n_42),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_42),
.B(n_84),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_42),
.B(n_57),
.C(n_237),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_42),
.B(n_246),
.C(n_250),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_45),
.A2(n_56),
.B1(n_57),
.B2(n_249),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_45),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_55),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_85),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_51),
.B(n_55),
.Y(n_70)
);

AO21x2_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_51),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_49),
.Y(n_50)
);

OA22x2_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_51),
.Y(n_165)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_52),
.B(n_159),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_56),
.A2(n_57),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_68),
.B(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_58),
.A2(n_68),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_63),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_59),
.A2(n_63),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_94),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_65),
.B(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_69),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_70),
.B(n_71),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_255),
.B(n_260),
.Y(n_72)
);

AOI21x1_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_229),
.B(n_252),
.Y(n_73)
);

OAI21x1_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_209),
.B(n_228),
.Y(n_74)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_189),
.B(n_208),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_136),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_122),
.B(n_135),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_SL g136 ( 
.A(n_78),
.B(n_137),
.C(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_110),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_110),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_97),
.C(n_106),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_96),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_82),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_81),
.A2(n_82),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_83),
.A2(n_84),
.B1(n_102),
.B2(n_103),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_83),
.A2(n_84),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_83),
.A2(n_103),
.B(n_109),
.C(n_180),
.Y(n_183)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_102),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_91),
.C(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_84),
.A2(n_221),
.B(n_224),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_84),
.B(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_90),
.A2(n_91),
.B1(n_133),
.B2(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_90),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_90),
.A2(n_91),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_90),
.B(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_90),
.A2(n_91),
.B1(n_146),
.B2(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_91),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_91),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_91),
.B(n_102),
.C(n_164),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_93),
.B(n_120),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_106),
.B1(n_107),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_103),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_103),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_141),
.C(n_145),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_102),
.A2(n_103),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_102),
.A2(n_103),
.B1(n_157),
.B2(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_102),
.A2(n_103),
.B1(n_145),
.B2(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_103),
.B(n_119),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_111),
.B(n_115),
.C(n_118),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_112),
.A2(n_113),
.B(n_116),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_112),
.A2(n_113),
.B(n_196),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_132),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_128),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_130),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_152),
.B(n_188),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_149),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_182),
.B(n_187),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_176),
.B(n_181),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_166),
.B(n_175),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_160),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_184),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_191),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_207),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_198),
.B1(n_205),
.B2(n_206),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_205),
.C(n_207),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_204),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_201),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_211),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_219),
.B2(n_220),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_219),
.C(n_225),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_224),
.A2(n_233),
.B1(n_234),
.B2(n_239),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_224),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_242),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_241),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_241),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_240),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_239),
.C(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_251),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_251),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_259),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);


endmodule