module real_aes_6537_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_0), .A2(n_168), .B(n_171), .C(n_175), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_1), .B(n_159), .Y(n_178) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_3), .B(n_169), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_4), .A2(n_132), .B(n_135), .C(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_5), .A2(n_127), .B(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_6), .A2(n_127), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_7), .B(n_159), .Y(n_530) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_8), .A2(n_161), .B(n_233), .Y(n_232) );
AND2x6_ASAP7_75t_L g132 ( .A(n_9), .B(n_133), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_10), .A2(n_132), .B(n_135), .C(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g490 ( .A(n_11), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_12), .B(n_39), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_13), .B(n_174), .Y(n_501) );
INVx1_ASAP7_75t_L g153 ( .A(n_14), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_15), .B(n_169), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_16), .A2(n_170), .B(n_510), .C(n_512), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_17), .B(n_159), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_18), .B(n_147), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_19), .A2(n_135), .B(n_138), .C(n_146), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_20), .A2(n_173), .B(n_241), .C(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_21), .B(n_174), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_22), .B(n_174), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_23), .Y(n_471) );
INVx1_ASAP7_75t_L g451 ( .A(n_24), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_25), .A2(n_135), .B(n_146), .C(n_236), .Y(n_235) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_26), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_27), .Y(n_497) );
INVx1_ASAP7_75t_L g465 ( .A(n_28), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_29), .A2(n_127), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g130 ( .A(n_30), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_31), .A2(n_185), .B(n_186), .C(n_190), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_32), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_33), .A2(n_744), .B1(n_749), .B2(n_750), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_33), .Y(n_749) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_34), .A2(n_173), .B(n_527), .C(n_529), .Y(n_526) );
INVxp67_ASAP7_75t_L g466 ( .A(n_35), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_36), .B(n_238), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_37), .A2(n_135), .B(n_146), .C(n_450), .Y(n_449) );
CKINVDCx14_ASAP7_75t_R g525 ( .A(n_38), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_40), .A2(n_175), .B(n_488), .C(n_489), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_41), .B(n_126), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_42), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_43), .B(n_169), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_44), .B(n_127), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_45), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_46), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_47), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_48), .A2(n_185), .B(n_190), .C(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g172 ( .A(n_49), .Y(n_172) );
INVx1_ASAP7_75t_L g216 ( .A(n_50), .Y(n_216) );
INVx1_ASAP7_75t_L g538 ( .A(n_51), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_52), .B(n_127), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_53), .Y(n_155) );
CKINVDCx14_ASAP7_75t_R g486 ( .A(n_54), .Y(n_486) );
INVx1_ASAP7_75t_L g133 ( .A(n_55), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_56), .B(n_127), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_57), .B(n_159), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_58), .A2(n_145), .B(n_201), .C(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g152 ( .A(n_59), .Y(n_152) );
INVx1_ASAP7_75t_SL g528 ( .A(n_60), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_61), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_62), .B(n_169), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_63), .B(n_159), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_64), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_65), .B(n_170), .Y(n_251) );
INVx1_ASAP7_75t_L g474 ( .A(n_66), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_67), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_68), .B(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_69), .A2(n_135), .B(n_190), .C(n_199), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g225 ( .A(n_70), .Y(n_225) );
INVx1_ASAP7_75t_L g764 ( .A(n_71), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_72), .A2(n_127), .B(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_73), .A2(n_95), .B1(n_747), .B2(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_73), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_74), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_75), .A2(n_127), .B(n_507), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_76), .A2(n_102), .B1(n_725), .B2(n_726), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_76), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_77), .A2(n_126), .B(n_461), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g448 ( .A(n_78), .Y(n_448) );
INVx1_ASAP7_75t_L g508 ( .A(n_79), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_80), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_80), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_81), .B(n_143), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_82), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_83), .A2(n_127), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g511 ( .A(n_84), .Y(n_511) );
INVx2_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
INVx1_ASAP7_75t_L g500 ( .A(n_86), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_87), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_88), .B(n_174), .Y(n_252) );
OR2x2_ASAP7_75t_L g110 ( .A(n_89), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g440 ( .A(n_89), .Y(n_440) );
OR2x2_ASAP7_75t_L g755 ( .A(n_89), .B(n_736), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_90), .A2(n_135), .B(n_190), .C(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_91), .B(n_127), .Y(n_183) );
INVx1_ASAP7_75t_L g187 ( .A(n_92), .Y(n_187) );
AOI22xp33_ASAP7_75t_SL g103 ( .A1(n_93), .A2(n_104), .B1(n_760), .B2(n_766), .Y(n_103) );
INVxp67_ASAP7_75t_L g228 ( .A(n_94), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_95), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_96), .B(n_161), .Y(n_491) );
INVx1_ASAP7_75t_L g200 ( .A(n_97), .Y(n_200) );
INVx1_ASAP7_75t_L g247 ( .A(n_98), .Y(n_247) );
INVx2_ASAP7_75t_L g541 ( .A(n_99), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_100), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g218 ( .A(n_101), .B(n_149), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_102), .Y(n_725) );
AO221x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_738), .B1(n_743), .B2(n_751), .C(n_756), .Y(n_104) );
OAI222xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_721), .B1(n_727), .B2(n_731), .C1(n_732), .C2(n_737), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OAI22xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_114), .B1(n_437), .B2(n_441), .Y(n_107) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_108), .A2(n_115), .B1(n_729), .B2(n_730), .Y(n_728) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g439 ( .A(n_111), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g736 ( .A(n_111), .Y(n_736) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_114), .A2(n_115), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_SL g115 ( .A(n_116), .B(n_392), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_327), .Y(n_116) );
NAND4xp25_ASAP7_75t_SL g117 ( .A(n_118), .B(n_272), .C(n_296), .D(n_319), .Y(n_117) );
AOI221xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_209), .B1(n_243), .B2(n_256), .C(n_259), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_179), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_121), .A2(n_157), .B1(n_210), .B2(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_121), .B(n_180), .Y(n_330) );
AND2x2_ASAP7_75t_L g349 ( .A(n_121), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_121), .B(n_333), .Y(n_419) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_157), .Y(n_121) );
AND2x2_ASAP7_75t_L g287 ( .A(n_122), .B(n_180), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_122), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g310 ( .A(n_122), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g315 ( .A(n_122), .B(n_158), .Y(n_315) );
INVx2_ASAP7_75t_L g347 ( .A(n_122), .Y(n_347) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_122), .Y(n_391) );
AND2x2_ASAP7_75t_L g408 ( .A(n_122), .B(n_285), .Y(n_408) );
INVx5_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g326 ( .A(n_123), .B(n_285), .Y(n_326) );
AND2x4_ASAP7_75t_L g340 ( .A(n_123), .B(n_157), .Y(n_340) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_123), .Y(n_344) );
AND2x2_ASAP7_75t_L g364 ( .A(n_123), .B(n_279), .Y(n_364) );
AND2x2_ASAP7_75t_L g414 ( .A(n_123), .B(n_181), .Y(n_414) );
AND2x2_ASAP7_75t_L g424 ( .A(n_123), .B(n_158), .Y(n_424) );
OR2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_154), .Y(n_123) );
AOI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_134), .B(n_147), .Y(n_124) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
NAND2x1p5_ASAP7_75t_L g248 ( .A(n_128), .B(n_132), .Y(n_248) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx1_ASAP7_75t_L g242 ( .A(n_130), .Y(n_242) );
INVx1_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_131), .Y(n_141) );
INVx3_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
INVx1_ASAP7_75t_L g238 ( .A(n_131), .Y(n_238) );
BUFx3_ASAP7_75t_L g146 ( .A(n_132), .Y(n_146) );
INVx4_ASAP7_75t_SL g177 ( .A(n_132), .Y(n_177) );
INVx5_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx3_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_136), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_142), .B(n_144), .Y(n_138) );
INVx2_ASAP7_75t_L g143 ( .A(n_140), .Y(n_143) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_143), .A2(n_187), .B(n_188), .C(n_189), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_143), .A2(n_189), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_143), .A2(n_474), .B(n_475), .C(n_476), .Y(n_473) );
O2A1O1Ixp5_ASAP7_75t_L g499 ( .A1(n_143), .A2(n_476), .B(n_500), .C(n_501), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_144), .A2(n_169), .B(n_451), .C(n_452), .Y(n_450) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_145), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_148), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_149), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_149), .A2(n_213), .B(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_149), .A2(n_248), .B(n_448), .C(n_449), .Y(n_447) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_149), .A2(n_484), .B(n_491), .Y(n_483) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_L g162 ( .A(n_150), .B(n_151), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_156), .A2(n_496), .B(n_502), .Y(n_495) );
AND2x2_ASAP7_75t_L g280 ( .A(n_157), .B(n_180), .Y(n_280) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_157), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_157), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g370 ( .A(n_157), .Y(n_370) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g258 ( .A(n_158), .B(n_195), .Y(n_258) );
AND2x2_ASAP7_75t_L g285 ( .A(n_158), .B(n_196), .Y(n_285) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_163), .B(n_178), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_160), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_160), .A2(n_197), .B(n_207), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_160), .B(n_208), .Y(n_207) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_160), .A2(n_246), .B(n_253), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_160), .B(n_454), .Y(n_453) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_160), .A2(n_470), .B(n_477), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_160), .B(n_503), .Y(n_502) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_161), .A2(n_234), .B(n_235), .Y(n_233) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g255 ( .A(n_162), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_177), .Y(n_164) );
INVx2_ASAP7_75t_L g185 ( .A(n_166), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_166), .A2(n_177), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_SL g461 ( .A1(n_166), .A2(n_177), .B(n_462), .C(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_166), .A2(n_177), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_166), .A2(n_177), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_166), .A2(n_177), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_SL g537 ( .A1(n_166), .A2(n_177), .B(n_538), .C(n_539), .Y(n_537) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_169), .B(n_228), .Y(n_227) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_169), .A2(n_202), .B1(n_465), .B2(n_466), .Y(n_464) );
INVx5_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_170), .B(n_490), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_173), .B(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g488 ( .A(n_174), .Y(n_488) );
INVx2_ASAP7_75t_L g476 ( .A(n_175), .Y(n_476) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_176), .Y(n_189) );
INVx1_ASAP7_75t_L g512 ( .A(n_176), .Y(n_512) );
INVx1_ASAP7_75t_L g190 ( .A(n_177), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_179), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_193), .Y(n_179) );
OR2x2_ASAP7_75t_L g311 ( .A(n_180), .B(n_194), .Y(n_311) );
AND2x2_ASAP7_75t_L g348 ( .A(n_180), .B(n_258), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_180), .B(n_279), .Y(n_359) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_180), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_180), .B(n_315), .Y(n_432) );
INVx5_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx2_ASAP7_75t_L g257 ( .A(n_181), .Y(n_257) );
AND2x2_ASAP7_75t_L g266 ( .A(n_181), .B(n_194), .Y(n_266) );
AND2x2_ASAP7_75t_L g382 ( .A(n_181), .B(n_277), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_181), .B(n_315), .Y(n_404) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_191), .Y(n_181) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_194), .Y(n_350) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_195), .Y(n_302) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_L g279 ( .A(n_196), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_206), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_203), .C(n_204), .Y(n_199) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_202), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_202), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g529 ( .A(n_205), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_219), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_210), .B(n_292), .Y(n_411) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_211), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g263 ( .A(n_211), .B(n_264), .Y(n_263) );
INVx5_ASAP7_75t_SL g271 ( .A(n_211), .Y(n_271) );
OR2x2_ASAP7_75t_L g294 ( .A(n_211), .B(n_264), .Y(n_294) );
OR2x2_ASAP7_75t_L g304 ( .A(n_211), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g367 ( .A(n_211), .B(n_221), .Y(n_367) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_211), .B(n_220), .Y(n_405) );
NOR4xp25_ASAP7_75t_L g426 ( .A(n_211), .B(n_347), .C(n_427), .D(n_428), .Y(n_426) );
AND2x2_ASAP7_75t_L g436 ( .A(n_211), .B(n_268), .Y(n_436) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_218), .Y(n_211) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g261 ( .A(n_220), .B(n_257), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_220), .B(n_263), .Y(n_430) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
OR2x2_ASAP7_75t_L g270 ( .A(n_221), .B(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g277 ( .A(n_221), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_221), .B(n_245), .Y(n_289) );
INVxp67_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_221), .B(n_264), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_221), .B(n_231), .Y(n_358) );
AND2x2_ASAP7_75t_L g373 ( .A(n_221), .B(n_268), .Y(n_373) );
OR2x2_ASAP7_75t_L g402 ( .A(n_221), .B(n_231), .Y(n_402) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_229), .Y(n_221) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_222), .A2(n_506), .B(n_513), .Y(n_505) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_222), .A2(n_523), .B(n_530), .Y(n_522) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_222), .A2(n_536), .B(n_542), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_230), .B(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_230), .B(n_271), .Y(n_410) );
OR2x2_ASAP7_75t_L g431 ( .A(n_230), .B(n_308), .Y(n_431) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g244 ( .A(n_231), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g268 ( .A(n_231), .B(n_264), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_231), .B(n_245), .Y(n_283) );
AND2x2_ASAP7_75t_L g353 ( .A(n_231), .B(n_277), .Y(n_353) );
AND2x2_ASAP7_75t_L g387 ( .A(n_231), .B(n_271), .Y(n_387) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_232), .B(n_271), .Y(n_290) );
AND2x2_ASAP7_75t_L g318 ( .A(n_232), .B(n_245), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B(n_240), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_240), .A2(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_243), .B(n_326), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_244), .A2(n_333), .B1(n_369), .B2(n_386), .C(n_388), .Y(n_385) );
INVx5_ASAP7_75t_SL g264 ( .A(n_245), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_249), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_248), .A2(n_471), .B(n_472), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_248), .A2(n_497), .B(n_498), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g459 ( .A(n_255), .Y(n_459) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OAI33xp33_ASAP7_75t_L g284 ( .A1(n_257), .A2(n_285), .A3(n_286), .B1(n_288), .B2(n_291), .B3(n_295), .Y(n_284) );
OR2x2_ASAP7_75t_L g300 ( .A(n_257), .B(n_301), .Y(n_300) );
AOI322xp5_ASAP7_75t_L g409 ( .A1(n_257), .A2(n_326), .A3(n_333), .B1(n_410), .B2(n_411), .C1(n_412), .C2(n_415), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_257), .B(n_285), .Y(n_427) );
A2O1A1Ixp33_ASAP7_75t_SL g433 ( .A1(n_257), .A2(n_285), .B(n_434), .C(n_436), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_258), .A2(n_273), .B1(n_278), .B2(n_281), .C(n_284), .Y(n_272) );
INVx1_ASAP7_75t_L g365 ( .A(n_258), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_258), .B(n_414), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_262), .B1(n_265), .B2(n_267), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g342 ( .A(n_263), .B(n_277), .Y(n_342) );
AND2x2_ASAP7_75t_L g400 ( .A(n_263), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g308 ( .A(n_264), .B(n_271), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_264), .B(n_277), .Y(n_336) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_266), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_266), .B(n_344), .Y(n_398) );
OAI321xp33_ASAP7_75t_L g417 ( .A1(n_266), .A2(n_339), .A3(n_418), .B1(n_419), .B2(n_420), .C(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g384 ( .A(n_267), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_268), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g323 ( .A(n_268), .B(n_271), .Y(n_323) );
AOI321xp33_ASAP7_75t_L g381 ( .A1(n_268), .A2(n_285), .A3(n_382), .B1(n_383), .B2(n_384), .C(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g298 ( .A(n_270), .B(n_283), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_271), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_271), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_271), .B(n_357), .Y(n_394) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g317 ( .A(n_275), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g282 ( .A(n_276), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g390 ( .A(n_277), .Y(n_390) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_280), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_287), .B(n_322), .Y(n_371) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
OR2x2_ASAP7_75t_L g335 ( .A(n_290), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g380 ( .A(n_290), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_291), .A2(n_338), .B1(n_341), .B2(n_343), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g435 ( .A(n_294), .B(n_358), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_299), .B1(n_303), .B2(n_309), .C(n_312), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_SL g379 ( .A(n_305), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_307), .B(n_357), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_307), .A2(n_375), .B(n_377), .Y(n_374) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g420 ( .A(n_308), .B(n_402), .Y(n_420) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_SL g322 ( .A(n_311), .Y(n_322) );
AOI21xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B(n_316), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g366 ( .A(n_318), .B(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g428 ( .A(n_318), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B(n_324), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_322), .B(n_340), .Y(n_376) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g397 ( .A(n_326), .Y(n_397) );
NAND5xp2_ASAP7_75t_L g327 ( .A(n_328), .B(n_345), .C(n_354), .D(n_374), .E(n_381), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B(n_334), .C(n_337), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g369 ( .A(n_333), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_341), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
OAI21xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_349), .B(n_351), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_346), .A2(n_400), .B1(n_403), .B2(n_405), .C(n_406), .Y(n_399) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AOI321xp33_ASAP7_75t_L g354 ( .A1(n_347), .A2(n_355), .A3(n_359), .B1(n_360), .B2(n_366), .C(n_368), .Y(n_354) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g425 ( .A(n_359), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_361), .B(n_365), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g377 ( .A(n_362), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NOR2xp67_ASAP7_75t_SL g389 ( .A(n_363), .B(n_370), .Y(n_389) );
AOI321xp33_ASAP7_75t_SL g421 ( .A1(n_366), .A2(n_422), .A3(n_423), .B1(n_424), .B2(n_425), .C(n_426), .Y(n_421) );
O2A1O1Ixp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B(n_371), .C(n_372), .Y(n_368) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_379), .B(n_387), .Y(n_416) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .C(n_391), .Y(n_388) );
NOR3xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_417), .C(n_429), .Y(n_392) );
OAI211xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_395), .B(n_399), .C(n_409), .Y(n_393) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_398), .A2(n_430), .B1(n_431), .B2(n_432), .C(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g422 ( .A(n_420), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
CKINVDCx14_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g730 ( .A(n_438), .Y(n_730) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_440), .B(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g729 ( .A(n_441), .Y(n_729) );
OR4x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_611), .C(n_658), .D(n_698), .Y(n_441) );
NAND3xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_557), .C(n_586), .Y(n_442) );
AOI211xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_479), .B(n_514), .C(n_550), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_444), .A2(n_570), .B(n_587), .C(n_591), .Y(n_586) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_455), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_446), .B(n_549), .Y(n_548) );
INVx3_ASAP7_75t_SL g553 ( .A(n_446), .Y(n_553) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_446), .Y(n_565) );
AND2x4_ASAP7_75t_L g569 ( .A(n_446), .B(n_521), .Y(n_569) );
AND2x2_ASAP7_75t_L g580 ( .A(n_446), .B(n_469), .Y(n_580) );
OR2x2_ASAP7_75t_L g604 ( .A(n_446), .B(n_517), .Y(n_604) );
AND2x2_ASAP7_75t_L g617 ( .A(n_446), .B(n_522), .Y(n_617) );
AND2x2_ASAP7_75t_L g657 ( .A(n_446), .B(n_643), .Y(n_657) );
AND2x2_ASAP7_75t_L g664 ( .A(n_446), .B(n_627), .Y(n_664) );
AND2x2_ASAP7_75t_L g694 ( .A(n_446), .B(n_456), .Y(n_694) );
OR2x6_ASAP7_75t_L g446 ( .A(n_447), .B(n_453), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_455), .B(n_621), .Y(n_633) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_468), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_456), .B(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g571 ( .A(n_456), .B(n_468), .Y(n_571) );
BUFx3_ASAP7_75t_L g579 ( .A(n_456), .Y(n_579) );
OR2x2_ASAP7_75t_L g600 ( .A(n_456), .B(n_482), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_456), .B(n_621), .Y(n_711) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_460), .B(n_467), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_458), .A2(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g518 ( .A(n_460), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_467), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_468), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g564 ( .A(n_468), .Y(n_564) );
AND2x2_ASAP7_75t_L g627 ( .A(n_468), .B(n_522), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_468), .A2(n_630), .B1(n_632), .B2(n_634), .C(n_635), .Y(n_629) );
AND2x2_ASAP7_75t_L g643 ( .A(n_468), .B(n_517), .Y(n_643) );
AND2x2_ASAP7_75t_L g669 ( .A(n_468), .B(n_553), .Y(n_669) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g549 ( .A(n_469), .B(n_522), .Y(n_549) );
BUFx2_ASAP7_75t_L g683 ( .A(n_469), .Y(n_683) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI32xp33_ASAP7_75t_L g649 ( .A1(n_480), .A2(n_610), .A3(n_624), .B1(n_650), .B2(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
AND2x2_ASAP7_75t_L g590 ( .A(n_481), .B(n_534), .Y(n_590) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g572 ( .A(n_482), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_482), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g644 ( .A(n_482), .B(n_534), .Y(n_644) );
AND2x2_ASAP7_75t_L g655 ( .A(n_482), .B(n_547), .Y(n_655) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g556 ( .A(n_483), .B(n_535), .Y(n_556) );
AND2x2_ASAP7_75t_L g560 ( .A(n_483), .B(n_535), .Y(n_560) );
AND2x2_ASAP7_75t_L g595 ( .A(n_483), .B(n_546), .Y(n_595) );
AND2x2_ASAP7_75t_L g602 ( .A(n_483), .B(n_504), .Y(n_602) );
OAI211xp5_ASAP7_75t_L g607 ( .A1(n_483), .A2(n_553), .B(n_564), .C(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g661 ( .A(n_483), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_483), .B(n_494), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_492), .B(n_544), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_492), .B(n_560), .Y(n_650) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g555 ( .A(n_493), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
AND2x2_ASAP7_75t_L g547 ( .A(n_494), .B(n_505), .Y(n_547) );
OR2x2_ASAP7_75t_L g562 ( .A(n_494), .B(n_505), .Y(n_562) );
AND2x2_ASAP7_75t_L g585 ( .A(n_494), .B(n_546), .Y(n_585) );
INVx1_ASAP7_75t_L g589 ( .A(n_494), .Y(n_589) );
AND2x2_ASAP7_75t_L g608 ( .A(n_494), .B(n_545), .Y(n_608) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_494), .A2(n_573), .B1(n_619), .B2(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_494), .B(n_661), .Y(n_685) );
AND2x2_ASAP7_75t_L g700 ( .A(n_494), .B(n_560), .Y(n_700) );
INVx4_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx3_ASAP7_75t_L g532 ( .A(n_495), .Y(n_532) );
AND2x2_ASAP7_75t_L g574 ( .A(n_495), .B(n_505), .Y(n_574) );
AND2x2_ASAP7_75t_L g576 ( .A(n_495), .B(n_534), .Y(n_576) );
AND3x2_ASAP7_75t_L g638 ( .A(n_495), .B(n_602), .C(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g673 ( .A(n_504), .B(n_545), .Y(n_673) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g534 ( .A(n_505), .B(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_505), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_505), .B(n_544), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_505), .B(n_585), .C(n_661), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_531), .B1(n_543), .B2(n_548), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_520), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_517), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g625 ( .A(n_517), .Y(n_625) );
OAI31xp33_ASAP7_75t_L g641 ( .A1(n_520), .A2(n_642), .A3(n_643), .B(n_644), .Y(n_641) );
AND2x2_ASAP7_75t_L g666 ( .A(n_520), .B(n_553), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_520), .B(n_579), .Y(n_712) );
AND2x2_ASAP7_75t_L g621 ( .A(n_521), .B(n_553), .Y(n_621) );
AND2x2_ASAP7_75t_L g682 ( .A(n_521), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g552 ( .A(n_522), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g610 ( .A(n_522), .Y(n_610) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g631 ( .A(n_532), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_533), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AOI221x1_ASAP7_75t_SL g598 ( .A1(n_534), .A2(n_599), .B1(n_601), .B2(n_603), .C(n_605), .Y(n_598) );
INVx2_ASAP7_75t_L g546 ( .A(n_535), .Y(n_546) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_535), .Y(n_640) );
INVx1_ASAP7_75t_L g628 ( .A(n_543), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_547), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_544), .B(n_561), .Y(n_653) );
INVx1_ASAP7_75t_SL g716 ( .A(n_544), .Y(n_716) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g634 ( .A(n_547), .B(n_560), .Y(n_634) );
INVx1_ASAP7_75t_L g702 ( .A(n_548), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_548), .B(n_631), .Y(n_715) );
INVx2_ASAP7_75t_SL g554 ( .A(n_549), .Y(n_554) );
AND2x2_ASAP7_75t_L g597 ( .A(n_549), .B(n_553), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_549), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_549), .B(n_624), .Y(n_651) );
AOI21xp33_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_554), .B(n_555), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_552), .B(n_624), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_552), .B(n_579), .Y(n_720) );
OR2x2_ASAP7_75t_L g592 ( .A(n_553), .B(n_571), .Y(n_592) );
AND2x2_ASAP7_75t_L g691 ( .A(n_553), .B(n_682), .Y(n_691) );
OAI22xp5_ASAP7_75t_SL g566 ( .A1(n_554), .A2(n_567), .B1(n_572), .B2(n_575), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_554), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g614 ( .A(n_556), .B(n_562), .Y(n_614) );
INVx1_ASAP7_75t_L g678 ( .A(n_556), .Y(n_678) );
AOI311xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_563), .A3(n_565), .B(n_566), .C(n_577), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_561), .A2(n_693), .B1(n_705), .B2(n_708), .C(n_710), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_561), .B(n_716), .Y(n_718) );
INVx2_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g615 ( .A(n_563), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_564), .A2(n_606), .B(n_607), .C(n_609), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
O2A1O1Ixp33_ASAP7_75t_SL g674 ( .A1(n_568), .A2(n_570), .B(n_675), .C(n_676), .Y(n_674) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_569), .B(n_643), .Y(n_709) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g591 ( .A1(n_572), .A2(n_592), .B1(n_593), .B2(n_596), .C(n_598), .Y(n_591) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g594 ( .A(n_574), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g677 ( .A(n_574), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_578), .A2(n_636), .B(n_637), .C(n_641), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_579), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_579), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
INVxp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g601 ( .A(n_585), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_589), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g703 ( .A(n_592), .Y(n_703) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_595), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g630 ( .A(n_595), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g707 ( .A(n_595), .Y(n_707) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g648 ( .A(n_597), .B(n_624), .Y(n_648) );
INVx1_ASAP7_75t_SL g642 ( .A(n_604), .Y(n_642) );
INVx1_ASAP7_75t_L g619 ( .A(n_610), .Y(n_619) );
NAND3xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_629), .C(n_645), .Y(n_611) );
AOI322xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .A3(n_616), .B1(n_618), .B2(n_622), .C1(n_626), .C2(n_628), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_613), .A2(n_666), .B(n_667), .C(n_674), .Y(n_665) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_616), .A2(n_637), .B1(n_668), .B2(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g626 ( .A(n_624), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g663 ( .A(n_624), .B(n_664), .Y(n_663) );
AOI32xp33_ASAP7_75t_L g714 ( .A1(n_624), .A2(n_715), .A3(n_716), .B1(n_717), .B2(n_719), .Y(n_714) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g636 ( .A(n_627), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_627), .A2(n_680), .B1(n_684), .B2(n_686), .C(n_689), .Y(n_679) );
AND2x2_ASAP7_75t_L g693 ( .A(n_627), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g696 ( .A(n_631), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g706 ( .A(n_631), .B(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g697 ( .A(n_640), .B(n_661), .Y(n_697) );
AOI211xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_648), .B(n_649), .C(n_652), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI21xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI211xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_662), .B(n_665), .C(n_679), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_673), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g688 ( .A(n_685), .Y(n_688) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B(n_695), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_701), .B(n_704), .C(n_714), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g731 ( .A(n_721), .Y(n_731) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
BUFx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g752 ( .A(n_742), .Y(n_752) );
INVx1_ASAP7_75t_L g750 ( .A(n_744), .Y(n_750) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g759 ( .A(n_755), .Y(n_759) );
INVx1_ASAP7_75t_SL g765 ( .A(n_755), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g767 ( .A(n_761), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_765), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
endmodule