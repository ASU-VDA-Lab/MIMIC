module fake_jpeg_26733_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_0),
.B(n_1),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_39),
.B(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_50),
.Y(n_85)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_16),
.B1(n_25),
.B2(n_22),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_69),
.B1(n_36),
.B2(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_27),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_30),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_43),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_16),
.B1(n_22),
.B2(n_26),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_21),
.B(n_18),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_27),
.B(n_44),
.C(n_21),
.Y(n_89)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_16),
.B1(n_26),
.B2(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_78),
.B1(n_81),
.B2(n_47),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_36),
.B1(n_42),
.B2(n_40),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_87),
.B1(n_89),
.B2(n_35),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_76),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_26),
.B1(n_31),
.B2(n_23),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_19),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_83),
.Y(n_98)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_37),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_40),
.B1(n_37),
.B2(n_35),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_44),
.Y(n_119)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_95),
.Y(n_106)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_52),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_96),
.A2(n_81),
.B(n_95),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_105),
.Y(n_128)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_113),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_119),
.B(n_91),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_80),
.Y(n_112)
);

BUFx4f_ASAP7_75t_SL g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_53),
.C(n_55),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_82),
.C(n_76),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_77),
.B(n_31),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_53),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_60),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_146),
.B(n_150),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_91),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_91),
.B1(n_82),
.B2(n_74),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_98),
.B1(n_113),
.B2(n_111),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_149),
.Y(n_171)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_148),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_116),
.C(n_109),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_83),
.B(n_70),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_96),
.B1(n_81),
.B2(n_71),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_104),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_154),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_153),
.A2(n_92),
.B1(n_68),
.B2(n_65),
.Y(n_204)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_100),
.B(n_108),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_175),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_108),
.B(n_119),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_157),
.B(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_165),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_145),
.B(n_116),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_109),
.B(n_79),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_164),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_148),
.C(n_144),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_109),
.B(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_129),
.B1(n_102),
.B2(n_127),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_105),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_131),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_61),
.B1(n_60),
.B2(n_71),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_173),
.B1(n_97),
.B2(n_102),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_70),
.B1(n_92),
.B2(n_49),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_29),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_140),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_186),
.C(n_203),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_187),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_131),
.C(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_151),
.B1(n_154),
.B2(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_194),
.B1(n_170),
.B2(n_168),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_128),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_199),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_29),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_201),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_49),
.B1(n_143),
.B2(n_88),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_204),
.B1(n_176),
.B2(n_102),
.Y(n_214)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_152),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_125),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_135),
.C(n_126),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_112),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_51),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_156),
.B(n_177),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_216),
.B(n_192),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_214),
.A2(n_215),
.B1(n_225),
.B2(n_212),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_155),
.B1(n_157),
.B2(n_165),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_180),
.A2(n_164),
.B(n_155),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_218),
.A2(n_228),
.B1(n_230),
.B2(n_44),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_174),
.C(n_170),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_197),
.C(n_192),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_205),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_132),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_178),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_226),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_135),
.B1(n_126),
.B2(n_120),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_125),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_227),
.B(n_24),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_188),
.A2(n_183),
.B1(n_182),
.B2(n_202),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_44),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_132),
.B1(n_86),
.B2(n_84),
.Y(n_230)
);

AO22x1_ASAP7_75t_L g231 ( 
.A1(n_208),
.A2(n_190),
.B1(n_204),
.B2(n_179),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_237),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_240),
.C(n_244),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_226),
.Y(n_237)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_50),
.B(n_19),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_211),
.B(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_158),
.C(n_86),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_84),
.B1(n_94),
.B2(n_32),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_94),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_243),
.B(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_44),
.C(n_21),
.Y(n_244)
);

INVxp33_ASAP7_75t_SL g245 ( 
.A(n_229),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_245),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_24),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_249),
.C(n_252),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_247),
.A2(n_210),
.B1(n_207),
.B2(n_224),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_220),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_17),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_24),
.CI(n_17),
.CON(n_251),
.SN(n_251)
);

OAI321xp33_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_222),
.A3(n_206),
.B1(n_215),
.B2(n_227),
.C(n_207),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_33),
.C(n_32),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_206),
.B1(n_213),
.B2(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_231),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_237),
.B1(n_210),
.B2(n_235),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_267),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_225),
.C(n_32),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_252),
.C(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_245),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_269),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_283),
.C(n_258),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_233),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_265),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_236),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_249),
.B1(n_246),
.B2(n_17),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_282),
.B1(n_6),
.B2(n_13),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_7),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_9),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_254),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_9),
.C(n_13),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_292),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_261),
.B(n_255),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_290),
.B(n_283),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_255),
.B(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_282),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_267),
.B(n_254),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_294),
.B(n_5),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_269),
.B(n_253),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_14),
.B(n_6),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_295),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_271),
.B(n_279),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_306),
.B(n_293),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_273),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_291),
.B(n_10),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_5),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_310),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_285),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_312),
.A2(n_315),
.B(n_11),
.C(n_12),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_14),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_5),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_2),
.B(n_3),
.Y(n_319)
);

OAI211xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_317),
.B(n_319),
.C(n_3),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_SL g317 ( 
.A(n_308),
.B(n_12),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_311),
.C(n_308),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_SL g323 ( 
.A(n_321),
.B(n_322),
.C(n_316),
.Y(n_323)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_318),
.B(n_4),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_4),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_4),
.Y(n_326)
);


endmodule