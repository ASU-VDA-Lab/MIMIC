module fake_jpeg_16517_n_321 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx9p33_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_22),
.B1(n_28),
.B2(n_20),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_54),
.B1(n_36),
.B2(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_20),
.B1(n_28),
.B2(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_61),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_36),
.B1(n_31),
.B2(n_37),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_70),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_36),
.B1(n_20),
.B2(n_28),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_51),
.B1(n_31),
.B2(n_14),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_39),
.B1(n_33),
.B2(n_37),
.Y(n_76)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_38),
.B1(n_33),
.B2(n_48),
.Y(n_96)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_52),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_21),
.B(n_16),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_14),
.B1(n_18),
.B2(n_16),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_28),
.B1(n_19),
.B2(n_27),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_82)
);

OAI22x1_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_19),
.B1(n_24),
.B2(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_93),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_94),
.B1(n_96),
.B2(n_105),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_47),
.B1(n_37),
.B2(n_31),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_92),
.B1(n_59),
.B2(n_77),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_37),
.B1(n_31),
.B2(n_33),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_99),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_73),
.B(n_79),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_60),
.Y(n_110)
);

OA22x2_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_38),
.B1(n_40),
.B2(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_83),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_124),
.B1(n_85),
.B2(n_128),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_123),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_120),
.B(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_74),
.B1(n_73),
.B2(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_68),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_91),
.A2(n_99),
.B1(n_93),
.B2(n_86),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_127),
.B1(n_130),
.B2(n_107),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_76),
.C(n_77),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_40),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_69),
.B1(n_67),
.B2(n_58),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_76),
.B1(n_38),
.B2(n_40),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_89),
.B1(n_96),
.B2(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_76),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_105),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_50),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_50),
.Y(n_151)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_137),
.A2(n_138),
.B(n_149),
.Y(n_192)
);

XOR2x2_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_107),
.B1(n_101),
.B2(n_108),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_147),
.B1(n_156),
.B2(n_160),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_144),
.B1(n_114),
.B2(n_23),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_130),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_142),
.B(n_145),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_108),
.B1(n_100),
.B2(n_102),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_100),
.B1(n_106),
.B2(n_87),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_109),
.B(n_106),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_53),
.C(n_40),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_155),
.C(n_17),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_152),
.A2(n_163),
.B1(n_21),
.B2(n_64),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_18),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_30),
.B1(n_24),
.B2(n_53),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_123),
.B(n_65),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_68),
.C(n_65),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_18),
.B1(n_16),
.B2(n_25),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_17),
.Y(n_159)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_11),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_0),
.B(n_1),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_112),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_164),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_126),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_169),
.A2(n_182),
.B(n_188),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_125),
.B(n_122),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_171),
.A2(n_156),
.B(n_160),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_29),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_127),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_183),
.C(n_191),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_184),
.B1(n_190),
.B2(n_196),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_179),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_136),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_121),
.B1(n_112),
.B2(n_123),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_193),
.B1(n_195),
.B2(n_149),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_112),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_17),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_154),
.A2(n_17),
.B1(n_29),
.B2(n_66),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_155),
.B(n_42),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_154),
.A2(n_29),
.B1(n_8),
.B2(n_2),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_8),
.B1(n_12),
.B2(n_3),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_137),
.A2(n_144),
.B(n_140),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_154),
.B1(n_147),
.B2(n_139),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_207),
.B1(n_176),
.B2(n_173),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_204),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_168),
.B(n_148),
.CI(n_159),
.CON(n_205),
.SN(n_205)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_182),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_150),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_210),
.C(n_215),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_172),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_161),
.B1(n_145),
.B2(n_143),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_211),
.A2(n_213),
.B1(n_180),
.B2(n_181),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_198),
.A2(n_143),
.B1(n_136),
.B2(n_158),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_158),
.C(n_161),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_175),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_169),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_8),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g228 ( 
.A(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_228),
.B(n_233),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_221),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_231),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_177),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_197),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_170),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_240),
.B1(n_242),
.B2(n_217),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_184),
.B1(n_176),
.B2(n_189),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_203),
.B1(n_169),
.B2(n_209),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_192),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_241),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_189),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_180),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_167),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_245),
.A2(n_200),
.B(n_167),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_215),
.C(n_212),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_253),
.C(n_256),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_209),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_260),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_212),
.C(n_208),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_260),
.B1(n_232),
.B2(n_227),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_211),
.B(n_188),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_223),
.C(n_205),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_261),
.B1(n_232),
.B2(n_244),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_217),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_247),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_205),
.C(n_222),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_263),
.C(n_231),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_195),
.B1(n_193),
.B2(n_3),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_42),
.C(n_29),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_252),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_268),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_234),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_250),
.C(n_248),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_253),
.C(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_274),
.C(n_275),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_259),
.C(n_258),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_241),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_233),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_277),
.C(n_266),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_230),
.C(n_244),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_278),
.A2(n_263),
.B1(n_243),
.B2(n_3),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_282),
.B1(n_275),
.B2(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_9),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_276),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_243),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_29),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_7),
.B1(n_13),
.B2(n_3),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_289),
.B1(n_10),
.B2(n_12),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_290),
.Y(n_293)
);

OAI321xp33_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_9),
.A3(n_13),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_29),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_264),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_264),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_296),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_7),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_283),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_299),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_300),
.B1(n_0),
.B2(n_1),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_274),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_285),
.C(n_286),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_305),
.C(n_300),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_285),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_282),
.B1(n_7),
.B2(n_4),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.C(n_5),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_311),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_5),
.C(n_6),
.Y(n_311)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_308),
.B(n_304),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_302),
.Y(n_315)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_313),
.C(n_310),
.Y(n_316)
);

OAI211xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_5),
.B(n_10),
.C(n_11),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_11),
.B(n_12),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_12),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_0),
.B(n_1),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_1),
.C(n_311),
.Y(n_321)
);


endmodule