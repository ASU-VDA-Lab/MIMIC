module fake_jpeg_12465_n_532 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_532);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_532;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_76),
.Y(n_113)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_55),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_85),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_93),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_94),
.B(n_96),
.Y(n_155)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_30),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_101),
.Y(n_123)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_21),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_111),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_131),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_85),
.A2(n_28),
.B1(n_37),
.B2(n_32),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_125),
.A2(n_127),
.B1(n_128),
.B2(n_138),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_28),
.B1(n_36),
.B2(n_45),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_28),
.B1(n_36),
.B2(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_54),
.B(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_133),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_52),
.A2(n_38),
.B1(n_24),
.B2(n_43),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_130),
.A2(n_140),
.B1(n_157),
.B2(n_39),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_64),
.A2(n_83),
.B1(n_65),
.B2(n_58),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_131),
.A2(n_149),
.B1(n_158),
.B2(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_24),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_66),
.A2(n_36),
.B1(n_31),
.B2(n_45),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_77),
.A2(n_36),
.B1(n_31),
.B2(n_45),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_38),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_161),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_102),
.A2(n_21),
.B1(n_31),
.B2(n_43),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_99),
.A2(n_31),
.B1(n_41),
.B2(n_43),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_53),
.A2(n_41),
.B1(n_43),
.B2(n_38),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_96),
.B(n_49),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_59),
.A2(n_41),
.B1(n_49),
.B2(n_39),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_60),
.A2(n_41),
.B1(n_46),
.B2(n_44),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_44),
.B1(n_25),
.B2(n_29),
.Y(n_195)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_165),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_33),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_169),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_167),
.B(n_215),
.Y(n_266)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_110),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_108),
.A2(n_101),
.B1(n_69),
.B2(n_68),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_170),
.A2(n_171),
.B1(n_195),
.B2(n_222),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_108),
.A2(n_80),
.B1(n_72),
.B2(n_75),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_172),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_182),
.Y(n_227)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_179),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_100),
.C(n_91),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_186),
.C(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_39),
.Y(n_183)
);

NOR2xp67_ASAP7_75t_R g240 ( 
.A(n_183),
.B(n_187),
.Y(n_240)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_184),
.Y(n_262)
);

AO22x2_ASAP7_75t_L g185 ( 
.A1(n_106),
.A2(n_82),
.B1(n_74),
.B2(n_57),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_185),
.B(n_216),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_94),
.C(n_90),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_107),
.B(n_49),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_120),
.Y(n_190)
);

OR2x4_ASAP7_75t_L g191 ( 
.A(n_107),
.B(n_117),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_191),
.A2(n_0),
.B(n_1),
.Y(n_260)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_198),
.Y(n_249)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_194),
.A2(n_136),
.B1(n_150),
.B2(n_148),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_119),
.B(n_56),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_119),
.B(n_22),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_123),
.A2(n_71),
.B1(n_44),
.B2(n_25),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_200),
.A2(n_208),
.B1(n_210),
.B2(n_213),
.Y(n_232)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_202),
.Y(n_235)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_22),
.B(n_25),
.C(n_29),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_205),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_108),
.B(n_56),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_206),
.B(n_207),
.C(n_0),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_0),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_116),
.A2(n_46),
.B1(n_29),
.B2(n_22),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_106),
.A2(n_95),
.B1(n_55),
.B2(n_46),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_214),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_105),
.B(n_33),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_217),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_116),
.A2(n_33),
.B1(n_34),
.B2(n_11),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_105),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_114),
.B(n_11),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_115),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_218),
.Y(n_230)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_219),
.A2(n_220),
.B1(n_147),
.B2(n_122),
.Y(n_238)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_114),
.B(n_11),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_221),
.B(n_17),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_122),
.A2(n_33),
.B1(n_34),
.B2(n_11),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_112),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_234),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_231),
.A2(n_203),
.B1(n_195),
.B2(n_197),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_176),
.B(n_134),
.Y(n_234)
);

AOI32xp33_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_136),
.A3(n_109),
.B1(n_153),
.B2(n_132),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_237),
.A2(n_245),
.B(n_260),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_238),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_153),
.B1(n_132),
.B2(n_150),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_241),
.A2(n_261),
.B1(n_177),
.B2(n_218),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_189),
.A2(n_121),
.B1(n_148),
.B2(n_146),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_244),
.A2(n_253),
.B1(n_268),
.B2(n_235),
.Y(n_285)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_191),
.A2(n_121),
.A3(n_34),
.B1(n_144),
.B2(n_126),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_186),
.A2(n_12),
.B(n_18),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_254),
.C(n_204),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_154),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_264),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_189),
.A2(n_154),
.B1(n_146),
.B2(n_144),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_7),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_207),
.C(n_206),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_200),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_207),
.B(n_1),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_167),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_SL g293 ( 
.A1(n_265),
.A2(n_267),
.B(n_173),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_167),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_269),
.B(n_227),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_2),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_255),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_276),
.B(n_278),
.Y(n_352)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_224),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_277),
.Y(n_342)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_282),
.A2(n_312),
.B1(n_240),
.B2(n_245),
.Y(n_331)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_249),
.B(n_180),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_284),
.B(n_286),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_285),
.A2(n_291),
.B1(n_292),
.B2(n_296),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_249),
.B(n_226),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_225),
.A2(n_185),
.B1(n_215),
.B2(n_193),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_287),
.A2(n_289),
.B1(n_293),
.B2(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_225),
.A2(n_185),
.B1(n_178),
.B2(n_164),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_236),
.Y(n_290)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_290),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_244),
.A2(n_210),
.B1(n_208),
.B2(n_185),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_253),
.A2(n_196),
.B1(n_199),
.B2(n_201),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_227),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_294),
.B(n_298),
.Y(n_349)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_236),
.Y(n_295)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

AO21x2_ASAP7_75t_L g296 ( 
.A1(n_251),
.A2(n_165),
.B(n_217),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_233),
.B(n_234),
.Y(n_298)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_229),
.B(n_196),
.C(n_209),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_254),
.C(n_260),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_229),
.A2(n_184),
.B(n_175),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_302),
.A2(n_305),
.B(n_319),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_263),
.B(n_172),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_303),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_179),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_168),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_246),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_309),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_310),
.B(n_262),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_266),
.A2(n_219),
.B1(n_211),
.B2(n_220),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_313),
.B1(n_247),
.B2(n_228),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_237),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_266),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_248),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_316),
.Y(n_328)
);

CKINVDCx12_ASAP7_75t_R g315 ( 
.A(n_263),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_2),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_230),
.B(n_14),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_318),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_230),
.B(n_2),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_256),
.B(n_3),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_320),
.A2(n_331),
.B1(n_343),
.B2(n_350),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_285),
.A2(n_231),
.B1(n_232),
.B2(n_240),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_323),
.A2(n_346),
.B1(n_315),
.B2(n_297),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_354),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_333),
.C(n_334),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_282),
.A2(n_270),
.B1(n_232),
.B2(n_256),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_252),
.C(n_258),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_252),
.C(n_258),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_250),
.C(n_242),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_356),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_319),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_340),
.B(n_281),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_287),
.A2(n_271),
.B1(n_273),
.B2(n_243),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_306),
.A2(n_242),
.B(n_247),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_345),
.A2(n_360),
.B(n_305),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_296),
.A2(n_271),
.B1(n_250),
.B2(n_273),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_289),
.A2(n_243),
.B1(n_262),
.B2(n_228),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_294),
.A2(n_262),
.B1(n_259),
.B2(n_5),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_353),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_284),
.B(n_3),
.C(n_4),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_274),
.B(n_3),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_275),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_276),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_361),
.A2(n_377),
.B1(n_378),
.B2(n_383),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_331),
.A2(n_296),
.B1(n_297),
.B2(n_274),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_362),
.A2(n_392),
.B1(n_357),
.B2(n_348),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_336),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_364),
.B(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_335),
.Y(n_368)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_341),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_354),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_371),
.B(n_379),
.C(n_333),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_349),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_372),
.B(n_375),
.Y(n_420)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_346),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_334),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_339),
.A2(n_279),
.B1(n_314),
.B2(n_296),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_339),
.A2(n_279),
.B1(n_296),
.B2(n_310),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_275),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_352),
.B(n_286),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_380),
.B(n_382),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_381),
.A2(n_351),
.B(n_393),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_321),
.B(n_288),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_323),
.A2(n_296),
.B1(n_280),
.B2(n_304),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_322),
.A2(n_308),
.B1(n_291),
.B2(n_316),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_384),
.A2(n_388),
.B1(n_389),
.B2(n_361),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_322),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_385),
.B(n_326),
.Y(n_426)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_337),
.A2(n_292),
.B1(n_309),
.B2(n_307),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_332),
.A2(n_295),
.B1(n_290),
.B2(n_283),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_320),
.A2(n_278),
.B1(n_318),
.B2(n_317),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_321),
.B(n_277),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_394),
.B(n_395),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_396),
.B(n_403),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_369),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_397),
.B(n_407),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_391),
.Y(n_398)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_398),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_371),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_401),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_366),
.B(n_327),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_404),
.A2(n_411),
.B1(n_414),
.B2(n_370),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_328),
.C(n_344),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_409),
.C(n_365),
.Y(n_428)
);

OAI22x1_ASAP7_75t_L g407 ( 
.A1(n_383),
.A2(n_345),
.B1(n_338),
.B2(n_329),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_328),
.C(n_344),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_325),
.Y(n_410)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_410),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_378),
.A2(n_338),
.B1(n_329),
.B2(n_340),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_377),
.A2(n_343),
.B1(n_350),
.B2(n_347),
.Y(n_414)
);

NAND4xp25_ASAP7_75t_SL g415 ( 
.A(n_364),
.B(n_351),
.C(n_325),
.D(n_300),
.Y(n_415)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

AND2x2_ASAP7_75t_SL g435 ( 
.A(n_417),
.B(n_389),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_379),
.B(n_347),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_424),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_369),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_422),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_356),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_425),
.A2(n_393),
.B1(n_384),
.B2(n_381),
.Y(n_430)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_428),
.B(n_429),
.C(n_444),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_365),
.C(n_388),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_440),
.B1(n_452),
.B2(n_414),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_362),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_441),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_426),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_432),
.B(n_442),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_434),
.A2(n_437),
.B1(n_448),
.B2(n_449),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_439),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_375),
.B1(n_385),
.B2(n_392),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_403),
.B(n_368),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_425),
.A2(n_363),
.B1(n_394),
.B2(n_367),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_396),
.B(n_390),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_420),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_387),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_404),
.A2(n_363),
.B1(n_373),
.B2(n_374),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_411),
.A2(n_358),
.B1(n_326),
.B2(n_342),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_401),
.B(n_358),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_450),
.B(n_402),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_420),
.A2(n_360),
.B1(n_342),
.B2(n_6),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_451),
.Y(n_455)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_438),
.Y(n_457)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_457),
.Y(n_490)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_438),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_458),
.A2(n_460),
.B1(n_472),
.B2(n_419),
.Y(n_481)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_461),
.A2(n_418),
.B1(n_419),
.B2(n_416),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_434),
.A2(n_407),
.B1(n_413),
.B2(n_422),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_464),
.A2(n_467),
.B1(n_471),
.B2(n_473),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_428),
.B(n_409),
.C(n_424),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_466),
.C(n_443),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_429),
.B(n_413),
.C(n_417),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_437),
.A2(n_397),
.B1(n_405),
.B2(n_398),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_427),
.B(n_405),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_469),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_446),
.A2(n_449),
.B(n_435),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_470),
.A2(n_435),
.B(n_430),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_446),
.A2(n_423),
.B1(n_412),
.B2(n_408),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_448),
.A2(n_423),
.B1(n_412),
.B2(n_408),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_431),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_479),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_466),
.A2(n_450),
.B(n_415),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_475),
.B(n_478),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_443),
.Y(n_479)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_473),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_463),
.B(n_444),
.C(n_447),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_483),
.C(n_485),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_463),
.B(n_447),
.C(n_433),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_484),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_433),
.C(n_441),
.Y(n_485)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_460),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_454),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_472),
.C(n_439),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_459),
.C(n_471),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_477),
.A2(n_470),
.B(n_453),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_501),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_458),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_492),
.B(n_495),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_477),
.A2(n_461),
.B1(n_455),
.B2(n_468),
.Y(n_494)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_494),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_499),
.B(n_500),
.Y(n_512)
);

OAI321xp33_ASAP7_75t_L g500 ( 
.A1(n_488),
.A2(n_490),
.A3(n_484),
.B1(n_476),
.B2(n_457),
.C(n_464),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_480),
.A2(n_489),
.B1(n_462),
.B2(n_467),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_4),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_486),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_SL g513 ( 
.A1(n_504),
.A2(n_452),
.B1(n_418),
.B2(n_342),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_502),
.A2(n_478),
.B(n_485),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_506),
.A2(n_493),
.B(n_503),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_498),
.A2(n_483),
.B(n_482),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_511),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_496),
.B(n_462),
.Y(n_510)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_510),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_498),
.A2(n_479),
.B(n_474),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_513),
.B(n_514),
.Y(n_519)
);

AOI21xp33_ASAP7_75t_L g515 ( 
.A1(n_512),
.A2(n_496),
.B(n_491),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_515),
.B(n_520),
.Y(n_524)
);

A2O1A1O1Ixp25_ASAP7_75t_L g518 ( 
.A1(n_508),
.A2(n_499),
.B(n_497),
.C(n_494),
.D(n_493),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_518),
.A2(n_509),
.B(n_510),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_519),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_521),
.A2(n_522),
.B(n_523),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_516),
.A2(n_509),
.B(n_505),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_524),
.A2(n_517),
.B(n_518),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_4),
.C(n_5),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_525),
.A2(n_513),
.B(n_514),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_527),
.A2(n_528),
.B1(n_4),
.B2(n_5),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_6),
.Y(n_530)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_530),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_6),
.Y(n_532)
);


endmodule