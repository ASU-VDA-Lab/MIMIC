module fake_jpeg_5099_n_177 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_20),
.A2(n_3),
.B(n_4),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_35),
.Y(n_40)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_30),
.A2(n_15),
.B1(n_17),
.B2(n_25),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_15),
.B1(n_17),
.B2(n_13),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_14),
.Y(n_46)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_64),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_15),
.B1(n_13),
.B2(n_33),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_23),
.B(n_19),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_40),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_45),
.B(n_43),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_62),
.C(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_77),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_35),
.B1(n_33),
.B2(n_50),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_83),
.B1(n_35),
.B2(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_80),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_51),
.B1(n_33),
.B2(n_35),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_91),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_66),
.B1(n_67),
.B2(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_74),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_57),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_116),
.C(n_87),
.Y(n_118)
);

AOI221xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_74),
.B1(n_84),
.B2(n_79),
.C(n_81),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_110),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_76),
.B1(n_83),
.B2(n_46),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_25),
.C(n_14),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_24),
.C(n_16),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_82),
.B1(n_63),
.B2(n_40),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_128),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_121),
.Y(n_133)
);

AOI321xp33_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_32),
.A3(n_20),
.B1(n_36),
.B2(n_39),
.C(n_48),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_96),
.C(n_89),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_129),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_88),
.A3(n_91),
.B1(n_99),
.B2(n_94),
.C(n_32),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_115),
.A3(n_110),
.B1(n_130),
.B2(n_104),
.C1(n_120),
.C2(n_109),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_106),
.C(n_107),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_107),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_104),
.B(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_24),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_63),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_131),
.A2(n_137),
.B(n_141),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_140),
.B(n_142),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_16),
.C(n_26),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_57),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_142),
.B(n_132),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_124),
.B1(n_122),
.B2(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_58),
.B1(n_56),
.B2(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_36),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_136),
.B(n_36),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_26),
.B(n_23),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_147),
.C(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_4),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_152),
.B(n_12),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_52),
.B1(n_27),
.B2(n_21),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_16),
.C(n_52),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_135),
.C(n_139),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_52),
.B1(n_27),
.B2(n_21),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_5),
.C(n_6),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_27),
.B1(n_21),
.B2(n_12),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_158),
.C(n_9),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_5),
.B(n_6),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_26),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_164),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_23),
.B(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_16),
.C(n_10),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_156),
.B(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_159),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_9),
.B(n_10),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_11),
.C(n_173),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_168),
.B(n_9),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);


endmodule