module fake_jpeg_29535_n_411 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_411);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_12),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_3),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_47),
.B(n_55),
.Y(n_126)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_52),
.Y(n_94)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_26),
.B(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_61),
.Y(n_127)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_71),
.Y(n_87)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_86)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_83),
.B1(n_30),
.B2(n_20),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_85),
.B(n_102),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_20),
.B1(n_30),
.B2(n_35),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_93),
.A2(n_63),
.B1(n_76),
.B2(n_54),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_45),
.A2(n_30),
.B1(n_22),
.B2(n_31),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_96),
.A2(n_100),
.B1(n_113),
.B2(n_117),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_123),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_51),
.A2(n_30),
.B1(n_22),
.B2(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_41),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_41),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_121),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_64),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_67),
.A2(n_28),
.B1(n_41),
.B2(n_34),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_34),
.C(n_27),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_21),
.C(n_27),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_41),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_16),
.B(n_13),
.C(n_14),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_139),
.Y(n_190)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_88),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_138),
.B(n_140),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_73),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_91),
.A2(n_69),
.B1(n_68),
.B2(n_75),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_145),
.B1(n_87),
.B2(n_84),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_146),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_159),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_75),
.B1(n_74),
.B2(n_81),
.Y(n_148)
);

OAI22x1_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_93),
.B1(n_21),
.B2(n_34),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_71),
.B(n_73),
.C(n_21),
.Y(n_149)
);

NOR2x1_ASAP7_75t_R g182 ( 
.A(n_149),
.B(n_27),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_103),
.C(n_119),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_98),
.A2(n_71),
.B1(n_74),
.B2(n_27),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_125),
.A3(n_112),
.B1(n_103),
.B2(n_124),
.Y(n_185)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_156),
.Y(n_189)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_157),
.B(n_162),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_27),
.B1(n_34),
.B2(n_21),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_87),
.B1(n_105),
.B2(n_102),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_95),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_160),
.B(n_161),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_87),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_107),
.B1(n_111),
.B2(n_106),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_170),
.B1(n_173),
.B2(n_183),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_151),
.B1(n_91),
.B2(n_110),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_166),
.A2(n_175),
.B1(n_186),
.B2(n_149),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_85),
.B(n_94),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_134),
.B(n_126),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_182),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_110),
.B1(n_109),
.B2(n_114),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_109),
.B1(n_114),
.B2(n_97),
.Y(n_183)
);

AOI22x1_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_149),
.B1(n_157),
.B2(n_153),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_107),
.B1(n_111),
.B2(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_135),
.B(n_112),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_135),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_149),
.C(n_137),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_196),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_152),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_200),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_128),
.B1(n_159),
.B2(n_158),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_202),
.B1(n_220),
.B2(n_184),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_184),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_168),
.B(n_134),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_201),
.A2(n_212),
.B(n_140),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_183),
.B1(n_170),
.B2(n_174),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_169),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_150),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_206),
.C(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_185),
.B(n_180),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_209),
.B1(n_217),
.B2(n_213),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_149),
.B1(n_162),
.B2(n_143),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_146),
.B(n_164),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_214),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_132),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_177),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_166),
.A2(n_156),
.B1(n_133),
.B2(n_144),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_136),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_174),
.A2(n_138),
.B1(n_161),
.B2(n_124),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_186),
.B1(n_175),
.B2(n_193),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_237),
.B1(n_240),
.B2(n_244),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_225),
.B(n_13),
.CI(n_12),
.CON(n_270),
.SN(n_270)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_199),
.B1(n_207),
.B2(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_231),
.C(n_238),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_233),
.B1(n_243),
.B2(n_220),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_190),
.C(n_180),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_195),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_208),
.B1(n_213),
.B2(n_217),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_171),
.B(n_179),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_236),
.A2(n_246),
.B(n_0),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_177),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_202),
.A2(n_188),
.B1(n_167),
.B2(n_178),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_172),
.C(n_178),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_211),
.C(n_215),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_184),
.B1(n_181),
.B2(n_187),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_187),
.B1(n_191),
.B2(n_181),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_194),
.A2(n_199),
.B1(n_213),
.B2(n_201),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_247),
.B1(n_215),
.B2(n_210),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_194),
.A2(n_140),
.B1(n_130),
.B2(n_108),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_249),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_237),
.A2(n_200),
.B1(n_218),
.B2(n_212),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_250),
.A2(n_243),
.B(n_235),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_253),
.B1(n_262),
.B2(n_267),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_201),
.B(n_203),
.C(n_216),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_252),
.B(n_268),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_230),
.A2(n_207),
.B1(n_219),
.B2(n_197),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_205),
.Y(n_257)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_223),
.B(n_207),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_260),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_241),
.C(n_222),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_215),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_17),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_269),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_233),
.A2(n_211),
.B1(n_16),
.B2(n_13),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_228),
.B(n_16),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_242),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_270),
.B(n_275),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_273),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_0),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_276),
.Y(n_299)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_1),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_224),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_227),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_281),
.C(n_293),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_236),
.Y(n_281)
);

XOR2x2_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_246),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_SL g311 ( 
.A(n_283),
.B(n_284),
.C(n_285),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_262),
.A2(n_245),
.B(n_260),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_268),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_238),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_259),
.B(n_226),
.Y(n_294)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_231),
.Y(n_295)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_250),
.B(n_225),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_247),
.C(n_226),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_253),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_278),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_258),
.B1(n_273),
.B2(n_249),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_307),
.A2(n_315),
.B1(n_320),
.B2(n_284),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_251),
.B1(n_285),
.B2(n_286),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_309),
.B(n_313),
.Y(n_346)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_267),
.B1(n_258),
.B2(n_249),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_282),
.A2(n_249),
.B1(n_248),
.B2(n_264),
.Y(n_315)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_316),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_257),
.Y(n_317)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_317),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_249),
.C(n_269),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_283),
.C(n_298),
.Y(n_330)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_277),
.B1(n_226),
.B2(n_254),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_322),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_304),
.A2(n_255),
.B1(n_271),
.B2(n_272),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_274),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_324),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_266),
.B1(n_276),
.B2(n_234),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_326),
.Y(n_341)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_300),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_330),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_302),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_336),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_293),
.C(n_283),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_338),
.C(n_343),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_332),
.A2(n_313),
.B1(n_309),
.B2(n_310),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_306),
.B(n_289),
.CI(n_287),
.CON(n_333),
.SN(n_333)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_333),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_311),
.A2(n_289),
.B1(n_294),
.B2(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_305),
.B(n_299),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_299),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_322),
.C(n_317),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_305),
.B(n_270),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_345),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_346),
.A2(n_311),
.B(n_308),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_350),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_334),
.A2(n_307),
.B1(n_315),
.B2(n_320),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_352),
.A2(n_357),
.B1(n_358),
.B2(n_360),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_354),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_324),
.C(n_280),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_338),
.C(n_330),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_340),
.A2(n_292),
.B1(n_290),
.B2(n_297),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_335),
.A2(n_290),
.B1(n_297),
.B2(n_270),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_344),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_361),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_337),
.A2(n_332),
.B(n_346),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_362),
.A2(n_339),
.B(n_3),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_365),
.Y(n_377)
);

FAx1_ASAP7_75t_SL g364 ( 
.A(n_357),
.B(n_331),
.CI(n_333),
.CON(n_364),
.SN(n_364)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_364),
.B(n_351),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_327),
.C(n_328),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_333),
.C(n_342),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_370),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_358),
.Y(n_376)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_349),
.Y(n_370)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_359),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_374),
.Y(n_379)
);

OAI321xp33_ASAP7_75t_L g374 ( 
.A1(n_362),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_8),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_350),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_376),
.B(n_382),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_368),
.A2(n_352),
.B1(n_356),
.B2(n_351),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_380),
.A2(n_371),
.B1(n_367),
.B2(n_364),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_355),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_386),
.C(n_6),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_366),
.A2(n_356),
.B(n_347),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_383),
.A2(n_384),
.B(n_6),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_363),
.A2(n_347),
.B(n_354),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_6),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_360),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_388),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_365),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_379),
.A2(n_1),
.B(n_4),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_389),
.A2(n_392),
.B(n_8),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_5),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_376),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_393),
.B(n_394),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_R g395 ( 
.A(n_378),
.B(n_8),
.Y(n_395)
);

OAI21xp33_ASAP7_75t_L g400 ( 
.A1(n_395),
.A2(n_9),
.B(n_10),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_396),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_397),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_SL g402 ( 
.A1(n_400),
.A2(n_390),
.B(n_389),
.C(n_11),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_381),
.Y(n_401)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_401),
.A2(n_386),
.B(n_10),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_402),
.A2(n_9),
.B(n_10),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_405),
.A2(n_399),
.B(n_404),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_407),
.C(n_403),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_398),
.C(n_10),
.Y(n_409)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_409),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_11),
.Y(n_411)
);


endmodule