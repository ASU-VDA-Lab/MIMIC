module fake_netlist_5_1380_n_1829 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1829);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1829;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_SL g182 ( 
.A(n_49),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_65),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_37),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_70),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_31),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_49),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_58),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_47),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_142),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_63),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_6),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_36),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_18),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_7),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_131),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_153),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_94),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_143),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_31),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_117),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_101),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_130),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_59),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_72),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_123),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_128),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_105),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_39),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_55),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_109),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_154),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_134),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_96),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_107),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_25),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_4),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_126),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_58),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_106),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_54),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_4),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_135),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_102),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_53),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_71),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_36),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_47),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_50),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_33),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_64),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_122),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_5),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_62),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_17),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_43),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_44),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_164),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_147),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_56),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_6),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_57),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_55),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_136),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_33),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_114),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_119),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_179),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_3),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_9),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_12),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_90),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_22),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_50),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_74),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_39),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_93),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_60),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_35),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_166),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_15),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_2),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_99),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_8),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_91),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_89),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_124),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_21),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_41),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_22),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_177),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_133),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_149),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_82),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_1),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_167),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_125),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_12),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_155),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_44),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_32),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_29),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_67),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_38),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_98),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_23),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_24),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_181),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_169),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_113),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_110),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_27),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_54),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_11),
.Y(n_317)
);

BUFx4f_ASAP7_75t_SL g318 ( 
.A(n_56),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_25),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_27),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_180),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_46),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_129),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_32),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_150),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_172),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_61),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_86),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_3),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_21),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_57),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_8),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_40),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_178),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_139),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_61),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_42),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_84),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_112),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_11),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_24),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_38),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_111),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_176),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_5),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_0),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_62),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_116),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_26),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_29),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_78),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_28),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_81),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_9),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_157),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_137),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_69),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_46),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_14),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_250),
.B(n_0),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_183),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_185),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_233),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_289),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_183),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_186),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_7),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_209),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_234),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_188),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_189),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_186),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_193),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_218),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_193),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_190),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_314),
.Y(n_377)
);

BUFx6f_ASAP7_75t_SL g378 ( 
.A(n_232),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_199),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_199),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_191),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_321),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_218),
.B(n_10),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_196),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_333),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_344),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_195),
.B(n_10),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_184),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_197),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_201),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_220),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_227),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_229),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_236),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_237),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_211),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_211),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_211),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_240),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_232),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_243),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_201),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_244),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_251),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_205),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_205),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_252),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_207),
.B(n_13),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_255),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_195),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_210),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_256),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_258),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_200),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_210),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_192),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_215),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_207),
.B(n_13),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_259),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_268),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_213),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_213),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_274),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_216),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_276),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_200),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_216),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_224),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_198),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_266),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_279),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_204),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_206),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_224),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_202),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_194),
.B(n_15),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_230),
.B(n_16),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_208),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_232),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_215),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_282),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_202),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_228),
.B(n_16),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_230),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_284),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_235),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_212),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_285),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_235),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_431),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_431),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_308),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_401),
.B(n_266),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_385),
.B(n_266),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_265),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_362),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_361),
.A2(n_242),
.B(n_239),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_418),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_365),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_368),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_366),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_372),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_450),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_375),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_388),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_379),
.Y(n_471)
);

AND2x6_ASAP7_75t_L g472 ( 
.A(n_409),
.B(n_194),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_380),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_419),
.B(n_266),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_403),
.B(n_266),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_362),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_417),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_430),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_406),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_433),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_407),
.B(n_272),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_412),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_434),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_416),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_439),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_448),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

BUFx8_ASAP7_75t_L g489 ( 
.A(n_378),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_423),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_425),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_383),
.B(n_194),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_428),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_435),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_441),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_445),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_R g498 ( 
.A(n_386),
.B(n_214),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_440),
.B(n_272),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_272),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_441),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_387),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_370),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_387),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_R g505 ( 
.A(n_370),
.B(n_217),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_444),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_369),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_367),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_444),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_438),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_411),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_415),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_371),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_363),
.B(n_308),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_364),
.B(n_296),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_360),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_371),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_374),
.B(n_272),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_436),
.B(n_265),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_376),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_449),
.B(n_296),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_376),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_408),
.B(n_231),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_505),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_381),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_468),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_516),
.B(n_426),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_381),
.Y(n_531)
);

BUFx4f_ASAP7_75t_L g532 ( 
.A(n_460),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_472),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_501),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_468),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_397),
.Y(n_536)
);

NOR3xp33_ASAP7_75t_L g537 ( 
.A(n_525),
.B(n_399),
.C(n_398),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_489),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_501),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_468),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_461),
.B(n_389),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_501),
.B(n_239),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_451),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_455),
.B(n_242),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_502),
.B(n_389),
.Y(n_545)
);

AO22x2_ASAP7_75t_L g546 ( 
.A1(n_510),
.A2(n_182),
.B1(n_358),
.B2(n_228),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_457),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_455),
.B(n_248),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_498),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_503),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_468),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_452),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_462),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_462),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_508),
.B(n_391),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_496),
.B(n_391),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_453),
.B(n_248),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_453),
.B(n_392),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_182),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_520),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_453),
.B(n_392),
.Y(n_562)
);

NAND2x1p5_ASAP7_75t_L g563 ( 
.A(n_521),
.B(n_261),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_457),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_508),
.B(n_393),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_465),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_466),
.Y(n_567)
);

OR2x2_ASAP7_75t_SL g568 ( 
.A(n_458),
.B(n_249),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_464),
.B(n_393),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_521),
.B(n_338),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_453),
.B(n_338),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_466),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_520),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_474),
.B(n_395),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_468),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_467),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_480),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_467),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_502),
.B(n_356),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_465),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_510),
.A2(n_384),
.B1(n_446),
.B2(n_442),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_470),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_460),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_469),
.Y(n_585)
);

BUFx8_ASAP7_75t_SL g586 ( 
.A(n_463),
.Y(n_586)
);

INVxp33_ASAP7_75t_L g587 ( 
.A(n_502),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_504),
.B(n_395),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_469),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_473),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_454),
.B(n_396),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_480),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_473),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_480),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_480),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_475),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_521),
.B(n_356),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_475),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_515),
.B(n_519),
.C(n_512),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_474),
.B(n_396),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_491),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_522),
.B(n_402),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_499),
.A2(n_413),
.B1(n_446),
.B2(n_442),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_460),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_504),
.B(n_402),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_491),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_504),
.B(n_267),
.Y(n_607)
);

BUFx4f_ASAP7_75t_L g608 ( 
.A(n_460),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_465),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_483),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_521),
.B(n_249),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_493),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_480),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_510),
.B(n_404),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_521),
.B(n_264),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_506),
.B(n_404),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_507),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_493),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_492),
.A2(n_272),
.B1(n_303),
.B2(n_262),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_495),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_506),
.B(n_405),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_480),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_506),
.B(n_405),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_495),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_509),
.B(n_410),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_472),
.B(n_410),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_509),
.B(n_413),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_509),
.B(n_414),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_519),
.B(n_414),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_483),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_483),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_514),
.B(n_420),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_471),
.B(n_420),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_497),
.B(n_267),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_492),
.B(n_328),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_472),
.B(n_421),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_497),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_471),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_471),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_471),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_492),
.A2(n_303),
.B1(n_262),
.B2(n_358),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_485),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_472),
.B(n_421),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_488),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_485),
.B(n_424),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_485),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_485),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_511),
.B(n_283),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_492),
.A2(n_303),
.B1(n_264),
.B2(n_273),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_485),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_511),
.B(n_278),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_512),
.B(n_424),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_517),
.B(n_432),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_517),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_524),
.B(n_449),
.C(n_432),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_488),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_488),
.Y(n_658)
);

INVxp67_ASAP7_75t_SL g659 ( 
.A(n_476),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_472),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_490),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_492),
.A2(n_303),
.B1(n_315),
.B2(n_281),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_490),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_490),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_524),
.B(n_278),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_477),
.B(n_273),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_478),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_492),
.A2(n_472),
.B1(n_518),
.B2(n_513),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_494),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_494),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_494),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_479),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_492),
.B(n_328),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_SL g674 ( 
.A1(n_523),
.A2(n_247),
.B1(n_257),
.B2(n_277),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_527),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_584),
.A2(n_492),
.B1(n_472),
.B2(n_335),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_587),
.B(n_456),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_659),
.B(n_472),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_575),
.B(n_456),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_630),
.A2(n_377),
.B1(n_382),
.B2(n_187),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_561),
.B(n_481),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_587),
.B(n_484),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_574),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_527),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_633),
.B(n_602),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_545),
.B(n_486),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_584),
.A2(n_302),
.B1(n_323),
.B2(n_343),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_543),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_548),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_545),
.B(n_487),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_532),
.A2(n_482),
.B(n_476),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_548),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_600),
.B(n_459),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_626),
.B(n_489),
.C(n_292),
.Y(n_694)
);

INVxp33_ASAP7_75t_L g695 ( 
.A(n_588),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_614),
.B(n_378),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_531),
.A2(n_335),
.B1(n_302),
.B2(n_357),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_630),
.B(n_459),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_530),
.B(n_378),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_564),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_569),
.B(n_489),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_544),
.B(n_295),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_543),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_616),
.B(n_203),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_536),
.B(n_591),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_538),
.B(n_295),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_564),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_547),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_554),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_547),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_544),
.B(n_297),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_544),
.B(n_297),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_555),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_567),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_549),
.B(n_482),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_549),
.B(n_323),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_528),
.A2(n_271),
.B1(n_219),
.B2(n_221),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_549),
.B(n_343),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_619),
.B(n_348),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_541),
.B(n_489),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_572),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_533),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_577),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_558),
.B(n_348),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_533),
.B(n_328),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_553),
.Y(n_726)
);

O2A1O1Ixp5_ASAP7_75t_L g727 ( 
.A1(n_532),
.A2(n_500),
.B(n_357),
.C(n_355),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_604),
.A2(n_355),
.B1(n_303),
.B2(n_222),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_656),
.B(n_603),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_553),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_668),
.A2(n_269),
.B1(n_353),
.B2(n_351),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_579),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_655),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_616),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_585),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_566),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_557),
.B(n_582),
.Y(n_737)
);

NOR3xp33_ASAP7_75t_L g738 ( 
.A(n_674),
.B(n_263),
.C(n_301),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_586),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_558),
.B(n_500),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_533),
.B(n_660),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_566),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_558),
.B(n_223),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_589),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_623),
.B(n_318),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_642),
.B(n_225),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_533),
.B(n_328),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_650),
.B(n_226),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_588),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_623),
.B(n_305),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_533),
.B(n_328),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_590),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_593),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_655),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_596),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_662),
.B(n_238),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_532),
.A2(n_281),
.B(n_287),
.C(n_352),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_528),
.B(n_241),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_628),
.B(n_350),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_611),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_653),
.B(n_605),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_581),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_598),
.B(n_245),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_604),
.A2(n_328),
.B1(n_287),
.B2(n_352),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_550),
.B(n_320),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_601),
.B(n_246),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_606),
.B(n_253),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_581),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_605),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_653),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_636),
.A2(n_328),
.B1(n_317),
.B2(n_322),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_612),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_538),
.B(n_315),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_660),
.B(n_608),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_618),
.B(n_254),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_609),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_628),
.B(n_291),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_660),
.B(n_328),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_634),
.A2(n_260),
.B1(n_270),
.B2(n_275),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_608),
.B(n_280),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_636),
.A2(n_324),
.B1(n_317),
.B2(n_322),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_608),
.A2(n_324),
.B(n_346),
.C(n_349),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_620),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_627),
.B(n_286),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_609),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_624),
.B(n_288),
.Y(n_786)
);

OAI221xp5_ASAP7_75t_L g787 ( 
.A1(n_599),
.A2(n_346),
.B1(n_354),
.B2(n_347),
.C(n_359),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_526),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_638),
.B(n_290),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_563),
.B(n_639),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_534),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_634),
.A2(n_621),
.B1(n_562),
.B2(n_559),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_637),
.B(n_294),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_537),
.B(n_345),
.C(n_342),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_610),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_586),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_539),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_542),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_629),
.A2(n_299),
.B1(n_300),
.B2(n_339),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_644),
.B(n_306),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_563),
.B(n_311),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_640),
.B(n_312),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_610),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_673),
.A2(n_341),
.B1(n_340),
.B2(n_337),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_641),
.B(n_649),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_556),
.B(n_293),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_607),
.B(n_570),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_611),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_611),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_607),
.B(n_313),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_629),
.B(n_298),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_649),
.B(n_325),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_607),
.B(n_326),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_570),
.B(n_334),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_542),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_654),
.B(n_336),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_542),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_597),
.B(n_332),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_556),
.B(n_331),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_597),
.B(n_652),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_565),
.B(n_330),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_635),
.B(n_83),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_652),
.B(n_329),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_654),
.B(n_327),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_652),
.B(n_319),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_631),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_652),
.B(n_316),
.Y(n_827)
);

INVx8_ASAP7_75t_L g828 ( 
.A(n_560),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_652),
.B(n_310),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_632),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_652),
.B(n_309),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_568),
.B(n_307),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_632),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_565),
.B(n_304),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_611),
.B(n_76),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_551),
.B(n_17),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_645),
.B(n_77),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_538),
.B(n_73),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_645),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_646),
.B(n_18),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_673),
.A2(n_19),
.B(n_20),
.C(n_23),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_663),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_676),
.A2(n_535),
.B(n_540),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_685),
.A2(n_646),
.B1(n_560),
.B2(n_571),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_741),
.A2(n_535),
.B(n_540),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_741),
.A2(n_678),
.B(n_722),
.Y(n_846)
);

AO21x1_ASAP7_75t_L g847 ( 
.A1(n_840),
.A2(n_648),
.B(n_635),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_705),
.B(n_615),
.Y(n_848)
);

INVx11_ASAP7_75t_L g849 ( 
.A(n_788),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_691),
.A2(n_592),
.B(n_552),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_727),
.A2(n_571),
.B(n_615),
.Y(n_851)
);

AO21x1_ASAP7_75t_L g852 ( 
.A1(n_780),
.A2(n_665),
.B(n_670),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_722),
.A2(n_535),
.B(n_540),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_722),
.A2(n_625),
.B(n_573),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_798),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_677),
.B(n_615),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_778),
.A2(n_571),
.B(n_615),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_774),
.A2(n_625),
.B(n_573),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_774),
.A2(n_573),
.B(n_595),
.Y(n_859)
);

AO21x2_ASAP7_75t_L g860 ( 
.A1(n_780),
.A2(n_665),
.B(n_661),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_L g861 ( 
.A1(n_778),
.A2(n_820),
.B(n_807),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_687),
.A2(n_580),
.B1(n_546),
.B2(n_571),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_761),
.B(n_551),
.Y(n_863)
);

AO32x1_ASAP7_75t_L g864 ( 
.A1(n_731),
.A2(n_791),
.A3(n_797),
.B1(n_708),
.B2(n_710),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_677),
.B(n_560),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_740),
.A2(n_790),
.B(n_715),
.Y(n_866)
);

AO21x2_ASAP7_75t_L g867 ( 
.A1(n_784),
.A2(n_664),
.B(n_658),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_683),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_715),
.A2(n_595),
.B(n_573),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_SL g870 ( 
.A1(n_757),
.A2(n_657),
.B(n_669),
.C(n_663),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_782),
.A2(n_560),
.B(n_671),
.C(n_666),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_698),
.A2(n_595),
.B(n_622),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_679),
.A2(n_595),
.B(n_622),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_693),
.B(n_580),
.Y(n_874)
);

AO21x1_ASAP7_75t_L g875 ( 
.A1(n_737),
.A2(n_671),
.B(n_546),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_707),
.B(n_551),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_784),
.A2(n_622),
.B(n_529),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_750),
.A2(n_594),
.B(n_552),
.C(n_576),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_733),
.B(n_666),
.Y(n_879)
);

AOI21x1_ASAP7_75t_L g880 ( 
.A1(n_793),
.A2(n_666),
.B(n_546),
.Y(n_880)
);

NAND2x1p5_ASAP7_75t_L g881 ( 
.A(n_822),
.B(n_529),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_792),
.B(n_580),
.Y(n_882)
);

BUFx12f_ASAP7_75t_L g883 ( 
.A(n_739),
.Y(n_883)
);

AOI21x1_ASAP7_75t_L g884 ( 
.A1(n_793),
.A2(n_666),
.B(n_571),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_800),
.A2(n_622),
.B(n_529),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_758),
.B(n_580),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_800),
.A2(n_594),
.B(n_576),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_782),
.A2(n_552),
.B(n_651),
.C(n_576),
.Y(n_888)
);

OA22x2_ASAP7_75t_L g889 ( 
.A1(n_770),
.A2(n_672),
.B1(n_667),
.B2(n_583),
.Y(n_889)
);

AOI21x1_ASAP7_75t_L g890 ( 
.A1(n_725),
.A2(n_571),
.B(n_651),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_689),
.B(n_580),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_689),
.B(n_580),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_817),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_707),
.B(n_672),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_675),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_L g896 ( 
.A(n_760),
.B(n_667),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_692),
.B(n_651),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_805),
.A2(n_647),
.B(n_643),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_695),
.B(n_617),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_733),
.B(n_617),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_805),
.A2(n_647),
.B(n_643),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_749),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_695),
.B(n_647),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_757),
.A2(n_643),
.B(n_613),
.C(n_594),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_802),
.A2(n_613),
.B(n_592),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_725),
.A2(n_613),
.B(n_592),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_675),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_747),
.A2(n_578),
.B(n_80),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_760),
.A2(n_578),
.B1(n_87),
.B2(n_88),
.Y(n_909)
);

BUFx12f_ASAP7_75t_L g910 ( 
.A(n_739),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_754),
.B(n_578),
.Y(n_911)
);

AOI21x1_ASAP7_75t_L g912 ( 
.A1(n_747),
.A2(n_68),
.B(n_170),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_682),
.B(n_19),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_SL g914 ( 
.A(n_765),
.B(n_79),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_707),
.B(n_66),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_751),
.A2(n_95),
.B(n_168),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_777),
.A2(n_811),
.B(n_816),
.C(n_824),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_751),
.A2(n_174),
.B(n_160),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_808),
.A2(n_158),
.B(n_156),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_808),
.A2(n_152),
.B(n_148),
.Y(n_920)
);

AO22x1_ASAP7_75t_L g921 ( 
.A1(n_738),
.A2(n_20),
.B1(n_26),
.B2(n_28),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_692),
.B(n_30),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_769),
.B(n_30),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_809),
.A2(n_146),
.B(n_121),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_764),
.A2(n_728),
.B(n_771),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_815),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_700),
.B(n_34),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_700),
.B(n_34),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_809),
.A2(n_120),
.B(n_115),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_702),
.A2(n_108),
.B(n_104),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_729),
.A2(n_103),
.B1(n_100),
.B2(n_97),
.Y(n_931)
);

OAI22xp33_ASAP7_75t_L g932 ( 
.A1(n_759),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_932)
);

NOR2x1_ASAP7_75t_L g933 ( 
.A(n_694),
.B(n_43),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_681),
.B(n_45),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_734),
.B(n_59),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_684),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_711),
.A2(n_45),
.B(n_48),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_781),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_810),
.A2(n_813),
.B(n_815),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_684),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_788),
.Y(n_941)
);

AOI21xp33_ASAP7_75t_L g942 ( 
.A1(n_834),
.A2(n_53),
.B(n_745),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_688),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_709),
.B(n_713),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_822),
.A2(n_814),
.B(n_724),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_686),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_822),
.B(n_707),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_714),
.B(n_721),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_690),
.B(n_704),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_746),
.A2(n_743),
.B(n_716),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_723),
.B(n_732),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_795),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_841),
.A2(n_712),
.B(n_718),
.C(n_719),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_754),
.B(n_735),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_744),
.B(n_752),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_753),
.B(n_755),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_787),
.A2(n_696),
.B(n_699),
.C(n_783),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_806),
.B(n_819),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_717),
.B(n_720),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_819),
.B(n_821),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_772),
.B(n_730),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_818),
.A2(n_701),
.B(n_812),
.C(n_801),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_680),
.B(n_786),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_748),
.A2(n_756),
.B(n_789),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_773),
.B(n_838),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_688),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_763),
.A2(n_767),
.B(n_766),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_703),
.B(n_730),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_775),
.B(n_779),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_703),
.B(n_726),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_708),
.B(n_726),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_710),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_799),
.B(n_812),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_736),
.B(n_776),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_736),
.A2(n_768),
.B(n_785),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_801),
.A2(n_835),
.B(n_825),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_697),
.A2(n_803),
.B1(n_785),
.B2(n_742),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_795),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_826),
.A2(n_842),
.B(n_839),
.Y(n_979)
);

AO21x1_ASAP7_75t_L g980 ( 
.A1(n_837),
.A2(n_827),
.B(n_823),
.Y(n_980)
);

O2A1O1Ixp5_ASAP7_75t_L g981 ( 
.A1(n_742),
.A2(n_776),
.B(n_803),
.C(n_762),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_829),
.A2(n_831),
.B(n_830),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_762),
.B(n_768),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_838),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_795),
.B(n_833),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_828),
.A2(n_838),
.B1(n_821),
.B2(n_706),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_794),
.A2(n_828),
.B1(n_838),
.B2(n_836),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_837),
.A2(n_832),
.B(n_706),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_828),
.A2(n_706),
.B(n_773),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_804),
.B(n_828),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_841),
.B(n_706),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_773),
.A2(n_840),
.B(n_780),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_796),
.A2(n_533),
.B(n_660),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_685),
.A2(n_737),
.B1(n_705),
.B2(n_792),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_691),
.A2(n_608),
.B(n_532),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_815),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_676),
.A2(n_533),
.B(n_660),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_685),
.B(n_705),
.Y(n_998)
);

NOR2xp67_ASAP7_75t_L g999 ( 
.A(n_694),
.B(n_656),
.Y(n_999)
);

INVx5_ASAP7_75t_L g1000 ( 
.A(n_722),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_685),
.A2(n_750),
.B(n_840),
.C(n_737),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_683),
.Y(n_1002)
);

O2A1O1Ixp5_ASAP7_75t_L g1003 ( 
.A1(n_727),
.A2(n_570),
.B(n_597),
.C(n_691),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_676),
.A2(n_533),
.B(n_660),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_778),
.A2(n_793),
.B(n_784),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_L g1006 ( 
.A(n_685),
.B(n_750),
.C(n_816),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_683),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_798),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_685),
.A2(n_750),
.B(n_840),
.C(n_737),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_782),
.A2(n_757),
.B(n_841),
.C(n_711),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_685),
.B(n_705),
.Y(n_1011)
);

OA22x2_ASAP7_75t_L g1012 ( 
.A1(n_761),
.A2(n_770),
.B1(n_749),
.B2(n_769),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_685),
.B(n_705),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_675),
.Y(n_1014)
);

NOR2xp67_ASAP7_75t_SL g1015 ( 
.A(n_760),
.B(n_533),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_676),
.A2(n_533),
.B(n_660),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_782),
.A2(n_757),
.B(n_841),
.C(n_711),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_685),
.B(n_705),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_675),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_676),
.A2(n_533),
.B(n_660),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_685),
.A2(n_750),
.B(n_840),
.C(n_737),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_815),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_676),
.A2(n_533),
.B(n_660),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_676),
.A2(n_685),
.B1(n_668),
.B2(n_792),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_695),
.B(n_685),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_798),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_676),
.A2(n_685),
.B1(n_668),
.B2(n_792),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_685),
.B(n_705),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_798),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_695),
.B(n_685),
.Y(n_1030)
);

NOR2xp67_ASAP7_75t_L g1031 ( 
.A(n_694),
.B(n_656),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1018),
.B(n_1028),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_954),
.B(n_879),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_L g1036 ( 
.A1(n_917),
.A2(n_1021),
.B(n_1009),
.C(n_1001),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_994),
.A2(n_1006),
.B1(n_1024),
.B2(n_1027),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1025),
.B(n_1030),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_981),
.A2(n_859),
.B(n_858),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_998),
.B(n_1025),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_SL g1041 ( 
.A1(n_995),
.A2(n_857),
.B(n_947),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_961),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_1000),
.A2(n_1004),
.B(n_997),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_SL g1044 ( 
.A1(n_947),
.A2(n_965),
.B(n_851),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_913),
.A2(n_942),
.B(n_925),
.C(n_1030),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_887),
.A2(n_905),
.B(n_885),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_1000),
.A2(n_1020),
.B(n_1016),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_949),
.B(n_963),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_877),
.A2(n_982),
.B(n_901),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_849),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_898),
.A2(n_979),
.B(n_890),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_975),
.A2(n_872),
.B(n_845),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_861),
.A2(n_866),
.B(n_1003),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_855),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_911),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_958),
.B(n_856),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1000),
.A2(n_1023),
.B(n_945),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1014),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1000),
.A2(n_843),
.B(n_967),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_893),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_869),
.A2(n_1005),
.B(n_906),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1008),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_853),
.A2(n_1003),
.B(n_904),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_976),
.A2(n_886),
.B(n_884),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_954),
.B(n_879),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_904),
.A2(n_854),
.B(n_873),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_847),
.A2(n_852),
.A3(n_992),
.B(n_875),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_950),
.A2(n_939),
.B(n_970),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_968),
.A2(n_971),
.B(n_964),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_969),
.A2(n_882),
.B(n_874),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_941),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_952),
.A2(n_973),
.B(n_953),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_946),
.B(n_868),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_984),
.B(n_965),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_1002),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_848),
.B(n_960),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_938),
.A2(n_984),
.B1(n_862),
.B2(n_844),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_980),
.A2(n_878),
.A3(n_962),
.B(n_991),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_1002),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_952),
.A2(n_953),
.B(n_865),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_984),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1026),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_974),
.A2(n_983),
.B(n_888),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_957),
.A2(n_909),
.A3(n_903),
.B(n_864),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_891),
.A2(n_892),
.B(n_881),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_934),
.A2(n_871),
.B(n_959),
.C(n_1017),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_944),
.B(n_948),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1010),
.A2(n_1017),
.B(n_888),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_984),
.B(n_926),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_999),
.A2(n_1031),
.B1(n_986),
.B2(n_899),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_SL g1091 ( 
.A1(n_937),
.A2(n_932),
.B1(n_1010),
.B2(n_938),
.C(n_871),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_903),
.B(n_1029),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_895),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_881),
.A2(n_897),
.B(n_990),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_911),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_977),
.A2(n_870),
.B(n_936),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_926),
.B(n_1022),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_900),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_985),
.A2(n_956),
.B(n_951),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_L g1100 ( 
.A1(n_988),
.A2(n_1015),
.B(n_880),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_955),
.A2(n_993),
.B(n_860),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_977),
.A2(n_940),
.B(n_907),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_862),
.A2(n_1012),
.B1(n_987),
.B2(n_932),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_996),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_943),
.B(n_972),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_860),
.A2(n_867),
.B(n_930),
.Y(n_1106)
);

AO21x1_ASAP7_75t_L g1107 ( 
.A1(n_931),
.A2(n_927),
.B(n_922),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_902),
.B(n_1007),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_864),
.A2(n_928),
.A3(n_966),
.B(n_1019),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_867),
.A2(n_978),
.B(n_989),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_978),
.A2(n_915),
.B(n_908),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_902),
.B(n_923),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_SL g1113 ( 
.A(n_876),
.B(n_894),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_883),
.B(n_910),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_914),
.A2(n_933),
.B(n_896),
.C(n_929),
.Y(n_1115)
);

AOI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_889),
.A2(n_863),
.B(n_935),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_919),
.A2(n_920),
.B(n_924),
.C(n_918),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_912),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_900),
.B(n_889),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_921),
.B(n_916),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1025),
.B(n_761),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1014),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1124)
);

AO21x2_ASAP7_75t_L g1125 ( 
.A1(n_917),
.A2(n_992),
.B(n_847),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1126)
);

OAI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1011),
.A2(n_1018),
.B1(n_1028),
.B2(n_1013),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1001),
.A2(n_1021),
.B(n_1009),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_917),
.A2(n_1009),
.B(n_1021),
.C(n_1001),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_947),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_847),
.A2(n_852),
.A3(n_992),
.B(n_875),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_954),
.B(n_879),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_L g1141 ( 
.A1(n_917),
.A2(n_1009),
.B(n_1021),
.C(n_1001),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_917),
.A2(n_1009),
.B(n_1021),
.C(n_1001),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1006),
.B(n_917),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_941),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_984),
.Y(n_1150)
);

AO21x1_ASAP7_75t_L g1151 ( 
.A1(n_1024),
.A2(n_1027),
.B(n_994),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1006),
.B(n_917),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1025),
.B(n_761),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_868),
.Y(n_1154)
);

OA22x2_ASAP7_75t_L g1155 ( 
.A1(n_994),
.A2(n_1011),
.B1(n_1018),
.B2(n_1013),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_1003),
.A2(n_995),
.B(n_882),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_994),
.A2(n_1001),
.B1(n_1021),
.B2(n_1009),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_868),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1025),
.B(n_761),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_984),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_847),
.A2(n_852),
.A3(n_992),
.B(n_875),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_850),
.A2(n_846),
.B(n_981),
.Y(n_1168)
);

AO21x1_ASAP7_75t_L g1169 ( 
.A1(n_1024),
.A2(n_1027),
.B(n_994),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1170)
);

O2A1O1Ixp5_ASAP7_75t_L g1171 ( 
.A1(n_917),
.A2(n_1009),
.B(n_1021),
.C(n_1001),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_917),
.A2(n_1009),
.B(n_1021),
.C(n_1001),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1173)
);

INVx6_ASAP7_75t_L g1174 ( 
.A(n_900),
.Y(n_1174)
);

OAI222xp33_ASAP7_75t_L g1175 ( 
.A1(n_994),
.A2(n_1013),
.B1(n_1018),
.B2(n_1028),
.C1(n_1011),
.C2(n_932),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_L g1176 ( 
.A(n_1006),
.B(n_917),
.C(n_1001),
.Y(n_1176)
);

AOI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1005),
.A2(n_780),
.B(n_979),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_SL g1181 ( 
.A1(n_875),
.A2(n_880),
.B(n_937),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1006),
.B(n_917),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1006),
.B(n_917),
.C(n_685),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_1000),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_847),
.A2(n_852),
.A3(n_992),
.B(n_875),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1000),
.A2(n_660),
.B(n_533),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_984),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1038),
.B(n_1034),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1175),
.B(n_1128),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1121),
.B(n_1153),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1059),
.A2(n_1057),
.B(n_1041),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1184),
.A2(n_1037),
.B(n_1072),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_1184),
.Y(n_1194)
);

CKINVDCx16_ASAP7_75t_R g1195 ( 
.A(n_1071),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1054),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1164),
.B(n_1112),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1060),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1149),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1127),
.B(n_1038),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1032),
.B(n_1170),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1154),
.Y(n_1202)
);

BUFx2_ASAP7_75t_SL g1203 ( 
.A(n_1050),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1184),
.A2(n_1037),
.B(n_1106),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1081),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1058),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1062),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1082),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1184),
.A2(n_1053),
.B(n_1133),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1048),
.A2(n_1183),
.B1(n_1090),
.B2(n_1151),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1108),
.B(n_1126),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1035),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_1081),
.B(n_1150),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1122),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1053),
.A2(n_1172),
.B(n_1142),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1169),
.A2(n_1160),
.B1(n_1130),
.B2(n_1176),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1113),
.A2(n_1137),
.B1(n_1145),
.B2(n_1126),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1131),
.A2(n_1145),
.B1(n_1162),
.B2(n_1137),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1099),
.A2(n_1152),
.B(n_1146),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1105),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1035),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1131),
.A2(n_1157),
.B1(n_1158),
.B2(n_1178),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1157),
.A2(n_1162),
.B1(n_1173),
.B2(n_1158),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1173),
.B(n_1178),
.Y(n_1224)
);

NOR2xp67_ASAP7_75t_L g1225 ( 
.A(n_1050),
.B(n_1073),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1114),
.B(n_1075),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1081),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1081),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1042),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1040),
.B(n_1087),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1045),
.A2(n_1077),
.B1(n_1086),
.B2(n_1074),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1098),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1036),
.A2(n_1171),
.B(n_1141),
.C(n_1091),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1076),
.B(n_1056),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1092),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1075),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1056),
.B(n_1092),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1155),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1083),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1074),
.B(n_1044),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1182),
.A2(n_1101),
.B(n_1047),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1065),
.B(n_1140),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1065),
.B(n_1140),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1160),
.B(n_1155),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1161),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1091),
.A2(n_1077),
.B(n_1130),
.C(n_1088),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1079),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1079),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1055),
.B(n_1095),
.Y(n_1249)
);

AOI21xp33_ASAP7_75t_L g1250 ( 
.A1(n_1120),
.A2(n_1103),
.B(n_1125),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1097),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1043),
.A2(n_1070),
.B(n_1117),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1088),
.A2(n_1080),
.B(n_1102),
.C(n_1096),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1055),
.B(n_1095),
.Y(n_1254)
);

AO22x1_ASAP7_75t_L g1255 ( 
.A1(n_1150),
.A2(n_1188),
.B1(n_1166),
.B2(n_1120),
.Y(n_1255)
);

AND2x6_ASAP7_75t_L g1256 ( 
.A(n_1150),
.B(n_1166),
.Y(n_1256)
);

AO21x2_ASAP7_75t_L g1257 ( 
.A1(n_1181),
.A2(n_1064),
.B(n_1110),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1097),
.B(n_1116),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1166),
.A2(n_1188),
.B1(n_1089),
.B2(n_1115),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1174),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1109),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1188),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1174),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1104),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1116),
.B(n_1119),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1104),
.Y(n_1266)
);

NAND2xp33_ASAP7_75t_L g1267 ( 
.A(n_1135),
.B(n_1187),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1063),
.A2(n_1033),
.B(n_1148),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1069),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1125),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1094),
.B(n_1111),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1156),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1107),
.A2(n_1156),
.B1(n_1085),
.B2(n_1118),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1067),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1100),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1066),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1078),
.B(n_1139),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1118),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1067),
.B(n_1185),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1068),
.B(n_1061),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1052),
.A2(n_1039),
.B(n_1168),
.C(n_1165),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1132),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1138),
.A2(n_1143),
.B1(n_1180),
.B2(n_1179),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1067),
.Y(n_1284)
);

AO21x2_ASAP7_75t_L g1285 ( 
.A1(n_1123),
.A2(n_1129),
.B(n_1163),
.Y(n_1285)
);

OAI31xp33_ASAP7_75t_L g1286 ( 
.A1(n_1144),
.A2(n_1186),
.A3(n_1159),
.B(n_1084),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1167),
.B(n_1185),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1177),
.A2(n_1167),
.B1(n_1084),
.B2(n_1124),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1049),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1046),
.B(n_1134),
.Y(n_1290)
);

INVx5_ASAP7_75t_L g1291 ( 
.A(n_1136),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1147),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1054),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1128),
.B(n_1011),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1093),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1081),
.B(n_1184),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1151),
.A2(n_1169),
.B1(n_1037),
.B2(n_1006),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1081),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1175),
.A2(n_1009),
.B(n_1021),
.C(n_1001),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1074),
.B(n_1044),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1121),
.B(n_1153),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1071),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1071),
.Y(n_1303)
);

NAND2xp33_ASAP7_75t_L g1304 ( 
.A(n_1077),
.B(n_917),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1053),
.A2(n_1130),
.B(n_1063),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1051),
.A2(n_850),
.B(n_1033),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1128),
.B(n_1011),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1059),
.A2(n_660),
.B(n_533),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1054),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1093),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1093),
.Y(n_1311)
);

INVx5_ASAP7_75t_L g1312 ( 
.A(n_1184),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1081),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1175),
.A2(n_1009),
.B(n_1021),
.C(n_1001),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1128),
.A2(n_1009),
.B(n_1021),
.C(n_1001),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1054),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1071),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1054),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_SL g1319 ( 
.A(n_1050),
.B(n_583),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1050),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1128),
.A2(n_1006),
.B1(n_1009),
.B2(n_1001),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1128),
.A2(n_1006),
.B1(n_1009),
.B2(n_1001),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1071),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1059),
.A2(n_660),
.B(n_533),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1154),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1128),
.B(n_1011),
.Y(n_1326)
);

NAND2xp33_ASAP7_75t_L g1327 ( 
.A(n_1077),
.B(n_917),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1128),
.B(n_1011),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1038),
.B(n_1034),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1093),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1035),
.B(n_1065),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1054),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1054),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1059),
.A2(n_660),
.B(n_533),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1121),
.B(n_1153),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1071),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1081),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1241),
.A2(n_1281),
.B(n_1250),
.Y(n_1338)
);

INVx4_ASAP7_75t_L g1339 ( 
.A(n_1194),
.Y(n_1339)
);

BUFx4f_ASAP7_75t_SL g1340 ( 
.A(n_1303),
.Y(n_1340)
);

BUFx10_ASAP7_75t_L g1341 ( 
.A(n_1302),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1190),
.A2(n_1327),
.B1(n_1304),
.B2(n_1200),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1236),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1303),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1196),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1198),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1190),
.A2(n_1327),
.B1(n_1304),
.B2(n_1200),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1217),
.B(n_1238),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1194),
.Y(n_1349)
);

OAI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1294),
.A2(n_1326),
.B1(n_1328),
.B2(n_1307),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1210),
.A2(n_1222),
.B1(n_1223),
.B2(n_1218),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1201),
.A2(n_1224),
.B1(n_1189),
.B2(n_1329),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1231),
.A2(n_1322),
.B1(n_1321),
.B2(n_1265),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1234),
.B(n_1191),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1207),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1208),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1202),
.Y(n_1357)
);

INVx8_ASAP7_75t_L g1358 ( 
.A(n_1256),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1306),
.A2(n_1192),
.B(n_1252),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1283),
.A2(n_1280),
.B(n_1290),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1325),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1293),
.Y(n_1362)
);

AO21x1_ASAP7_75t_L g1363 ( 
.A1(n_1299),
.A2(n_1314),
.B(n_1219),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1301),
.B(n_1335),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1297),
.A2(n_1216),
.B(n_1246),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1309),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1316),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1315),
.A2(n_1193),
.B(n_1215),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1194),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1318),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1226),
.A2(n_1230),
.B1(n_1284),
.B2(n_1263),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1266),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1320),
.Y(n_1373)
);

BUFx12f_ASAP7_75t_L g1374 ( 
.A(n_1320),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1284),
.A2(n_1263),
.B1(n_1244),
.B2(n_1319),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1332),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1333),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1295),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1274),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1312),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1199),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1235),
.B(n_1220),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1211),
.B(n_1237),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1232),
.A2(n_1197),
.B1(n_1258),
.B2(n_1225),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1310),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1311),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1212),
.A2(n_1221),
.B1(n_1243),
.B2(n_1331),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1281),
.A2(n_1253),
.B(n_1204),
.Y(n_1388)
);

BUFx2_ASAP7_75t_R g1389 ( 
.A(n_1336),
.Y(n_1389)
);

CKINVDCx6p67_ASAP7_75t_R g1390 ( 
.A(n_1195),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1273),
.A2(n_1209),
.B(n_1253),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1330),
.Y(n_1392)
);

BUFx2_ASAP7_75t_R g1393 ( 
.A(n_1199),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1247),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1266),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1248),
.Y(n_1396)
);

NAND2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1312),
.B(n_1278),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1296),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1229),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1206),
.Y(n_1400)
);

NAND2x1p5_ASAP7_75t_L g1401 ( 
.A(n_1337),
.B(n_1272),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1279),
.B(n_1214),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1240),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1206),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1245),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1277),
.B(n_1274),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1240),
.B(n_1300),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1251),
.Y(n_1408)
);

AO21x1_ASAP7_75t_L g1409 ( 
.A1(n_1288),
.A2(n_1287),
.B(n_1271),
.Y(n_1409)
);

CKINVDCx6p67_ASAP7_75t_R g1410 ( 
.A(n_1317),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1254),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1269),
.A2(n_1239),
.B(n_1292),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1300),
.B(n_1249),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1259),
.A2(n_1260),
.B1(n_1242),
.B2(n_1203),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1317),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1296),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1257),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1276),
.A2(n_1289),
.B(n_1324),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1323),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1256),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1323),
.Y(n_1421)
);

CKINVDCx11_ASAP7_75t_R g1422 ( 
.A(n_1264),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1270),
.A2(n_1233),
.B(n_1261),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1205),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1264),
.Y(n_1425)
);

BUFx2_ASAP7_75t_R g1426 ( 
.A(n_1282),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1256),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1255),
.B(n_1275),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1262),
.A2(n_1267),
.B1(n_1227),
.B2(n_1228),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1262),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1305),
.B(n_1268),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1227),
.B(n_1228),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1213),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1267),
.A2(n_1313),
.B1(n_1298),
.B2(n_1289),
.Y(n_1434)
);

AOI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1268),
.A2(n_1308),
.B(n_1334),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1286),
.A2(n_1285),
.B(n_1291),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1298),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1291),
.A2(n_765),
.B1(n_1190),
.B2(n_1006),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1291),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1291),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1294),
.A2(n_1011),
.B1(n_1018),
.B2(n_1013),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1194),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1190),
.A2(n_1006),
.B1(n_1327),
.B2(n_1304),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1320),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1190),
.A2(n_1006),
.B1(n_1327),
.B2(n_1304),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1241),
.A2(n_1281),
.B(n_1250),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1190),
.A2(n_674),
.B1(n_1128),
.B2(n_1006),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1274),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1196),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1303),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1350),
.B(n_1352),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_SL g1452 ( 
.A(n_1374),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1407),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1407),
.B(n_1413),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1413),
.B(n_1403),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1379),
.B(n_1448),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1343),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1368),
.A2(n_1359),
.B(n_1409),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1381),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1402),
.B(n_1383),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1360),
.A2(n_1412),
.B(n_1435),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1344),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1413),
.B(n_1403),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1423),
.Y(n_1464)
);

BUFx2_ASAP7_75t_R g1465 ( 
.A(n_1444),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1423),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1394),
.Y(n_1467)
);

OR2x2_ASAP7_75t_SL g1468 ( 
.A(n_1388),
.B(n_1396),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1417),
.A2(n_1351),
.B(n_1365),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1418),
.A2(n_1363),
.B(n_1391),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1421),
.Y(n_1471)
);

BUFx4f_ASAP7_75t_SL g1472 ( 
.A(n_1374),
.Y(n_1472)
);

AO21x2_ASAP7_75t_L g1473 ( 
.A1(n_1363),
.A2(n_1391),
.B(n_1440),
.Y(n_1473)
);

BUFx8_ASAP7_75t_L g1474 ( 
.A(n_1357),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1344),
.Y(n_1475)
);

INVxp67_ASAP7_75t_L g1476 ( 
.A(n_1364),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1354),
.B(n_1364),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1349),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1383),
.B(n_1353),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1354),
.B(n_1342),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1347),
.A2(n_1391),
.B(n_1445),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1401),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1384),
.B(n_1441),
.Y(n_1483)
);

INVx4_ASAP7_75t_SL g1484 ( 
.A(n_1428),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1357),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1431),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1405),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1436),
.A2(n_1338),
.B(n_1446),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1406),
.B(n_1431),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1382),
.Y(n_1490)
);

AOI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1439),
.A2(n_1436),
.B(n_1428),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1443),
.B(n_1348),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1338),
.A2(n_1446),
.B(n_1434),
.Y(n_1493)
);

AO21x2_ASAP7_75t_L g1494 ( 
.A1(n_1429),
.A2(n_1367),
.B(n_1449),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1382),
.B(n_1411),
.Y(n_1495)
);

AO21x2_ASAP7_75t_L g1496 ( 
.A1(n_1345),
.A2(n_1362),
.B(n_1377),
.Y(n_1496)
);

NAND2x1_ASAP7_75t_L g1497 ( 
.A(n_1420),
.B(n_1339),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1378),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1385),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1447),
.B(n_1340),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1386),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1392),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1399),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1430),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1346),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1355),
.A2(n_1356),
.B(n_1376),
.Y(n_1506)
);

OR2x6_ASAP7_75t_L g1507 ( 
.A(n_1428),
.B(n_1358),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1397),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1438),
.A2(n_1375),
.B1(n_1371),
.B2(n_1414),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1366),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1388),
.B(n_1401),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1370),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1397),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1400),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1404),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1401),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1408),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1361),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1428),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1426),
.B(n_1450),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1390),
.A2(n_1450),
.B1(n_1387),
.B2(n_1430),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1474),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1489),
.B(n_1419),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1489),
.B(n_1390),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1486),
.B(n_1395),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1460),
.B(n_1437),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1460),
.B(n_1437),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1451),
.B(n_1424),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1484),
.B(n_1432),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1503),
.Y(n_1530)
);

AO21x1_ASAP7_75t_L g1531 ( 
.A1(n_1483),
.A2(n_1339),
.B(n_1442),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1507),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1486),
.B(n_1432),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1464),
.B(n_1432),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1494),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1506),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1509),
.A2(n_1373),
.B1(n_1422),
.B2(n_1372),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1496),
.B(n_1398),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1518),
.B(n_1389),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1496),
.B(n_1416),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1468),
.B(n_1425),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1511),
.Y(n_1542)
);

OAI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1481),
.A2(n_1415),
.B1(n_1444),
.B2(n_1427),
.C(n_1433),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1464),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1468),
.B(n_1456),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1466),
.B(n_1369),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1511),
.Y(n_1547)
);

OR2x2_ASAP7_75t_SL g1548 ( 
.A(n_1519),
.B(n_1398),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1473),
.B(n_1369),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1467),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1494),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1494),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1473),
.B(n_1380),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1490),
.B(n_1469),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1487),
.Y(n_1555)
);

OAI221xp5_ASAP7_75t_L g1556 ( 
.A1(n_1537),
.A2(n_1521),
.B1(n_1500),
.B2(n_1492),
.C(n_1485),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1543),
.A2(n_1492),
.B1(n_1462),
.B2(n_1393),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1543),
.A2(n_1476),
.B1(n_1477),
.B2(n_1479),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1548),
.A2(n_1479),
.B1(n_1528),
.B2(n_1480),
.Y(n_1559)
);

NOR3xp33_ASAP7_75t_L g1560 ( 
.A(n_1528),
.B(n_1475),
.C(n_1478),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1555),
.B(n_1457),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1555),
.B(n_1469),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1534),
.B(n_1491),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1524),
.B(n_1504),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1534),
.B(n_1491),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1524),
.A2(n_1504),
.B1(n_1520),
.B2(n_1453),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1534),
.B(n_1458),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1550),
.B(n_1480),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1530),
.A2(n_1495),
.B1(n_1512),
.B2(n_1510),
.C(n_1505),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1546),
.B(n_1458),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1539),
.A2(n_1454),
.B(n_1463),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1550),
.B(n_1510),
.Y(n_1572)
);

AOI211xp5_ASAP7_75t_L g1573 ( 
.A1(n_1531),
.A2(n_1415),
.B(n_1516),
.C(n_1493),
.Y(n_1573)
);

OAI221xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1541),
.A2(n_1410),
.B1(n_1482),
.B2(n_1516),
.C(n_1513),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1523),
.B(n_1512),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1523),
.B(n_1517),
.Y(n_1576)
);

NAND4xp25_ASAP7_75t_SL g1577 ( 
.A(n_1531),
.B(n_1373),
.C(n_1465),
.D(n_1517),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1542),
.B(n_1470),
.Y(n_1578)
);

OAI21xp33_ASAP7_75t_L g1579 ( 
.A1(n_1554),
.A2(n_1471),
.B(n_1459),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1522),
.A2(n_1427),
.B(n_1442),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1536),
.A2(n_1488),
.B(n_1461),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1525),
.B(n_1499),
.Y(n_1582)
);

OA211x2_ASAP7_75t_L g1583 ( 
.A1(n_1538),
.A2(n_1497),
.B(n_1484),
.C(n_1472),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1533),
.B(n_1499),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1533),
.B(n_1501),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1542),
.B(n_1455),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1535),
.B(n_1552),
.C(n_1551),
.Y(n_1587)
);

AOI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1554),
.A2(n_1515),
.B1(n_1514),
.B2(n_1455),
.C(n_1508),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1526),
.B(n_1498),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1527),
.B(n_1498),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1527),
.B(n_1502),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1529),
.B(n_1484),
.Y(n_1592)
);

NOR3xp33_ASAP7_75t_L g1593 ( 
.A(n_1540),
.B(n_1478),
.C(n_1497),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1529),
.B(n_1484),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1562),
.B(n_1545),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1568),
.B(n_1545),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1564),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1563),
.B(n_1532),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1563),
.B(n_1547),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1565),
.Y(n_1601)
);

BUFx4f_ASAP7_75t_SL g1602 ( 
.A(n_1592),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1569),
.B(n_1549),
.Y(n_1603)
);

AND2x2_ASAP7_75t_SL g1604 ( 
.A(n_1560),
.B(n_1532),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1566),
.B(n_1522),
.Y(n_1605)
);

NAND2x1p5_ASAP7_75t_L g1606 ( 
.A(n_1594),
.B(n_1532),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1593),
.B(n_1532),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1582),
.Y(n_1608)
);

INVx4_ASAP7_75t_L g1609 ( 
.A(n_1581),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1556),
.B(n_1522),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1572),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1569),
.B(n_1549),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1575),
.Y(n_1613)
);

INVx4_ASAP7_75t_L g1614 ( 
.A(n_1581),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1576),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1567),
.B(n_1540),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1553),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1570),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1586),
.B(n_1578),
.Y(n_1619)
);

INVx3_ASAP7_75t_R g1620 ( 
.A(n_1583),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1588),
.B(n_1544),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1589),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1609),
.Y(n_1623)
);

NOR3xp33_ASAP7_75t_L g1624 ( 
.A(n_1610),
.B(n_1557),
.C(n_1577),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_L g1625 ( 
.A(n_1603),
.B(n_1558),
.C(n_1573),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1601),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1609),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1598),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1611),
.B(n_1615),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1609),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1618),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1618),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1603),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1599),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1604),
.A2(n_1558),
.B1(n_1559),
.B2(n_1573),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1611),
.B(n_1559),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1606),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1614),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1615),
.B(n_1590),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1598),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1598),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1612),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1608),
.B(n_1591),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1606),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1599),
.B(n_1607),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1608),
.B(n_1584),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1612),
.B(n_1585),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1595),
.B(n_1587),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1600),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1599),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1634),
.B(n_1599),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1629),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1629),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1644),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1626),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1626),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1647),
.B(n_1452),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1633),
.B(n_1595),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1633),
.B(n_1617),
.Y(n_1659)
);

OR2x6_ASAP7_75t_L g1660 ( 
.A(n_1644),
.B(n_1580),
.Y(n_1660)
);

AND2x2_ASAP7_75t_SL g1661 ( 
.A(n_1624),
.B(n_1625),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1642),
.B(n_1617),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1625),
.B(n_1613),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1642),
.B(n_1596),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1631),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1647),
.B(n_1622),
.Y(n_1666)
);

NAND2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1628),
.B(n_1604),
.Y(n_1667)
);

NAND2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1628),
.B(n_1604),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1650),
.B(n_1645),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1623),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1649),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1640),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1623),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1636),
.B(n_1596),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1623),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1636),
.B(n_1616),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1649),
.Y(n_1679)
);

INVx2_ASAP7_75t_SL g1680 ( 
.A(n_1650),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1645),
.B(n_1619),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1649),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1646),
.B(n_1622),
.Y(n_1683)
);

CKINVDCx16_ASAP7_75t_R g1684 ( 
.A(n_1635),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1624),
.A2(n_1606),
.B1(n_1571),
.B2(n_1605),
.C(n_1579),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1646),
.B(n_1640),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1648),
.B(n_1616),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1631),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1641),
.B(n_1639),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1680),
.Y(n_1690)
);

INVxp67_ASAP7_75t_SL g1691 ( 
.A(n_1674),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1673),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1669),
.B(n_1681),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1661),
.B(n_1684),
.C(n_1663),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1661),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1679),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1655),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1669),
.B(n_1644),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1654),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1682),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1652),
.B(n_1648),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1665),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1680),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1653),
.B(n_1648),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1676),
.B(n_1631),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1681),
.B(n_1645),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1657),
.B(n_1597),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1676),
.B(n_1632),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1667),
.B(n_1645),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1667),
.B(n_1637),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1665),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1671),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1654),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1671),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1656),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1678),
.B(n_1632),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1686),
.B(n_1641),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1675),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1678),
.B(n_1632),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1687),
.B(n_1639),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1689),
.B(n_1643),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1685),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1660),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1688),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1667),
.B(n_1637),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1694),
.A2(n_1635),
.B1(n_1668),
.B2(n_1621),
.C(n_1687),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1694),
.A2(n_1670),
.B1(n_1672),
.B2(n_1635),
.Y(n_1727)
);

NAND2x1_ASAP7_75t_L g1728 ( 
.A(n_1709),
.B(n_1670),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1691),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1695),
.A2(n_1668),
.B1(n_1621),
.B2(n_1666),
.C(n_1658),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1693),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1695),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1690),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1702),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1693),
.B(n_1670),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1702),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1699),
.B(n_1660),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1722),
.B(n_1683),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1709),
.B(n_1668),
.Y(n_1739)
);

NAND2xp33_ASAP7_75t_L g1740 ( 
.A(n_1725),
.B(n_1664),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1699),
.A2(n_1620),
.B1(n_1660),
.B2(n_1602),
.Y(n_1741)
);

OAI211xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1715),
.A2(n_1664),
.B(n_1658),
.C(n_1675),
.Y(n_1742)
);

OAI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1713),
.A2(n_1660),
.B1(n_1637),
.B2(n_1659),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1713),
.A2(n_1672),
.B1(n_1607),
.B2(n_1637),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_L g1745 ( 
.A(n_1697),
.B(n_1677),
.C(n_1662),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1711),
.Y(n_1746)
);

NAND4xp25_ASAP7_75t_L g1747 ( 
.A(n_1715),
.B(n_1672),
.C(n_1574),
.D(n_1662),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1710),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1724),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1724),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1729),
.Y(n_1752)
);

BUFx4f_ASAP7_75t_SL g1753 ( 
.A(n_1748),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1732),
.B(n_1717),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1734),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1738),
.B(n_1717),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1731),
.B(n_1726),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_R g1758 ( 
.A(n_1740),
.B(n_1341),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1726),
.B(n_1721),
.Y(n_1759)
);

CKINVDCx16_ASAP7_75t_R g1760 ( 
.A(n_1741),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1733),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1736),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_L g1763 ( 
.A(n_1737),
.B(n_1723),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1746),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1735),
.B(n_1706),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1728),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1745),
.B(n_1720),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1727),
.B(n_1721),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1739),
.B(n_1706),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1730),
.A2(n_1723),
.B1(n_1725),
.B2(n_1710),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1744),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1759),
.A2(n_1763),
.B(n_1770),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1760),
.A2(n_1730),
.B1(n_1742),
.B2(n_1747),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1757),
.A2(n_1742),
.B1(n_1743),
.B2(n_1701),
.C(n_1704),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1753),
.B(n_1707),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1771),
.B(n_1749),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1768),
.A2(n_1704),
.B1(n_1701),
.B2(n_1723),
.C(n_1720),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1767),
.A2(n_1703),
.B(n_1690),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1767),
.A2(n_1750),
.B(n_1751),
.C(n_1723),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1761),
.B(n_1698),
.Y(n_1780)
);

OAI21x1_ASAP7_75t_SL g1781 ( 
.A1(n_1766),
.A2(n_1703),
.B(n_1690),
.Y(n_1781)
);

NAND4xp25_ASAP7_75t_L g1782 ( 
.A(n_1754),
.B(n_1703),
.C(n_1698),
.D(n_1696),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1756),
.A2(n_1696),
.B(n_1692),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1775),
.B(n_1766),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1772),
.B(n_1752),
.C(n_1755),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1773),
.B(n_1765),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1780),
.Y(n_1787)
);

NAND5xp2_ASAP7_75t_L g1788 ( 
.A(n_1774),
.B(n_1769),
.C(n_1765),
.D(n_1764),
.E(n_1762),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1782),
.B(n_1769),
.Y(n_1789)
);

AOI211xp5_ASAP7_75t_L g1790 ( 
.A1(n_1777),
.A2(n_1758),
.B(n_1762),
.C(n_1692),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1781),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1776),
.B(n_1705),
.Y(n_1792)
);

INVx1_ASAP7_75t_SL g1793 ( 
.A(n_1778),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1783),
.Y(n_1794)
);

NOR4xp25_ASAP7_75t_L g1795 ( 
.A(n_1779),
.B(n_1700),
.C(n_1714),
.D(n_1712),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1784),
.B(n_1758),
.Y(n_1796)
);

OAI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1795),
.A2(n_1700),
.B(n_1422),
.C(n_1712),
.Y(n_1797)
);

NOR2x1_ASAP7_75t_L g1798 ( 
.A(n_1784),
.B(n_1712),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1786),
.B(n_1705),
.Y(n_1799)
);

NOR2x1_ASAP7_75t_L g1800 ( 
.A(n_1791),
.B(n_1714),
.Y(n_1800)
);

NOR4xp25_ASAP7_75t_L g1801 ( 
.A(n_1793),
.B(n_1714),
.C(n_1718),
.D(n_1677),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1798),
.Y(n_1802)
);

AOI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1799),
.A2(n_1787),
.B1(n_1792),
.B2(n_1785),
.Y(n_1803)
);

NOR2xp67_ASAP7_75t_L g1804 ( 
.A(n_1796),
.B(n_1794),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1800),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1797),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1801),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1798),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1805),
.Y(n_1809)
);

O2A1O1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1807),
.A2(n_1788),
.B(n_1789),
.C(n_1790),
.Y(n_1810)
);

NAND4xp75_ASAP7_75t_L g1811 ( 
.A(n_1804),
.B(n_1718),
.C(n_1583),
.D(n_1651),
.Y(n_1811)
);

CKINVDCx12_ASAP7_75t_R g1812 ( 
.A(n_1806),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1802),
.Y(n_1813)
);

CKINVDCx20_ASAP7_75t_R g1814 ( 
.A(n_1803),
.Y(n_1814)
);

NOR2x1_ASAP7_75t_L g1815 ( 
.A(n_1814),
.B(n_1808),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1813),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1811),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1815),
.Y(n_1818)
);

OR4x1_ASAP7_75t_L g1819 ( 
.A(n_1818),
.B(n_1809),
.C(n_1816),
.D(n_1812),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1819),
.B(n_1810),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1819),
.A2(n_1817),
.B1(n_1718),
.B2(n_1708),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1821),
.B(n_1817),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1820),
.A2(n_1708),
.B(n_1716),
.Y(n_1823)
);

NAND2xp33_ASAP7_75t_SL g1824 ( 
.A(n_1822),
.B(n_1716),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1823),
.A2(n_1719),
.B(n_1659),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1824),
.A2(n_1719),
.B(n_1627),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1825),
.B1(n_1688),
.B2(n_1630),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_SL g1828 ( 
.A1(n_1827),
.A2(n_1341),
.B1(n_1638),
.B2(n_1623),
.C(n_1627),
.Y(n_1828)
);

AOI211xp5_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1341),
.B(n_1627),
.C(n_1630),
.Y(n_1829)
);


endmodule