module fake_jpeg_11179_n_635 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_635);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_635;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_588;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_70),
.Y(n_184)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_75),
.Y(n_209)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_86),
.Y(n_134)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_17),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_29),
.B(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_29),
.B(n_17),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_97),
.Y(n_169)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_44),
.B(n_17),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_99),
.B(n_100),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_16),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_26),
.B(n_16),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_103),
.B(n_128),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_114),
.Y(n_193)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_119),
.Y(n_201)
);

INVx5_ASAP7_75t_SL g120 ( 
.A(n_55),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_120),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_20),
.Y(n_124)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_45),
.B(n_16),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_130),
.B(n_161),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_79),
.B(n_23),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_135),
.B(n_65),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_55),
.B1(n_33),
.B2(n_20),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_151),
.A2(n_78),
.B1(n_82),
.B2(n_87),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_66),
.A2(n_25),
.B1(n_21),
.B2(n_38),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_158),
.A2(n_178),
.B1(n_200),
.B2(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_69),
.B(n_46),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_93),
.A2(n_25),
.B1(n_38),
.B2(n_21),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_173),
.A2(n_176),
.B1(n_190),
.B2(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_76),
.B(n_28),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_175),
.B(n_194),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_68),
.A2(n_25),
.B1(n_38),
.B2(n_21),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_73),
.A2(n_38),
.B1(n_25),
.B2(n_43),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_179),
.B(n_56),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_77),
.A2(n_28),
.B1(n_60),
.B2(n_57),
.Y(n_182)
);

NAND2x1_ASAP7_75t_L g279 ( 
.A(n_182),
.B(n_19),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_79),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_75),
.B(n_33),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_187),
.B(n_51),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_83),
.A2(n_55),
.B1(n_60),
.B2(n_57),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_92),
.B(n_52),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_114),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_84),
.A2(n_62),
.B1(n_33),
.B2(n_55),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_85),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_117),
.Y(n_204)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_88),
.B(n_46),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_207),
.B(n_22),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_91),
.A2(n_62),
.B1(n_41),
.B2(n_52),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_96),
.A2(n_37),
.B1(n_51),
.B2(n_41),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_214),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_215),
.B(n_220),
.Y(n_289)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_217),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_131),
.B(n_124),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_221),
.B(n_240),
.Y(n_311)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_222),
.Y(n_303)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_137),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_223),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_133),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

NAND2x1p5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_129),
.Y(n_226)
);

NOR2x1_ASAP7_75t_SL g336 ( 
.A(n_226),
.B(n_30),
.Y(n_336)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_227),
.Y(n_297)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_228),
.Y(n_322)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_229),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_230),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

INVx8_ASAP7_75t_L g335 ( 
.A(n_231),
.Y(n_335)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_132),
.Y(n_232)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_143),
.Y(n_234)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_234),
.Y(n_302)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_156),
.Y(n_236)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_148),
.A2(n_80),
.B1(n_74),
.B2(n_67),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_238),
.A2(n_258),
.B1(n_280),
.B2(n_282),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_138),
.Y(n_239)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

AND2x2_ASAP7_75t_SL g240 ( 
.A(n_165),
.B(n_101),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_242),
.B(n_256),
.Y(n_295)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_245),
.B(n_259),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_157),
.Y(n_248)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_248),
.Y(n_318)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_190),
.A2(n_127),
.B1(n_125),
.B2(n_123),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_250),
.A2(n_252),
.B1(n_262),
.B2(n_206),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_212),
.A2(n_121),
.B1(n_118),
.B2(n_111),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_253),
.Y(n_327)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_254),
.Y(n_343)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_165),
.Y(n_255)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_255),
.Y(n_345)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_257),
.B(n_260),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_148),
.A2(n_110),
.B1(n_109),
.B2(n_104),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_162),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_158),
.A2(n_37),
.B1(n_50),
.B2(n_32),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_261),
.A2(n_180),
.B1(n_170),
.B2(n_163),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_139),
.A2(n_56),
.B1(n_50),
.B2(n_32),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_144),
.Y(n_263)
);

BUFx24_ASAP7_75t_L g321 ( 
.A(n_263),
.Y(n_321)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_145),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_265),
.Y(n_305)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_146),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_266),
.Y(n_329)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_168),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_267),
.Y(n_313)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_147),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_268),
.B(n_269),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_149),
.Y(n_269)
);

BUFx4f_ASAP7_75t_SL g270 ( 
.A(n_193),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_284),
.Y(n_290)
);

INVx4_ASAP7_75t_SL g271 ( 
.A(n_209),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_271),
.Y(n_328)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_197),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_272),
.B(n_273),
.Y(n_310)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_172),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_160),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_274),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_275),
.B(n_276),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_139),
.B(n_22),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_277),
.B(n_278),
.Y(n_339)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_164),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_279),
.A2(n_245),
.B1(n_240),
.B2(n_285),
.Y(n_325)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_159),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_177),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_281),
.B(n_283),
.Y(n_320)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_166),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_134),
.B(n_19),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_134),
.B(n_15),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_169),
.B(n_15),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_183),
.C(n_182),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_177),
.B(n_14),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_169),
.B(n_14),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_192),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_288),
.A2(n_201),
.B1(n_191),
.B2(n_204),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_151),
.B(n_187),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_291),
.A2(n_10),
.B(n_2),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_292),
.B(n_336),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_243),
.B(n_182),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_301),
.B(n_330),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_270),
.C(n_280),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_314),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_250),
.A2(n_206),
.B1(n_203),
.B2(n_168),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_315),
.A2(n_340),
.B1(n_231),
.B2(n_230),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_226),
.B(n_150),
.C(n_191),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_323),
.B(n_337),
.C(n_3),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_325),
.A2(n_338),
.B(n_246),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_225),
.B(n_140),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_247),
.A2(n_174),
.B1(n_198),
.B2(n_199),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_332),
.A2(n_347),
.B1(n_349),
.B2(n_221),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g337 ( 
.A(n_221),
.B(n_0),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_240),
.A2(n_141),
.B1(n_195),
.B2(n_198),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_251),
.A2(n_203),
.B1(n_188),
.B2(n_185),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_263),
.B(n_188),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_346),
.B(n_241),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_247),
.A2(n_237),
.B1(n_258),
.B2(n_261),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_224),
.A2(n_185),
.B1(n_180),
.B2(n_170),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_348),
.A2(n_239),
.B1(n_269),
.B2(n_249),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_277),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_350),
.B(n_377),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_326),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g352 ( 
.A(n_323),
.B(n_221),
.CI(n_233),
.CON(n_352),
.SN(n_352)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_352),
.B(n_376),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_340),
.A2(n_301),
.B1(n_292),
.B2(n_291),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_353),
.A2(n_356),
.B1(n_357),
.B2(n_360),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_218),
.B1(n_259),
.B2(n_267),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_354),
.A2(n_364),
.B1(n_365),
.B2(n_375),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_355),
.A2(n_358),
.B1(n_359),
.B2(n_361),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_307),
.A2(n_238),
.B1(n_154),
.B2(n_163),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_309),
.A2(n_153),
.B1(n_154),
.B2(n_223),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_282),
.B1(n_274),
.B2(n_268),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_309),
.A2(n_265),
.B1(n_222),
.B2(n_227),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_153),
.B1(n_254),
.B2(n_234),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_346),
.Y(n_362)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_326),
.Y(n_363)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_311),
.A2(n_214),
.B1(n_229),
.B2(n_219),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_311),
.A2(n_271),
.B(n_216),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_366),
.A2(n_386),
.B(n_394),
.Y(n_398)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_396),
.C(n_366),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_372),
.Y(n_397)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_345),
.Y(n_370)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_370),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_320),
.B(n_228),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_373),
.B(n_388),
.Y(n_418)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_311),
.A2(n_270),
.B1(n_30),
.B2(n_13),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_321),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_329),
.Y(n_377)
);

BUFx8_ASAP7_75t_L g378 ( 
.A(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_293),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_380),
.B(n_387),
.Y(n_405)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_381),
.A2(n_351),
.B1(n_363),
.B2(n_335),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_328),
.B(n_244),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_382),
.B(n_304),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_330),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_383),
.A2(n_384),
.B1(n_337),
.B2(n_356),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_325),
.A2(n_306),
.B1(n_338),
.B2(n_290),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_341),
.A2(n_13),
.B1(n_10),
.B2(n_9),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_385),
.A2(n_395),
.B1(n_317),
.B2(n_304),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_324),
.B(n_10),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_289),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_297),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_391),
.Y(n_410)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_297),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_321),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_393),
.Y(n_413)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_290),
.A2(n_10),
.B(n_3),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_337),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_396),
.B(n_298),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_400),
.B(n_403),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_389),
.B(n_341),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_377),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_404),
.B(n_406),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_350),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_408),
.B(n_409),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_382),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_412),
.A2(n_423),
.B1(n_435),
.B2(n_359),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_372),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_415),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_341),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_419),
.B(n_421),
.Y(n_439)
);

BUFx24_ASAP7_75t_SL g420 ( 
.A(n_388),
.Y(n_420)
);

BUFx24_ASAP7_75t_SL g462 ( 
.A(n_420),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_368),
.B(n_295),
.C(n_312),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_353),
.A2(n_313),
.B1(n_316),
.B2(n_308),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_366),
.A2(n_394),
.B(n_386),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_424),
.A2(n_398),
.B(n_418),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_384),
.A2(n_298),
.B1(n_313),
.B2(n_343),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_425),
.A2(n_319),
.B(n_317),
.Y(n_469)
);

OAI32xp33_ASAP7_75t_L g427 ( 
.A1(n_362),
.A2(n_299),
.A3(n_331),
.B1(n_305),
.B2(n_339),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_436),
.Y(n_449)
);

OR2x6_ASAP7_75t_L g458 ( 
.A(n_428),
.B(n_411),
.Y(n_458)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_432),
.B(n_387),
.C(n_310),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_355),
.A2(n_361),
.B1(n_371),
.B2(n_352),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_433),
.A2(n_371),
.B1(n_352),
.B2(n_360),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_368),
.B(n_316),
.C(n_312),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_434),
.B(n_373),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_371),
.A2(n_318),
.B1(n_343),
.B2(n_300),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_369),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_437),
.Y(n_486)
);

AO21x1_ASAP7_75t_L g479 ( 
.A1(n_438),
.A2(n_446),
.B(n_461),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_441),
.B(n_469),
.Y(n_494)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_413),
.Y(n_442)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

OAI32xp33_ASAP7_75t_L g443 ( 
.A1(n_426),
.A2(n_415),
.A3(n_402),
.B1(n_397),
.B2(n_417),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_445),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_444),
.A2(n_458),
.B1(n_464),
.B2(n_472),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_410),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_426),
.A2(n_352),
.B(n_374),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_429),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_450),
.A2(n_455),
.B(n_465),
.Y(n_475)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_429),
.Y(n_452)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_452),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_370),
.Y(n_453)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_453),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_454),
.A2(n_456),
.B1(n_460),
.B2(n_401),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_398),
.A2(n_379),
.B(n_351),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_407),
.A2(n_379),
.B1(n_358),
.B2(n_395),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_397),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_457),
.B(n_466),
.Y(n_493)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_459),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_407),
.A2(n_393),
.B1(n_385),
.B2(n_380),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_418),
.A2(n_391),
.B(n_390),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_383),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_463),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_433),
.A2(n_357),
.B1(n_367),
.B2(n_381),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_363),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_418),
.A2(n_392),
.B(n_376),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_467),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_418),
.A2(n_333),
.B(n_318),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_427),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_404),
.B(n_333),
.Y(n_472)
);

AO22x1_ASAP7_75t_SL g473 ( 
.A1(n_437),
.A2(n_402),
.B1(n_401),
.B2(n_423),
.Y(n_473)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_473),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_474),
.A2(n_477),
.B1(n_480),
.B2(n_303),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_448),
.A2(n_425),
.B1(n_408),
.B2(n_412),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_454),
.A2(n_424),
.B1(n_436),
.B2(n_400),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_478),
.A2(n_489),
.B1(n_492),
.B2(n_457),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_448),
.A2(n_411),
.B1(n_435),
.B2(n_405),
.Y(n_480)
);

XNOR2x1_ASAP7_75t_L g514 ( 
.A(n_481),
.B(n_504),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_439),
.C(n_441),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_482),
.B(n_488),
.C(n_468),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_444),
.A2(n_434),
.B1(n_421),
.B2(n_405),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_483),
.A2(n_499),
.B1(n_470),
.B2(n_461),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_419),
.C(n_403),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_460),
.A2(n_442),
.B1(n_456),
.B2(n_451),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_445),
.A2(n_403),
.B1(n_406),
.B2(n_432),
.Y(n_492)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_447),
.Y(n_496)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_496),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_419),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_501),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_449),
.A2(n_428),
.B1(n_422),
.B2(n_399),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_439),
.B(n_446),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_422),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_503),
.B(n_505),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_440),
.B(n_431),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_443),
.B(n_327),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_506),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_507),
.B(n_528),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_508),
.A2(n_479),
.B1(n_485),
.B2(n_500),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_453),
.C(n_468),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_509),
.B(n_517),
.C(n_521),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_511),
.A2(n_473),
.B1(n_502),
.B2(n_496),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_474),
.A2(n_458),
.B1(n_464),
.B2(n_440),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_513),
.A2(n_515),
.B1(n_518),
.B2(n_526),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_489),
.A2(n_458),
.B1(n_438),
.B2(n_465),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_493),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_516),
.B(n_519),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_498),
.B(n_467),
.C(n_472),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_492),
.A2(n_458),
.B1(n_465),
.B2(n_463),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_450),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_493),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_520),
.B(n_522),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_469),
.C(n_455),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_483),
.B(n_462),
.Y(n_522)
);

FAx1_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_458),
.CI(n_459),
.CON(n_523),
.SN(n_523)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_523),
.A2(n_529),
.B(n_506),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_493),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_525),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_466),
.C(n_452),
.Y(n_525)
);

AOI211xp5_ASAP7_75t_L g526 ( 
.A1(n_476),
.A2(n_458),
.B(n_431),
.C(n_416),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_494),
.B(n_319),
.C(n_416),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_478),
.B(n_458),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_504),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_327),
.C(n_334),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_503),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_531),
.A2(n_499),
.B1(n_481),
.B2(n_491),
.Y(n_547)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_497),
.Y(n_532)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_532),
.Y(n_536)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_484),
.Y(n_533)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_533),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_537),
.B(n_540),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_538),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_508),
.A2(n_475),
.B(n_490),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_542),
.A2(n_513),
.B1(n_515),
.B2(n_511),
.Y(n_565)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_512),
.Y(n_545)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_545),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_547),
.A2(n_558),
.B1(n_514),
.B2(n_527),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_534),
.A2(n_486),
.B1(n_487),
.B2(n_495),
.Y(n_548)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_548),
.Y(n_575)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_532),
.Y(n_549)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_549),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_530),
.Y(n_569)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_533),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_551),
.Y(n_578)
);

BUFx24_ASAP7_75t_SL g552 ( 
.A(n_523),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_552),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_553),
.A2(n_526),
.B1(n_520),
.B2(n_523),
.Y(n_561)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_512),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_557),
.Y(n_560)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_534),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_518),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_539),
.B(n_546),
.C(n_507),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_562),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_561),
.A2(n_571),
.B1(n_344),
.B2(n_322),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_539),
.B(n_509),
.C(n_525),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_565),
.A2(n_572),
.B1(n_576),
.B2(n_302),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_541),
.A2(n_521),
.B1(n_517),
.B2(n_473),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_569),
.B(n_573),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_528),
.C(n_510),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_570),
.B(n_537),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_541),
.A2(n_514),
.B1(n_527),
.B2(n_510),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_542),
.A2(n_544),
.B1(n_558),
.B2(n_547),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_550),
.B(n_540),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_574),
.B(n_553),
.C(n_535),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_544),
.A2(n_335),
.B1(n_342),
.B2(n_302),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_564),
.B(n_555),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_579),
.B(n_581),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_577),
.A2(n_554),
.B(n_538),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_580),
.A2(n_584),
.B(n_588),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_582),
.B(n_591),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_559),
.B(n_545),
.C(n_543),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_583),
.B(n_569),
.C(n_566),
.Y(n_604)
);

AOI21x1_ASAP7_75t_L g584 ( 
.A1(n_577),
.A2(n_536),
.B(n_334),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_587),
.A2(n_567),
.B1(n_563),
.B2(n_568),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_562),
.B(n_300),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_590),
.B(n_592),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_565),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_575),
.B(n_300),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_572),
.A2(n_296),
.B(n_378),
.Y(n_593)
);

NAND3xp33_ASAP7_75t_SL g599 ( 
.A(n_593),
.B(n_560),
.C(n_561),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_342),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_594),
.A2(n_578),
.B(n_560),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_578),
.B(n_378),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_595),
.A2(n_578),
.B1(n_563),
.B2(n_568),
.Y(n_597)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_597),
.Y(n_609)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_598),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_604),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_600),
.A2(n_587),
.B1(n_593),
.B2(n_589),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_586),
.A2(n_570),
.B(n_576),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_602),
.A2(n_606),
.B(n_583),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_566),
.C(n_571),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_585),
.A2(n_342),
.B1(n_344),
.B2(n_322),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_607),
.B(n_608),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_580),
.A2(n_321),
.B(n_378),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_608),
.A2(n_584),
.B(n_595),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_610),
.A2(n_615),
.B(n_617),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_611),
.B(n_612),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_605),
.A2(n_582),
.B(n_589),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_616),
.B(n_596),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_604),
.A2(n_294),
.B(n_296),
.Y(n_617)
);

AOI21x1_ASAP7_75t_L g618 ( 
.A1(n_601),
.A2(n_294),
.B(n_5),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_618),
.A2(n_4),
.B(n_5),
.Y(n_622)
);

INVx6_ASAP7_75t_L g619 ( 
.A(n_613),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_619),
.B(n_622),
.Y(n_626)
);

AOI31xp33_ASAP7_75t_L g620 ( 
.A1(n_614),
.A2(n_599),
.A3(n_606),
.B(n_600),
.Y(n_620)
);

AO221x1_ASAP7_75t_L g628 ( 
.A1(n_620),
.A2(n_623),
.B1(n_4),
.B2(n_6),
.C(n_7),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g623 ( 
.A(n_609),
.B(n_603),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_625),
.B(n_4),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_624),
.B(n_616),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_627),
.A2(n_628),
.B(n_629),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_626),
.B(n_621),
.C(n_623),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_630),
.B(n_6),
.Y(n_632)
);

BUFx24_ASAP7_75t_SL g633 ( 
.A(n_632),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_633),
.A2(n_631),
.B(n_7),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g635 ( 
.A1(n_634),
.A2(n_6),
.B1(n_8),
.B2(n_578),
.Y(n_635)
);


endmodule