module fake_jpeg_17101_n_358 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_358);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_358;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_16),
.B(n_15),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_23),
.CON(n_40),
.SN(n_40)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_40),
.A2(n_19),
.B1(n_35),
.B2(n_34),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_25),
.B1(n_29),
.B2(n_38),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_59),
.B1(n_62),
.B2(n_23),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_25),
.B1(n_37),
.B2(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_24),
.B1(n_29),
.B2(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_37),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_38),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_19),
.Y(n_84)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_99),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_37),
.B1(n_28),
.B2(n_31),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_69),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_34),
.B1(n_27),
.B2(n_26),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_27),
.B1(n_26),
.B2(n_68),
.Y(n_121)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_49),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_33),
.CI(n_30),
.CON(n_138),
.SN(n_138)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_32),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_113),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_65),
.B(n_79),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_115),
.A2(n_119),
.B(n_28),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_72),
.B(n_57),
.C(n_74),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_139),
.B(n_70),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_100),
.B(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_121),
.B(n_138),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_105),
.B1(n_58),
.B2(n_84),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_128),
.B1(n_103),
.B2(n_83),
.Y(n_144)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_132),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_86),
.A2(n_74),
.B1(n_63),
.B2(n_41),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_28),
.B1(n_33),
.B2(n_31),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_89),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_81),
.B1(n_37),
.B2(n_83),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_86),
.B(n_28),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_102),
.C(n_28),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_32),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_144),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_147),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_140),
.A2(n_90),
.B1(n_102),
.B2(n_81),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_150),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_127),
.B1(n_138),
.B2(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_149),
.A2(n_151),
.B1(n_162),
.B2(n_168),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_96),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_70),
.B1(n_41),
.B2(n_73),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_56),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_163),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_110),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_73),
.B1(n_98),
.B2(n_109),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_156),
.B1(n_132),
.B2(n_118),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_73),
.B1(n_93),
.B2(n_33),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_93),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_33),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_31),
.B(n_30),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_128),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_126),
.A2(n_31),
.B1(n_30),
.B2(n_22),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_174),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_173),
.A2(n_184),
.B(n_151),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_121),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_195),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_137),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_181),
.C(n_189),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_114),
.C(n_117),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_187),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_110),
.C(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_118),
.C(n_125),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_196),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_164),
.A2(n_136),
.B1(n_154),
.B2(n_159),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_156),
.B(n_141),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_158),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_198),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_165),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_210),
.C(n_217),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_150),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_191),
.Y(n_233)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_227),
.Y(n_228)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_178),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_214),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_152),
.C(n_144),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_142),
.Y(n_211)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_153),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_223),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_173),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_155),
.C(n_169),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_170),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_129),
.B1(n_120),
.B2(n_168),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_172),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_225),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_147),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_175),
.B(n_177),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_229),
.A2(n_230),
.B(n_246),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_196),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_203),
.B(n_211),
.C(n_200),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_189),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_185),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_185),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_175),
.B1(n_191),
.B2(n_188),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_241),
.B1(n_255),
.B2(n_205),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_146),
.B1(n_167),
.B2(n_136),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_199),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_204),
.A2(n_227),
.B(n_201),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_202),
.B(n_32),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_248),
.B(n_120),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_129),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_219),
.A2(n_217),
.B1(n_213),
.B2(n_210),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_216),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_270),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_246),
.B(n_215),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_207),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_6),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_199),
.C(n_224),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_228),
.C(n_238),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_30),
.B1(n_1),
.B2(n_4),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_279),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_275),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_240),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_254),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_295),
.C(n_296),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_256),
.A2(n_250),
.B1(n_232),
.B2(n_251),
.Y(n_284)
);

OAI22x1_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_274),
.B1(n_259),
.B2(n_257),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_256),
.A2(n_244),
.B1(n_230),
.B2(n_239),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_285),
.A2(n_293),
.B1(n_281),
.B2(n_269),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_251),
.B1(n_233),
.B2(n_230),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_241),
.B(n_228),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_293),
.A2(n_7),
.B(n_8),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_32),
.C(n_5),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_1),
.C(n_5),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_278),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_297),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_301),
.A2(n_310),
.B1(n_9),
.B2(n_10),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_286),
.B(n_261),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_309),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_304),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_285),
.B(n_270),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_268),
.B1(n_258),
.B2(n_263),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_283),
.C(n_295),
.Y(n_315)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_308),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_290),
.B(n_263),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_287),
.B(n_6),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_6),
.B(n_7),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_314),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_9),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_8),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_304),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_296),
.C(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_319),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_284),
.B(n_281),
.Y(n_320)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_305),
.A2(n_298),
.B1(n_292),
.B2(n_288),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_322),
.B(n_325),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_8),
.Y(n_323)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_323),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_326),
.B(n_328),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_335),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_336),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_320),
.A2(n_10),
.B(n_11),
.Y(n_333)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_333),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_10),
.B(n_11),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_319),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_337),
.A2(n_11),
.B(n_13),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g341 ( 
.A1(n_336),
.A2(n_316),
.B(n_327),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_341),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_321),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_343),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_318),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_344),
.A2(n_331),
.B(n_338),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_346),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_13),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_350),
.B(n_351),
.C(n_14),
.Y(n_354)
);

A2O1A1O1Ixp25_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_14),
.B(n_339),
.C(n_345),
.D(n_340),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_354),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_353),
.C(n_349),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_352),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_347),
.Y(n_358)
);


endmodule