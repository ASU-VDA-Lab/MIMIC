module fake_jpeg_6318_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_47),
.B1(n_28),
.B2(n_29),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_1),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_24),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_23),
.B(n_1),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_54),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_23),
.Y(n_52)
);

NAND2x1_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_17),
.Y(n_53)
);

AOI32xp33_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_17),
.A3(n_47),
.B1(n_35),
.B2(n_44),
.Y(n_92)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_59),
.B1(n_65),
.B2(n_39),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_47),
.B1(n_37),
.B2(n_44),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_27),
.B1(n_18),
.B2(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_66),
.Y(n_76)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_18),
.B1(n_32),
.B2(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_41),
.B1(n_20),
.B2(n_34),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_73),
.Y(n_129)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_75),
.B(n_81),
.Y(n_127)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_16),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_30),
.B1(n_31),
.B2(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_85),
.C(n_98),
.Y(n_108)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_87),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_97),
.B1(n_101),
.B2(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_93),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_51),
.A2(n_37),
.B1(n_44),
.B2(n_43),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_37),
.B1(n_59),
.B2(n_57),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_18),
.B1(n_43),
.B2(n_30),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_17),
.A3(n_43),
.B1(n_35),
.B2(n_36),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_35),
.Y(n_112)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_50),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_103),
.Y(n_143)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_116),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_128),
.B1(n_77),
.B2(n_82),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_67),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_79),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_120),
.B1(n_75),
.B2(n_20),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_84),
.A2(n_61),
.B1(n_50),
.B2(n_48),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_56),
.B(n_65),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_36),
.C(n_49),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_93),
.C(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_131),
.B(n_134),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_137),
.C(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_136),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_89),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_139),
.B(n_141),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_115),
.C(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_142),
.A2(n_146),
.B1(n_45),
.B2(n_24),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_89),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_71),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g180 ( 
.A(n_145),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_108),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_157),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_152),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_76),
.C(n_72),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_78),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_123),
.B(n_88),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_78),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_16),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_123),
.B(n_88),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_114),
.B(n_105),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_114),
.B(n_105),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_105),
.B1(n_112),
.B2(n_73),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_167),
.A2(n_171),
.B1(n_194),
.B2(n_158),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_191),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_54),
.B1(n_64),
.B2(n_116),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_126),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_178),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_125),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_64),
.B1(n_54),
.B2(n_91),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_193),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_100),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_185),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_31),
.B1(n_26),
.B2(n_103),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_183),
.B(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_74),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_36),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_131),
.C(n_135),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_45),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_133),
.B(n_74),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_133),
.B(n_45),
.CI(n_36),
.CON(n_195),
.SN(n_195)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_25),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_203),
.C(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_147),
.C(n_49),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_49),
.C(n_136),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_216),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_213),
.B(n_218),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_163),
.A2(n_150),
.B1(n_117),
.B2(n_21),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_173),
.B1(n_176),
.B2(n_25),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_169),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_219),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_168),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_225),
.Y(n_233)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_223),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_182),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_138),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_226),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_45),
.Y(n_225)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_25),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_181),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_230),
.B(n_248),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_191),
.B1(n_162),
.B2(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_162),
.B1(n_188),
.B2(n_193),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_232),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_205),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_237),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_164),
.B(n_167),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_243),
.B(n_244),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_195),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_220),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_207),
.B(n_198),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_198),
.A2(n_188),
.B1(n_189),
.B2(n_195),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_186),
.B(n_196),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_210),
.B(n_203),
.Y(n_258)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_186),
.A3(n_165),
.B1(n_173),
.B2(n_25),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_210),
.B(n_165),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_10),
.B1(n_14),
.B2(n_5),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_198),
.A2(n_176),
.B1(n_155),
.B2(n_154),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_21),
.B1(n_24),
.B2(n_22),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_261),
.C(n_268),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_271),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_246),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_258),
.A2(n_228),
.B(n_241),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_208),
.C(n_197),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_267),
.Y(n_286)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_22),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_266),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_2),
.C(n_3),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_9),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_242),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_270),
.B(n_244),
.Y(n_277)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_271),
.B1(n_269),
.B2(n_253),
.Y(n_292)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_242),
.C(n_248),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_254),
.C(n_257),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_238),
.B(n_235),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_289),
.B1(n_7),
.B2(n_8),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_236),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_252),
.B(n_235),
.Y(n_284)
);

AO221x1_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_227),
.B1(n_247),
.B2(n_229),
.C(n_243),
.Y(n_287)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_234),
.B1(n_239),
.B2(n_3),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_295),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_259),
.B1(n_253),
.B2(n_258),
.Y(n_293)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_297),
.C(n_299),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_257),
.C(n_265),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_3),
.C(n_4),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_4),
.B1(n_15),
.B2(n_7),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_6),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_302),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_282),
.C(n_276),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_282),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_296),
.B(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_306),
.B(n_311),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_295),
.C(n_297),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_285),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_308),
.B(n_316),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_285),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_278),
.B(n_290),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_288),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_281),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_310),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_324),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_320),
.B(n_321),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_294),
.C(n_303),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_322),
.A2(n_325),
.B1(n_309),
.B2(n_305),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_307),
.B(n_278),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_312),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_313),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_330),
.B(n_11),
.C(n_12),
.Y(n_334)
);

AO221x1_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_312),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_332),
.B(n_334),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_335),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_333),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_330),
.Y(n_339)
);


endmodule