module fake_jpeg_14409_n_38 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_5),
.B(n_7),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_21),
.B1(n_14),
.B2(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_19),
.B1(n_20),
.B2(n_14),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_0),
.C(n_1),
.Y(n_18)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_14),
.A3(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

OR2x2_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_16),
.A2(n_10),
.B1(n_12),
.B2(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_27),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_26),
.C(n_23),
.Y(n_35)
);

AOI322xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.A3(n_33),
.B1(n_24),
.B2(n_20),
.C1(n_17),
.C2(n_8),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_4),
.C(n_5),
.Y(n_38)
);


endmodule