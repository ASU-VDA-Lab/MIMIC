module fake_jpeg_19762_n_56 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx4_ASAP7_75t_SL g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_20),
.A2(n_14),
.B1(n_11),
.B2(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_17),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_13),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_18),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_35),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_9),
.C(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_4),
.Y(n_43)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_19),
.B1(n_12),
.B2(n_16),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_9),
.B1(n_16),
.B2(n_10),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_4),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_31),
.B1(n_37),
.B2(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_50),
.B(n_40),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_41),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_51),
.C(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);


endmodule