module fake_jpeg_14311_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

CKINVDCx14_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_19),
.B1(n_12),
.B2(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_18),
.B(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_5),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_8),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_25),
.Y(n_35)
);

BUFx24_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_9),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_32),
.B1(n_29),
.B2(n_24),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_17),
.B1(n_16),
.B2(n_12),
.Y(n_32)
);

AND2x6_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_7),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_28),
.B(n_29),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.C(n_35),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.C(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_34),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_40),
.B1(n_30),
.B2(n_24),
.Y(n_46)
);

MAJx2_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_7),
.C(n_37),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_7),
.Y(n_48)
);


endmodule