module real_aes_8780_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g171 ( .A1(n_0), .A2(n_172), .B(n_175), .C(n_179), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_1), .B(n_163), .Y(n_182) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_3), .B(n_173), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_4), .A2(n_136), .B(n_139), .C(n_503), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_5), .A2(n_131), .B(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_6), .A2(n_131), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_7), .B(n_163), .Y(n_534) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_8), .A2(n_165), .B(n_237), .Y(n_236) );
AND2x6_ASAP7_75t_L g136 ( .A(n_9), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_10), .A2(n_136), .B(n_139), .C(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g494 ( .A(n_11), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_12), .B(n_39), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_13), .B(n_178), .Y(n_505) );
INVx1_ASAP7_75t_L g157 ( .A(n_14), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_15), .B(n_173), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_16), .A2(n_174), .B(n_514), .C(n_516), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_17), .B(n_163), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_18), .B(n_151), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_19), .A2(n_139), .B(n_142), .C(n_150), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_20), .A2(n_177), .B(n_245), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_21), .B(n_178), .Y(n_479) );
AOI222xp33_ASAP7_75t_L g113 ( .A1(n_22), .A2(n_74), .B1(n_114), .B2(n_725), .C1(n_728), .C2(n_729), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_23), .B(n_178), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_24), .Y(n_475) );
INVx1_ASAP7_75t_L g455 ( .A(n_25), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_26), .A2(n_139), .B(n_150), .C(n_240), .Y(n_239) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_27), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_28), .Y(n_501) );
INVx1_ASAP7_75t_L g469 ( .A(n_29), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_30), .A2(n_131), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g134 ( .A(n_31), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_32), .A2(n_189), .B(n_190), .C(n_194), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_33), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_34), .A2(n_177), .B(n_531), .C(n_533), .Y(n_530) );
INVxp67_ASAP7_75t_L g470 ( .A(n_35), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_36), .B(n_242), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_37), .A2(n_139), .B(n_150), .C(n_454), .Y(n_453) );
CKINVDCx14_ASAP7_75t_R g529 ( .A(n_38), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_40), .A2(n_179), .B(n_492), .C(n_493), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_41), .B(n_130), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_42), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_43), .B(n_173), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_44), .B(n_131), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_45), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_46), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_47), .B(n_744), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_48), .A2(n_189), .B(n_194), .C(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g176 ( .A(n_49), .Y(n_176) );
INVx1_ASAP7_75t_L g220 ( .A(n_50), .Y(n_220) );
INVx1_ASAP7_75t_L g542 ( .A(n_51), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_52), .B(n_131), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_53), .Y(n_159) );
CKINVDCx14_ASAP7_75t_R g490 ( .A(n_54), .Y(n_490) );
INVx1_ASAP7_75t_L g137 ( .A(n_55), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_56), .B(n_131), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_57), .B(n_163), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_58), .A2(n_149), .B(n_205), .C(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g156 ( .A(n_59), .Y(n_156) );
INVx1_ASAP7_75t_SL g532 ( .A(n_60), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_61), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_62), .B(n_173), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_63), .B(n_163), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_64), .B(n_174), .Y(n_255) );
INVx1_ASAP7_75t_L g478 ( .A(n_65), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_66), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_67), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_68), .A2(n_139), .B(n_194), .C(n_203), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_69), .Y(n_229) );
INVx1_ASAP7_75t_L g103 ( .A(n_70), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_71), .A2(n_131), .B(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_72), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_73), .A2(n_131), .B(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_74), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_75), .A2(n_130), .B(n_465), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_76), .Y(n_452) );
INVx1_ASAP7_75t_L g512 ( .A(n_77), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_78), .B(n_147), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_79), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_80), .A2(n_131), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g515 ( .A(n_81), .Y(n_515) );
INVx2_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
INVx1_ASAP7_75t_L g504 ( .A(n_83), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_84), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_85), .B(n_178), .Y(n_256) );
OR2x2_ASAP7_75t_L g107 ( .A(n_86), .B(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g117 ( .A(n_86), .B(n_109), .Y(n_117) );
INVx2_ASAP7_75t_L g444 ( .A(n_86), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_87), .A2(n_139), .B(n_194), .C(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_88), .B(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g191 ( .A(n_89), .Y(n_191) );
INVxp67_ASAP7_75t_L g232 ( .A(n_90), .Y(n_232) );
AOI222xp33_ASAP7_75t_SL g98 ( .A1(n_91), .A2(n_99), .B1(n_112), .B2(n_732), .C1(n_737), .C2(n_746), .Y(n_98) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_91), .A2(n_119), .B1(n_739), .B2(n_740), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_91), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_92), .B(n_165), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_93), .B(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g204 ( .A(n_94), .Y(n_204) );
INVx1_ASAP7_75t_L g251 ( .A(n_95), .Y(n_251) );
INVx2_ASAP7_75t_L g545 ( .A(n_96), .Y(n_545) );
AND2x2_ASAP7_75t_L g222 ( .A(n_97), .B(n_153), .Y(n_222) );
INVx1_ASAP7_75t_SL g99 ( .A(n_100), .Y(n_99) );
NAND2xp33_ASAP7_75t_L g100 ( .A(n_101), .B(n_105), .Y(n_100) );
NOR2xp33_ASAP7_75t_SL g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx1_ASAP7_75t_SL g736 ( .A(n_102), .Y(n_736) );
INVx1_ASAP7_75t_L g735 ( .A(n_104), .Y(n_735) );
OA21x2_ASAP7_75t_L g747 ( .A1(n_104), .A2(n_736), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_107), .Y(n_742) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_107), .Y(n_745) );
BUFx2_ASAP7_75t_L g748 ( .A(n_107), .Y(n_748) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_108), .B(n_444), .Y(n_731) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g443 ( .A(n_109), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B1(n_441), .B2(n_445), .Y(n_114) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_115), .A2(n_119), .B1(n_726), .B2(n_727), .Y(n_725) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g740 ( .A(n_119), .Y(n_740) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_396), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_331), .Y(n_120) );
NAND4xp25_ASAP7_75t_SL g121 ( .A(n_122), .B(n_276), .C(n_300), .D(n_323), .Y(n_121) );
AOI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_213), .B1(n_247), .B2(n_260), .C(n_263), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_183), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_125), .A2(n_161), .B1(n_214), .B2(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_125), .B(n_184), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_125), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_125), .B(n_337), .Y(n_423) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
AND2x2_ASAP7_75t_L g291 ( .A(n_126), .B(n_184), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_126), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g314 ( .A(n_126), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_126), .B(n_162), .Y(n_319) );
INVx2_ASAP7_75t_L g351 ( .A(n_126), .Y(n_351) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_126), .Y(n_395) );
AND2x2_ASAP7_75t_L g412 ( .A(n_126), .B(n_289), .Y(n_412) );
INVx5_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g330 ( .A(n_127), .B(n_289), .Y(n_330) );
AND2x4_ASAP7_75t_L g344 ( .A(n_127), .B(n_161), .Y(n_344) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_127), .Y(n_348) );
AND2x2_ASAP7_75t_L g368 ( .A(n_127), .B(n_283), .Y(n_368) );
AND2x2_ASAP7_75t_L g418 ( .A(n_127), .B(n_185), .Y(n_418) );
AND2x2_ASAP7_75t_L g428 ( .A(n_127), .B(n_162), .Y(n_428) );
OR2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_158), .Y(n_127) );
AOI21xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_138), .B(n_151), .Y(n_128) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_132), .B(n_136), .Y(n_252) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx1_ASAP7_75t_L g246 ( .A(n_134), .Y(n_246) );
INVx1_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_135), .Y(n_145) );
INVx3_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g242 ( .A(n_135), .Y(n_242) );
BUFx3_ASAP7_75t_L g150 ( .A(n_136), .Y(n_150) );
INVx4_ASAP7_75t_SL g181 ( .A(n_136), .Y(n_181) );
INVx5_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx3_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_148), .Y(n_142) );
INVx2_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_147), .A2(n_191), .B(n_192), .C(n_193), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_147), .A2(n_193), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_147), .A2(n_478), .B(n_479), .C(n_480), .Y(n_477) );
O2A1O1Ixp5_ASAP7_75t_L g503 ( .A1(n_147), .A2(n_480), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_148), .A2(n_173), .B(n_455), .C(n_456), .Y(n_454) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_149), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_152), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g160 ( .A(n_153), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_153), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_153), .A2(n_217), .B(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_153), .A2(n_252), .B(n_452), .C(n_453), .Y(n_451) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_153), .A2(n_488), .B(n_495), .Y(n_487) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_L g166 ( .A(n_154), .B(n_155), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_160), .A2(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g284 ( .A(n_161), .B(n_184), .Y(n_284) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_161), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_161), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g374 ( .A(n_161), .Y(n_374) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g262 ( .A(n_162), .B(n_199), .Y(n_262) );
AND2x2_ASAP7_75t_L g289 ( .A(n_162), .B(n_200), .Y(n_289) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_167), .B(n_182), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_164), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_164), .A2(n_201), .B(n_211), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_164), .B(n_212), .Y(n_211) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_164), .A2(n_250), .B(n_257), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_164), .B(n_458), .Y(n_457) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_164), .A2(n_474), .B(n_481), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_164), .B(n_507), .Y(n_506) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_165), .A2(n_238), .B(n_239), .Y(n_237) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g259 ( .A(n_166), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_170), .B(n_171), .C(n_181), .Y(n_168) );
INVx2_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_170), .A2(n_181), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_170), .A2(n_181), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g489 ( .A1(n_170), .A2(n_181), .B(n_490), .C(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_170), .A2(n_181), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_170), .A2(n_181), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g541 ( .A1(n_170), .A2(n_181), .B(n_542), .C(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_173), .B(n_232), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g468 ( .A1(n_173), .A2(n_206), .B1(n_469), .B2(n_470), .Y(n_468) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_174), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_177), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g492 ( .A(n_178), .Y(n_492) );
INVx2_ASAP7_75t_L g480 ( .A(n_179), .Y(n_480) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_180), .Y(n_193) );
INVx1_ASAP7_75t_L g516 ( .A(n_180), .Y(n_516) );
INVx1_ASAP7_75t_L g194 ( .A(n_181), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_183), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_197), .Y(n_183) );
OR2x2_ASAP7_75t_L g315 ( .A(n_184), .B(n_198), .Y(n_315) );
AND2x2_ASAP7_75t_L g352 ( .A(n_184), .B(n_262), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_184), .B(n_283), .Y(n_363) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_184), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_184), .B(n_319), .Y(n_436) );
INVx5_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g261 ( .A(n_185), .Y(n_261) );
AND2x2_ASAP7_75t_L g270 ( .A(n_185), .B(n_198), .Y(n_270) );
AND2x2_ASAP7_75t_L g386 ( .A(n_185), .B(n_281), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_185), .B(n_319), .Y(n_408) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_195), .Y(n_185) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_198), .Y(n_354) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_199), .Y(n_306) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_L g283 ( .A(n_200), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_210), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .C(n_208), .Y(n_203) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_206), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_206), .B(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g533 ( .A(n_209), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_223), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_214), .B(n_296), .Y(n_415) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_215), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g267 ( .A(n_215), .B(n_268), .Y(n_267) );
INVx5_ASAP7_75t_SL g275 ( .A(n_215), .Y(n_275) );
OR2x2_ASAP7_75t_L g298 ( .A(n_215), .B(n_268), .Y(n_298) );
OR2x2_ASAP7_75t_L g308 ( .A(n_215), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g371 ( .A(n_215), .B(n_225), .Y(n_371) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_215), .B(n_224), .Y(n_409) );
NOR4xp25_ASAP7_75t_L g430 ( .A(n_215), .B(n_351), .C(n_431), .D(n_432), .Y(n_430) );
AND2x2_ASAP7_75t_L g440 ( .A(n_215), .B(n_272), .Y(n_440) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g265 ( .A(n_224), .B(n_261), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_224), .B(n_267), .Y(n_434) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_234), .Y(n_224) );
OR2x2_ASAP7_75t_L g274 ( .A(n_225), .B(n_275), .Y(n_274) );
INVx3_ASAP7_75t_L g281 ( .A(n_225), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_225), .B(n_249), .Y(n_293) );
INVxp67_ASAP7_75t_L g296 ( .A(n_225), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_225), .B(n_268), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_225), .B(n_235), .Y(n_362) );
AND2x2_ASAP7_75t_L g377 ( .A(n_225), .B(n_272), .Y(n_377) );
OR2x2_ASAP7_75t_L g406 ( .A(n_225), .B(n_235), .Y(n_406) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_233), .Y(n_225) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_226), .A2(n_510), .B(n_517), .Y(n_509) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_226), .A2(n_527), .B(n_534), .Y(n_526) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_226), .A2(n_540), .B(n_546), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_234), .B(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_234), .B(n_275), .Y(n_414) );
OR2x2_ASAP7_75t_L g435 ( .A(n_234), .B(n_312), .Y(n_435) );
INVx1_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g248 ( .A(n_235), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g272 ( .A(n_235), .B(n_268), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_235), .B(n_249), .Y(n_287) );
AND2x2_ASAP7_75t_L g357 ( .A(n_235), .B(n_281), .Y(n_357) );
AND2x2_ASAP7_75t_L g391 ( .A(n_235), .B(n_275), .Y(n_391) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_236), .B(n_275), .Y(n_294) );
AND2x2_ASAP7_75t_L g322 ( .A(n_236), .B(n_249), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_243), .B(n_244), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_244), .A2(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_247), .B(n_330), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_248), .A2(n_337), .B1(n_373), .B2(n_390), .C(n_392), .Y(n_389) );
INVx5_ASAP7_75t_SL g268 ( .A(n_249), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_253), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_252), .A2(n_475), .B(n_476), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_252), .A2(n_501), .B(n_502), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g463 ( .A(n_259), .Y(n_463) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OAI33xp33_ASAP7_75t_L g288 ( .A1(n_261), .A2(n_289), .A3(n_290), .B1(n_292), .B2(n_295), .B3(n_299), .Y(n_288) );
OR2x2_ASAP7_75t_L g304 ( .A(n_261), .B(n_305), .Y(n_304) );
AOI322xp5_ASAP7_75t_L g413 ( .A1(n_261), .A2(n_330), .A3(n_337), .B1(n_414), .B2(n_415), .C1(n_416), .C2(n_419), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_261), .B(n_289), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_SL g437 ( .A1(n_261), .A2(n_289), .B(n_438), .C(n_440), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_262), .A2(n_277), .B1(n_282), .B2(n_285), .C(n_288), .Y(n_276) );
INVx1_ASAP7_75t_L g369 ( .A(n_262), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_262), .B(n_418), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_266), .B1(n_269), .B2(n_271), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g346 ( .A(n_267), .B(n_281), .Y(n_346) );
AND2x2_ASAP7_75t_L g404 ( .A(n_267), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g312 ( .A(n_268), .B(n_275), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_268), .B(n_281), .Y(n_340) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_270), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_270), .B(n_348), .Y(n_402) );
OAI321xp33_ASAP7_75t_L g421 ( .A1(n_270), .A2(n_343), .A3(n_422), .B1(n_423), .B2(n_424), .C(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g388 ( .A(n_271), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_272), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g327 ( .A(n_272), .B(n_275), .Y(n_327) );
AOI321xp33_ASAP7_75t_L g385 ( .A1(n_272), .A2(n_289), .A3(n_386), .B1(n_387), .B2(n_388), .C(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g302 ( .A(n_274), .B(n_287), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_275), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_275), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_275), .B(n_361), .Y(n_398) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g321 ( .A(n_279), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g286 ( .A(n_280), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g394 ( .A(n_281), .Y(n_394) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_284), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g317 ( .A(n_289), .Y(n_317) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_291), .B(n_326), .Y(n_375) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OR2x2_ASAP7_75t_L g339 ( .A(n_294), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g384 ( .A(n_294), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_295), .A2(n_342), .B1(n_345), .B2(n_347), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g439 ( .A(n_298), .B(n_362), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B1(n_307), .B2(n_313), .C(n_316), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g337 ( .A(n_306), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_SL g383 ( .A(n_309), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_311), .B(n_361), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_311), .A2(n_379), .B(n_381), .Y(n_378) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g424 ( .A(n_312), .B(n_406), .Y(n_424) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_SL g326 ( .A(n_315), .Y(n_326) );
AOI21xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B(n_320), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g370 ( .A(n_322), .B(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g432 ( .A(n_322), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B(n_328), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_326), .B(n_344), .Y(n_380) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g401 ( .A(n_330), .Y(n_401) );
NAND5xp2_ASAP7_75t_L g331 ( .A(n_332), .B(n_349), .C(n_358), .D(n_378), .E(n_385), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_338), .C(n_341), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g373 ( .A(n_337), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_345), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_353), .B(n_355), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_350), .A2(n_404), .B1(n_407), .B2(n_409), .C(n_410), .Y(n_403) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AOI321xp33_ASAP7_75t_L g358 ( .A1(n_351), .A2(n_359), .A3(n_363), .B1(n_364), .B2(n_370), .C(n_372), .Y(n_358) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g429 ( .A(n_363), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_365), .B(n_369), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g381 ( .A(n_366), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NOR2xp67_ASAP7_75t_SL g393 ( .A(n_367), .B(n_374), .Y(n_393) );
AOI321xp33_ASAP7_75t_SL g425 ( .A1(n_370), .A2(n_426), .A3(n_427), .B1(n_428), .B2(n_429), .C(n_430), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B(n_375), .C(n_376), .Y(n_372) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_383), .B(n_391), .Y(n_420) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .C(n_395), .Y(n_392) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_421), .C(n_433), .Y(n_396) );
OAI211xp5_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_399), .B(n_403), .C(n_413), .Y(n_397) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_402), .A2(n_434), .B1(n_435), .B2(n_436), .C(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g422 ( .A(n_404), .Y(n_422) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g426 ( .A(n_424), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
CKINVDCx14_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g727 ( .A(n_442), .Y(n_727) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g726 ( .A(n_445), .Y(n_726) );
OR4x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_615), .C(n_662), .D(n_702), .Y(n_445) );
NAND3xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_561), .C(n_590), .Y(n_446) );
AOI211xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_483), .B(n_518), .C(n_554), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_448), .A2(n_574), .B(n_591), .C(n_595), .Y(n_590) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_459), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_450), .B(n_553), .Y(n_552) );
INVx3_ASAP7_75t_SL g557 ( .A(n_450), .Y(n_557) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_450), .Y(n_569) );
AND2x4_ASAP7_75t_L g573 ( .A(n_450), .B(n_525), .Y(n_573) );
AND2x2_ASAP7_75t_L g584 ( .A(n_450), .B(n_473), .Y(n_584) );
OR2x2_ASAP7_75t_L g608 ( .A(n_450), .B(n_521), .Y(n_608) );
AND2x2_ASAP7_75t_L g621 ( .A(n_450), .B(n_526), .Y(n_621) );
AND2x2_ASAP7_75t_L g661 ( .A(n_450), .B(n_647), .Y(n_661) );
AND2x2_ASAP7_75t_L g668 ( .A(n_450), .B(n_631), .Y(n_668) );
AND2x2_ASAP7_75t_L g698 ( .A(n_450), .B(n_460), .Y(n_698) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_457), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_459), .B(n_625), .Y(n_637) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_472), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_460), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g575 ( .A(n_460), .B(n_472), .Y(n_575) );
BUFx3_ASAP7_75t_L g583 ( .A(n_460), .Y(n_583) );
OR2x2_ASAP7_75t_L g604 ( .A(n_460), .B(n_486), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_460), .B(n_625), .Y(n_715) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_464), .B(n_471), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_462), .A2(n_522), .B(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g522 ( .A(n_464), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_471), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_472), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g568 ( .A(n_472), .Y(n_568) );
AND2x2_ASAP7_75t_L g631 ( .A(n_472), .B(n_526), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_472), .A2(n_634), .B1(n_636), .B2(n_638), .C(n_639), .Y(n_633) );
AND2x2_ASAP7_75t_L g647 ( .A(n_472), .B(n_521), .Y(n_647) );
AND2x2_ASAP7_75t_L g673 ( .A(n_472), .B(n_557), .Y(n_673) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g553 ( .A(n_473), .B(n_526), .Y(n_553) );
BUFx2_ASAP7_75t_L g687 ( .A(n_473), .Y(n_687) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI32xp33_ASAP7_75t_L g653 ( .A1(n_484), .A2(n_614), .A3(n_628), .B1(n_654), .B2(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_496), .Y(n_484) );
AND2x2_ASAP7_75t_L g594 ( .A(n_485), .B(n_538), .Y(n_594) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g576 ( .A(n_486), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_486), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g648 ( .A(n_486), .B(n_538), .Y(n_648) );
AND2x2_ASAP7_75t_L g659 ( .A(n_486), .B(n_551), .Y(n_659) );
BUFx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g560 ( .A(n_487), .B(n_539), .Y(n_560) );
AND2x2_ASAP7_75t_L g564 ( .A(n_487), .B(n_539), .Y(n_564) );
AND2x2_ASAP7_75t_L g599 ( .A(n_487), .B(n_550), .Y(n_599) );
AND2x2_ASAP7_75t_L g606 ( .A(n_487), .B(n_508), .Y(n_606) );
OAI211xp5_ASAP7_75t_L g611 ( .A1(n_487), .A2(n_557), .B(n_568), .C(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g665 ( .A(n_487), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_487), .B(n_498), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_496), .B(n_548), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_496), .B(n_564), .Y(n_654) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g559 ( .A(n_497), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_508), .Y(n_497) );
AND2x2_ASAP7_75t_L g551 ( .A(n_498), .B(n_509), .Y(n_551) );
OR2x2_ASAP7_75t_L g566 ( .A(n_498), .B(n_509), .Y(n_566) );
AND2x2_ASAP7_75t_L g589 ( .A(n_498), .B(n_550), .Y(n_589) );
INVx1_ASAP7_75t_L g593 ( .A(n_498), .Y(n_593) );
AND2x2_ASAP7_75t_L g612 ( .A(n_498), .B(n_549), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_498), .A2(n_577), .B1(n_623), .B2(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_498), .B(n_665), .Y(n_689) );
AND2x2_ASAP7_75t_L g704 ( .A(n_498), .B(n_564), .Y(n_704) );
INVx4_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx3_ASAP7_75t_L g536 ( .A(n_499), .Y(n_536) );
AND2x2_ASAP7_75t_L g578 ( .A(n_499), .B(n_509), .Y(n_578) );
AND2x2_ASAP7_75t_L g580 ( .A(n_499), .B(n_538), .Y(n_580) );
AND3x2_ASAP7_75t_L g642 ( .A(n_499), .B(n_606), .C(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g677 ( .A(n_508), .B(n_549), .Y(n_677) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g538 ( .A(n_509), .B(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_509), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_509), .B(n_548), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g717 ( .A(n_509), .B(n_589), .C(n_665), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_535), .B1(n_547), .B2(n_552), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_524), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_521), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g629 ( .A(n_521), .Y(n_629) );
OAI31xp33_ASAP7_75t_L g645 ( .A1(n_524), .A2(n_646), .A3(n_647), .B(n_648), .Y(n_645) );
AND2x2_ASAP7_75t_L g670 ( .A(n_524), .B(n_557), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_524), .B(n_583), .Y(n_716) );
AND2x2_ASAP7_75t_L g625 ( .A(n_525), .B(n_557), .Y(n_625) );
AND2x2_ASAP7_75t_L g686 ( .A(n_525), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g556 ( .A(n_526), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g614 ( .A(n_526), .Y(n_614) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g635 ( .A(n_536), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_537), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AOI221x1_ASAP7_75t_SL g602 ( .A1(n_538), .A2(n_603), .B1(n_605), .B2(n_607), .C(n_609), .Y(n_602) );
INVx2_ASAP7_75t_L g550 ( .A(n_539), .Y(n_550) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_539), .Y(n_644) );
INVx1_ASAP7_75t_L g632 ( .A(n_547), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_548), .B(n_565), .Y(n_657) );
INVx1_ASAP7_75t_SL g720 ( .A(n_548), .Y(n_720) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g638 ( .A(n_551), .B(n_564), .Y(n_638) );
INVx1_ASAP7_75t_L g706 ( .A(n_552), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_552), .B(n_635), .Y(n_719) );
INVx2_ASAP7_75t_SL g558 ( .A(n_553), .Y(n_558) );
AND2x2_ASAP7_75t_L g601 ( .A(n_553), .B(n_557), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_553), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_553), .B(n_628), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_558), .B(n_559), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_556), .B(n_628), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_556), .B(n_583), .Y(n_724) );
OR2x2_ASAP7_75t_L g596 ( .A(n_557), .B(n_575), .Y(n_596) );
AND2x2_ASAP7_75t_L g695 ( .A(n_557), .B(n_686), .Y(n_695) );
OAI22xp5_ASAP7_75t_SL g570 ( .A1(n_558), .A2(n_571), .B1(n_576), .B2(n_579), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_558), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g618 ( .A(n_560), .B(n_566), .Y(n_618) );
INVx1_ASAP7_75t_L g682 ( .A(n_560), .Y(n_682) );
AOI311xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_567), .A3(n_569), .B(n_570), .C(n_581), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_565), .A2(n_697), .B1(n_709), .B2(n_712), .C(n_714), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_565), .B(n_720), .Y(n_722) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g619 ( .A(n_567), .Y(n_619) );
AOI211xp5_ASAP7_75t_L g609 ( .A1(n_568), .A2(n_610), .B(n_611), .C(n_613), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_SL g678 ( .A1(n_572), .A2(n_574), .B(n_679), .C(n_680), .Y(n_678) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_573), .B(n_647), .Y(n_713) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_576), .A2(n_596), .B1(n_597), .B2(n_600), .C(n_602), .Y(n_595) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g598 ( .A(n_578), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g681 ( .A(n_578), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_582), .A2(n_640), .B(n_641), .C(n_645), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_583), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_583), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g605 ( .A(n_589), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_593), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g707 ( .A(n_596), .Y(n_707) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_599), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g634 ( .A(n_599), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g711 ( .A(n_599), .Y(n_711) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g652 ( .A(n_601), .B(n_628), .Y(n_652) );
INVx1_ASAP7_75t_SL g646 ( .A(n_608), .Y(n_646) );
INVx1_ASAP7_75t_L g623 ( .A(n_614), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g615 ( .A(n_616), .B(n_633), .C(n_649), .Y(n_615) );
AOI322xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .A3(n_620), .B1(n_622), .B2(n_626), .C1(n_630), .C2(n_632), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_617), .A2(n_670), .B(n_671), .C(n_678), .Y(n_669) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_620), .A2(n_641), .B1(n_672), .B2(n_674), .Y(n_671) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g630 ( .A(n_628), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g667 ( .A(n_628), .B(n_668), .Y(n_667) );
AOI32xp33_ASAP7_75t_L g718 ( .A1(n_628), .A2(n_719), .A3(n_720), .B1(n_721), .B2(n_723), .Y(n_718) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g640 ( .A(n_631), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_631), .A2(n_684), .B1(n_688), .B2(n_690), .C(n_693), .Y(n_683) );
AND2x2_ASAP7_75t_L g697 ( .A(n_631), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g700 ( .A(n_635), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g710 ( .A(n_635), .B(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g701 ( .A(n_644), .B(n_665), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B(n_653), .C(n_656), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI21xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B(n_660), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_666), .B(n_669), .C(n_683), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_677), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g692 ( .A(n_689), .Y(n_692) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B(n_699), .Y(n_693) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI211xp5_ASAP7_75t_SL g702 ( .A1(n_703), .A2(n_705), .B(n_708), .C(n_718), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OAI21xp5_ASAP7_75t_SL g737 ( .A1(n_738), .A2(n_741), .B(n_743), .Y(n_737) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
endmodule