module fake_jpeg_23476_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_8),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_30),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_42),
.Y(n_82)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_29),
.B1(n_24),
.B2(n_20),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_36),
.B1(n_27),
.B2(n_16),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_75),
.B1(n_79),
.B2(n_83),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_27),
.B1(n_25),
.B2(n_16),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_93),
.B1(n_31),
.B2(n_35),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_25),
.B1(n_16),
.B2(n_29),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_0),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_24),
.B1(n_29),
.B2(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_42),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_88),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_49),
.B(n_20),
.CI(n_31),
.CON(n_88),
.SN(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_24),
.B1(n_26),
.B2(n_20),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_26),
.B1(n_20),
.B2(n_25),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_22),
.B1(n_17),
.B2(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_31),
.B1(n_25),
.B2(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_56),
.B(n_34),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_94),
.B(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_97),
.A2(n_98),
.B1(n_118),
.B2(n_70),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_112),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_71),
.B1(n_78),
.B2(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_108),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_102),
.Y(n_143)
);

OR2x4_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_32),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_88),
.B(n_74),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_19),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_68),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_110),
.Y(n_148)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_17),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_118),
.Y(n_124)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_40),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_121),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_22),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_76),
.B(n_19),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_123),
.Y(n_145)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_78),
.B1(n_87),
.B2(n_74),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_91),
.C(n_77),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_149),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_73),
.B(n_51),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_139),
.B(n_122),
.Y(n_152)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_141),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_97),
.B1(n_112),
.B2(n_117),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_58),
.B(n_88),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_71),
.B1(n_72),
.B2(n_95),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_146),
.B1(n_107),
.B2(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_77),
.C(n_95),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_37),
.B(n_40),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_102),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_150),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_152),
.A2(n_131),
.B(n_137),
.Y(n_203)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_161),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_170),
.B1(n_144),
.B2(n_134),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_158),
.A2(n_165),
.B1(n_174),
.B2(n_135),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_121),
.A3(n_107),
.B1(n_115),
.B2(n_101),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_145),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_125),
.A2(n_111),
.B1(n_81),
.B2(n_99),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_32),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_128),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_61),
.C(n_41),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_128),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_87),
.B1(n_92),
.B2(n_22),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_105),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_105),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_81),
.B1(n_99),
.B2(n_87),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_81),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_176),
.B(n_125),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_133),
.C(n_130),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_179),
.C(n_188),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_136),
.B1(n_133),
.B2(n_148),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_190),
.B1(n_194),
.B2(n_154),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_150),
.C(n_143),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_198),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_143),
.C(n_141),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_163),
.A2(n_148),
.B1(n_140),
.B2(n_147),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_166),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_144),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_144),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_197),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_137),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_174),
.B1(n_160),
.B2(n_168),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_11),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_172),
.B(n_131),
.Y(n_213)
);

NAND2x1_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_169),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_207),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_156),
.CI(n_159),
.CON(n_206),
.SN(n_206)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_217),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_183),
.A2(n_164),
.B(n_151),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_216),
.B(n_23),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_194),
.B1(n_184),
.B2(n_180),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_218),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_170),
.B1(n_168),
.B2(n_135),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_193),
.A2(n_167),
.B(n_52),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_92),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_201),
.B1(n_185),
.B2(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_15),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_219),
.B(n_12),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_52),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_227),
.C(n_192),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_69),
.B1(n_67),
.B2(n_65),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_185),
.A2(n_54),
.B1(n_50),
.B2(n_61),
.Y(n_222)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_186),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_54),
.C(n_50),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_12),
.Y(n_243)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_233),
.C(n_215),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_192),
.C(n_201),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_235),
.A2(n_241),
.B(n_245),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

AO22x1_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_180),
.B1(n_195),
.B2(n_198),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_216),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_224),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_247),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_33),
.B1(n_28),
.B2(n_21),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_32),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_225),
.B1(n_229),
.B2(n_226),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_212),
.B1(n_227),
.B2(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_258),
.C(n_263),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_232),
.C(n_230),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_207),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_204),
.C(n_220),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_204),
.C(n_206),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_265),
.C(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_206),
.C(n_209),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_241),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_239),
.C(n_236),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_212),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_0),
.C(n_1),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_249),
.B1(n_231),
.B2(n_234),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_282),
.B1(n_2),
.B2(n_3),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_235),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_267),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_254),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_285),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_231),
.B1(n_234),
.B2(n_250),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_248),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_286),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_0),
.C(n_1),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_259),
.C(n_253),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_33),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_287),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_33),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_10),
.B(n_15),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_264),
.B1(n_257),
.B2(n_263),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_296),
.B1(n_21),
.B2(n_28),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_261),
.C(n_252),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_303),
.C(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

OAI321xp33_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_33),
.A3(n_28),
.B1(n_21),
.B2(n_18),
.C(n_7),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_301),
.B1(n_302),
.B2(n_7),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_23),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_3),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_277),
.A2(n_9),
.B1(n_10),
.B2(n_7),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_277),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_3),
.C(n_4),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_302),
.B(n_289),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_310),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_272),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_306),
.B(n_313),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_294),
.B(n_5),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_314),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_272),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_18),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_298),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_303),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_4),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_318),
.C(n_320),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_5),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_311),
.B(n_314),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_294),
.B1(n_21),
.B2(n_18),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_324),
.Y(n_326)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_327),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_6),
.C(n_18),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_322),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_23),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_23),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

AO21x2_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_326),
.B(n_334),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_333),
.B(n_28),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_333),
.C(n_6),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_6),
.C(n_337),
.Y(n_341)
);


endmodule