module fake_netlist_6_2090_n_2903 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2903);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2903;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_1371;
wire n_873;
wire n_1285;
wire n_2886;
wire n_1985;
wire n_2838;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2345;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_928;
wire n_1214;
wire n_835;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_627;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2307;
wire n_2069;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2900;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_1548;
wire n_799;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2888;
wire n_2793;
wire n_2715;
wire n_2885;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_1583;
wire n_832;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_771;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_2899;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_SL g625 ( 
.A(n_27),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_343),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_12),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_221),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_339),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_271),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_381),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_572),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_249),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_151),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_471),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_318),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_308),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_140),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_456),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_436),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_568),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_414),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_547),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_204),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_600),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_416),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_480),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_92),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_158),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_304),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_288),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_183),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_242),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_293),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_542),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_567),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_260),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_315),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_100),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_535),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_339),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_556),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_531),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_375),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_516),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_219),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_451),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_205),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_311),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_292),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_5),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_105),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_96),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_325),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_354),
.Y(n_675)
);

BUFx2_ASAP7_75t_SL g676 ( 
.A(n_491),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_458),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_125),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_574),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_172),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_573),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_115),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_462),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_319),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_393),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_342),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_91),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_313),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_41),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_566),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_28),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_120),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_343),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_576),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_183),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_581),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_319),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_451),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_46),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_162),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_162),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_148),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_308),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_601),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_538),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_1),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_466),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_582),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_88),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_257),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_617),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_571),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_37),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_565),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_543),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_46),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_583),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_598),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_219),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_258),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_220),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_298),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_205),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_226),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_580),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_449),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_493),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_53),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_267),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_405),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_518),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_55),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_250),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_483),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_352),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_523),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_564),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_215),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_459),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_192),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_359),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_163),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_116),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_4),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_555),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_575),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_376),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_473),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_375),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_606),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_600),
.Y(n_751)
);

BUFx10_ASAP7_75t_L g752 ( 
.A(n_570),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_73),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_279),
.Y(n_754)
);

CKINVDCx14_ASAP7_75t_R g755 ( 
.A(n_450),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_116),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_246),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_583),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_192),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_337),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_347),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_587),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_56),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_464),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_448),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_428),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_6),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_226),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_352),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_577),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_310),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_468),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_324),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_556),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_549),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_590),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_403),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_63),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_519),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_202),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_588),
.Y(n_781)
);

CKINVDCx16_ASAP7_75t_R g782 ( 
.A(n_133),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_24),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_223),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_521),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_286),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_258),
.Y(n_787)
);

BUFx10_ASAP7_75t_L g788 ( 
.A(n_113),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_562),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_599),
.Y(n_790)
);

CKINVDCx14_ASAP7_75t_R g791 ( 
.A(n_80),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_201),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_550),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_156),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_350),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_442),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_9),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_309),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_578),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_215),
.Y(n_800)
);

CKINVDCx16_ASAP7_75t_R g801 ( 
.A(n_214),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_107),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_576),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_260),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_298),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_441),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_331),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_182),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_578),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_299),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_127),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_579),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_23),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_245),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_20),
.Y(n_815)
);

BUFx10_ASAP7_75t_L g816 ( 
.A(n_623),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_186),
.Y(n_817)
);

BUFx10_ASAP7_75t_L g818 ( 
.A(n_315),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_409),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_466),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_55),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_75),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_259),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_64),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_178),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_185),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_142),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_124),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_273),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_172),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_134),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_233),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_347),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_587),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_379),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_208),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_146),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_98),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_541),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_149),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_563),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_422),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_406),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_98),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_22),
.Y(n_845)
);

BUFx10_ASAP7_75t_L g846 ( 
.A(n_479),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_401),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_394),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_588),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_238),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_552),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_104),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_474),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_248),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_558),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_395),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_28),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_462),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_198),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_357),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_387),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_622),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_23),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_360),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_373),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_301),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_22),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_569),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_489),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_25),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_565),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_124),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_563),
.Y(n_873)
);

INVxp33_ASAP7_75t_SL g874 ( 
.A(n_764),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_755),
.Y(n_875)
);

CKINVDCx16_ASAP7_75t_R g876 ( 
.A(n_782),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_670),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_791),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_802),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_670),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_708),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_708),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_737),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_737),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_796),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_796),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_820),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_820),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_801),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_833),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_833),
.Y(n_891)
);

CKINVDCx16_ASAP7_75t_R g892 ( 
.A(n_643),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_847),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_847),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_666),
.Y(n_895)
);

CKINVDCx14_ASAP7_75t_R g896 ( 
.A(n_775),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_853),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_674),
.Y(n_898)
);

INVxp33_ASAP7_75t_SL g899 ( 
.A(n_626),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_674),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_674),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_853),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_674),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_641),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_850),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_667),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_674),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_663),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_790),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_790),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_790),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_790),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_673),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_790),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_668),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_671),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_844),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_844),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_643),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_844),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_844),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_844),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_816),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_848),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_848),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_675),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_643),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_848),
.Y(n_928)
);

INVxp33_ASAP7_75t_SL g929 ( 
.A(n_626),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_848),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_652),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_848),
.Y(n_932)
);

CKINVDCx16_ASAP7_75t_R g933 ( 
.A(n_652),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_677),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_679),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_680),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_687),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_627),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_750),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_628),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_630),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_629),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_713),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_640),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_632),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_636),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_637),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_681),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_638),
.Y(n_949)
);

INVxp33_ASAP7_75t_L g950 ( 
.A(n_639),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_640),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_645),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_646),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_630),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_685),
.Y(n_955)
);

INVxp33_ASAP7_75t_L g956 ( 
.A(n_650),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_656),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_657),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_652),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_686),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_664),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_688),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_669),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_720),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_672),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_678),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_689),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_711),
.B(n_0),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_725),
.Y(n_969)
);

INVxp33_ASAP7_75t_L g970 ( 
.A(n_682),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_684),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_691),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_695),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_697),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_741),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_910),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_923),
.B(n_862),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_910),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_910),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_904),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_910),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_923),
.B(n_862),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_928),
.Y(n_983)
);

BUFx12f_ASAP7_75t_L g984 ( 
.A(n_875),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_875),
.B(n_816),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_877),
.B(n_683),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_927),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_941),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_880),
.B(n_683),
.Y(n_989)
);

CKINVDCx6p67_ASAP7_75t_R g990 ( 
.A(n_876),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_881),
.B(n_701),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_898),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_878),
.B(n_816),
.Y(n_993)
);

INVx5_ASAP7_75t_L g994 ( 
.A(n_928),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_939),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_927),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_898),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_928),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_882),
.B(n_701),
.Y(n_999)
);

BUFx8_ASAP7_75t_SL g1000 ( 
.A(n_904),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_889),
.Y(n_1001)
);

BUFx12f_ASAP7_75t_L g1002 ( 
.A(n_878),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_939),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_898),
.B(n_653),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_903),
.B(n_653),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_883),
.B(n_733),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_928),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_900),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_903),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_889),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_900),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_901),
.Y(n_1012)
);

INVx5_ASAP7_75t_L g1013 ( 
.A(n_903),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_884),
.B(n_860),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_885),
.B(n_733),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_901),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_886),
.B(n_759),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_939),
.Y(n_1018)
);

BUFx12f_ASAP7_75t_L g1019 ( 
.A(n_895),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_887),
.B(n_759),
.Y(n_1020)
);

AND2x6_ASAP7_75t_L g1021 ( 
.A(n_925),
.B(n_730),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_925),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_939),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_907),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_968),
.B(n_895),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_909),
.B(n_730),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_911),
.Y(n_1027)
);

INVx5_ASAP7_75t_L g1028 ( 
.A(n_944),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_888),
.B(n_890),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_944),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_891),
.B(n_784),
.Y(n_1031)
);

CKINVDCx6p67_ASAP7_75t_R g1032 ( 
.A(n_892),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_912),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_906),
.B(n_915),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_893),
.B(n_784),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_944),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_954),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_894),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_951),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_914),
.Y(n_1040)
);

INVx5_ASAP7_75t_L g1041 ( 
.A(n_951),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1009),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_987),
.B(n_905),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1014),
.B(n_897),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1009),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1009),
.B(n_917),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1005),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_1008),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1012),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1014),
.B(n_902),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_1038),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1005),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_987),
.B(n_879),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1030),
.B(n_918),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1005),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1005),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_992),
.B(n_920),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_976),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1012),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1024),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1024),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_976),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_976),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1030),
.B(n_921),
.Y(n_1064)
);

AND2x6_ASAP7_75t_L g1065 ( 
.A(n_1025),
.B(n_747),
.Y(n_1065)
);

AND2x6_ASAP7_75t_L g1066 ( 
.A(n_1004),
.B(n_747),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1004),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1004),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_L g1069 ( 
.A(n_988),
.B(n_1037),
.C(n_724),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1040),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_992),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1040),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_996),
.B(n_933),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1016),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1016),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_997),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_976),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_1008),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_997),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1026),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_996),
.B(n_906),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1038),
.B(n_1026),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1026),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1026),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_976),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1030),
.B(n_922),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_979),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_979),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_998),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1008),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_978),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_986),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_998),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1008),
.Y(n_1094)
);

AND3x2_ASAP7_75t_L g1095 ( 
.A(n_1001),
.B(n_931),
.C(n_919),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_1018),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1008),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1007),
.Y(n_1098)
);

INVxp33_ASAP7_75t_SL g1099 ( 
.A(n_985),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1007),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_989),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_977),
.B(n_899),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_983),
.B(n_924),
.Y(n_1103)
);

AND3x2_ASAP7_75t_L g1104 ( 
.A(n_1001),
.B(n_959),
.C(n_757),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1011),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_991),
.B(n_930),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1011),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_983),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1023),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1011),
.B(n_932),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1023),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1023),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1011),
.B(n_938),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1011),
.B(n_1022),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1022),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1022),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1023),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1022),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_999),
.B(n_940),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1023),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1022),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1027),
.Y(n_1122)
);

CKINVDCx8_ASAP7_75t_R g1123 ( 
.A(n_1010),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_978),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_978),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1006),
.B(n_942),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1027),
.Y(n_1127)
);

OA21x2_ASAP7_75t_L g1128 ( 
.A1(n_1015),
.A2(n_1020),
.B(n_1017),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1027),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1027),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_982),
.A2(n_946),
.B(n_945),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1066),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1082),
.Y(n_1133)
);

INVx6_ASAP7_75t_L g1134 ( 
.A(n_1057),
.Y(n_1134)
);

OAI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1092),
.A2(n_915),
.B1(n_926),
.B2(n_916),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1074),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1074),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1047),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1047),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1074),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1052),
.B(n_1034),
.C(n_1031),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1075),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1052),
.Y(n_1143)
);

NOR2x1p5_ASAP7_75t_L g1144 ( 
.A(n_1043),
.B(n_1032),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1065),
.B(n_993),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1102),
.B(n_1010),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1075),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1075),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1055),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1049),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_L g1151 ( 
.A(n_1073),
.B(n_1081),
.C(n_1069),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1082),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1049),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_1131),
.A2(n_1035),
.B(n_710),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1049),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1059),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1053),
.B(n_916),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1051),
.Y(n_1158)
);

CKINVDCx6p67_ASAP7_75t_R g1159 ( 
.A(n_1043),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1066),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1065),
.B(n_1055),
.Y(n_1161)
);

NOR2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1053),
.B(n_1032),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_1066),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1059),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1099),
.B(n_899),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1059),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1056),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1065),
.B(n_1056),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1060),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1092),
.B(n_926),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1065),
.B(n_995),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1080),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1060),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1051),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1060),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1061),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1101),
.B(n_934),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1066),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1101),
.B(n_929),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_SL g1180 ( 
.A(n_1119),
.B(n_934),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1119),
.B(n_935),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1061),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1065),
.A2(n_874),
.B1(n_929),
.B2(n_1021),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1061),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1080),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1071),
.B(n_935),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1070),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1065),
.B(n_1083),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1042),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1126),
.B(n_1029),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1083),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1044),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1084),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1070),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1065),
.B(n_995),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1084),
.Y(n_1196)
);

BUFx10_ASAP7_75t_L g1197 ( 
.A(n_1095),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_L g1198 ( 
.A(n_1065),
.B(n_1021),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1071),
.B(n_936),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1126),
.B(n_936),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1044),
.B(n_948),
.Y(n_1201)
);

INVx5_ASAP7_75t_L g1202 ( 
.A(n_1066),
.Y(n_1202)
);

NOR2x1p5_ASAP7_75t_L g1203 ( 
.A(n_1050),
.B(n_990),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1128),
.B(n_955),
.C(n_948),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1070),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1072),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1072),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1103),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1103),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1072),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1050),
.B(n_955),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1067),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1042),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1045),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1045),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1057),
.Y(n_1216)
);

CKINVDCx16_ASAP7_75t_R g1217 ( 
.A(n_1123),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1087),
.Y(n_1218)
);

INVx8_ASAP7_75t_L g1219 ( 
.A(n_1066),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1067),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1076),
.B(n_960),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1068),
.A2(n_960),
.B1(n_967),
.B2(n_962),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1087),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1057),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1088),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1068),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1057),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1088),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1089),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1046),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1078),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1089),
.Y(n_1232)
);

INVx8_ASAP7_75t_L g1233 ( 
.A(n_1066),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1128),
.B(n_1106),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_L g1235 ( 
.A(n_1066),
.B(n_1021),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1046),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1106),
.B(n_896),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1093),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1093),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1108),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1058),
.Y(n_1241)
);

INVx11_ASAP7_75t_L g1242 ( 
.A(n_1123),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1076),
.B(n_962),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1098),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1128),
.B(n_995),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_1078),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1098),
.Y(n_1247)
);

AND2x2_ASAP7_75t_SL g1248 ( 
.A(n_1128),
.B(n_751),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1108),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1128),
.A2(n_874),
.B1(n_1021),
.B2(n_676),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1079),
.B(n_1100),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1100),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1058),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1079),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1123),
.B(n_967),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1110),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1131),
.B(n_1054),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1131),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1054),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1110),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1064),
.B(n_1003),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1064),
.B(n_1003),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1086),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1113),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1113),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1078),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1086),
.B(n_1003),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1109),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1090),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1109),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1165),
.B(n_908),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1241),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1213),
.Y(n_1273)
);

XNOR2x2_ASAP7_75t_L g1274 ( 
.A(n_1255),
.B(n_625),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1213),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1138),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1138),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1179),
.B(n_908),
.Y(n_1278)
);

XNOR2x2_ASAP7_75t_L g1279 ( 
.A(n_1146),
.B(n_660),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1139),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1139),
.Y(n_1281)
);

NAND2x1p5_ASAP7_75t_L g1282 ( 
.A(n_1163),
.B(n_1048),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1143),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1157),
.B(n_1019),
.Y(n_1284)
);

AND2x6_ASAP7_75t_L g1285 ( 
.A(n_1132),
.B(n_1090),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1143),
.Y(n_1286)
);

INVxp33_ASAP7_75t_L g1287 ( 
.A(n_1237),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1149),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1234),
.A2(n_1114),
.B(n_1094),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1158),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1149),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1190),
.B(n_1069),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1167),
.Y(n_1293)
);

XOR2xp5_ASAP7_75t_L g1294 ( 
.A(n_1217),
.B(n_980),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1158),
.B(n_990),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1167),
.Y(n_1296)
);

XOR2xp5_ASAP7_75t_L g1297 ( 
.A(n_1217),
.B(n_980),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1174),
.B(n_1019),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1214),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1212),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1212),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1242),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1220),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1220),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1190),
.B(n_984),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1237),
.B(n_1104),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1159),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1192),
.B(n_1104),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1226),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1226),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1172),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1214),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1192),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1174),
.B(n_984),
.Y(n_1314)
);

INVxp67_ASAP7_75t_SL g1315 ( 
.A(n_1241),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1172),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1185),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1241),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1185),
.Y(n_1319)
);

XOR2xp5_ASAP7_75t_L g1320 ( 
.A(n_1141),
.B(n_913),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1191),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1191),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1193),
.Y(n_1323)
);

INVxp33_ASAP7_75t_L g1324 ( 
.A(n_1170),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1264),
.B(n_1090),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1159),
.B(n_734),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1193),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1196),
.Y(n_1328)
);

AND2x6_ASAP7_75t_L g1329 ( 
.A(n_1132),
.B(n_1094),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1245),
.A2(n_1114),
.B(n_1097),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1264),
.B(n_1094),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1196),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1218),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1181),
.B(n_1002),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1218),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1133),
.B(n_1095),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1200),
.B(n_1002),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1189),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1177),
.B(n_1201),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1180),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1189),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1223),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1135),
.B(n_913),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1223),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1189),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1245),
.A2(n_1107),
.B(n_1097),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1225),
.Y(n_1347)
);

XOR2xp5_ASAP7_75t_L g1348 ( 
.A(n_1141),
.B(n_937),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1225),
.Y(n_1349)
);

INVxp33_ASAP7_75t_L g1350 ( 
.A(n_1211),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1186),
.B(n_937),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1215),
.Y(n_1352)
);

XNOR2xp5_ASAP7_75t_L g1353 ( 
.A(n_1162),
.B(n_943),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1228),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1228),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1229),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1229),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1232),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1232),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1238),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1133),
.B(n_943),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1238),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1215),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1239),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1239),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1244),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1244),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1222),
.B(n_964),
.Y(n_1368)
);

INVxp33_ASAP7_75t_L g1369 ( 
.A(n_1199),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1247),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1247),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1252),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1252),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1240),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1203),
.B(n_829),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1221),
.B(n_947),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1240),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1249),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1249),
.Y(n_1379)
);

INVxp67_ASAP7_75t_SL g1380 ( 
.A(n_1241),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1268),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1268),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1270),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1265),
.B(n_1097),
.Y(n_1384)
);

XOR2xp5_ASAP7_75t_L g1385 ( 
.A(n_1204),
.B(n_964),
.Y(n_1385)
);

XNOR2xp5_ASAP7_75t_L g1386 ( 
.A(n_1162),
.B(n_969),
.Y(n_1386)
);

XOR2xp5_ASAP7_75t_L g1387 ( 
.A(n_1204),
.B(n_969),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1265),
.B(n_1107),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1270),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1243),
.B(n_1152),
.Y(n_1390)
);

XNOR2xp5_ASAP7_75t_L g1391 ( 
.A(n_1144),
.B(n_975),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1241),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1152),
.B(n_975),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1215),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1136),
.Y(n_1395)
);

XNOR2x1_ASAP7_75t_L g1396 ( 
.A(n_1144),
.B(n_631),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1136),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1137),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1137),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1140),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1140),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1254),
.B(n_768),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1234),
.A2(n_1115),
.B(n_1107),
.Y(n_1403)
);

XOR2xp5_ASAP7_75t_L g1404 ( 
.A(n_1183),
.B(n_1000),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1142),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1254),
.B(n_1216),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1142),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1147),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1147),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_1251),
.B(n_1208),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1197),
.Y(n_1411)
);

XNOR2x2_ASAP7_75t_L g1412 ( 
.A(n_1242),
.B(n_736),
.Y(n_1412)
);

XNOR2x2_ASAP7_75t_L g1413 ( 
.A(n_1145),
.B(n_745),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1259),
.B(n_772),
.Y(n_1414)
);

XNOR2xp5_ASAP7_75t_L g1415 ( 
.A(n_1203),
.B(n_1000),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1148),
.Y(n_1416)
);

AND2x6_ASAP7_75t_L g1417 ( 
.A(n_1132),
.B(n_1115),
.Y(n_1417)
);

XOR2x2_ASAP7_75t_L g1418 ( 
.A(n_1151),
.B(n_761),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1148),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1197),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1197),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1224),
.Y(n_1422)
);

NAND2x1p5_ASAP7_75t_L g1423 ( 
.A(n_1163),
.B(n_1048),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1224),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1224),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1227),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1230),
.B(n_1115),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1230),
.B(n_1116),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1227),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1227),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1169),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1197),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1236),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1169),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1173),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1173),
.Y(n_1436)
);

NOR2xp67_ASAP7_75t_L g1437 ( 
.A(n_1208),
.B(n_949),
.Y(n_1437)
);

BUFx2_ASAP7_75t_R g1438 ( 
.A(n_1154),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1253),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1209),
.B(n_950),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1236),
.B(n_1116),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1259),
.B(n_797),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1175),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1263),
.B(n_808),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1263),
.B(n_1209),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1154),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1256),
.Y(n_1447)
);

XOR2xp5_ASAP7_75t_L g1448 ( 
.A(n_1132),
.B(n_815),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1216),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1175),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1176),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_SL g1452 ( 
.A(n_1163),
.B(n_834),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1176),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1256),
.B(n_956),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1260),
.B(n_826),
.Y(n_1455)
);

NAND2x1p5_ASAP7_75t_L g1456 ( 
.A(n_1163),
.B(n_1048),
.Y(n_1456)
);

XOR2xp5_ASAP7_75t_L g1457 ( 
.A(n_1132),
.B(n_830),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1260),
.B(n_856),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1182),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1182),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1248),
.B(n_1116),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1184),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1184),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1134),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1187),
.Y(n_1465)
);

XNOR2x2_ASAP7_75t_L g1466 ( 
.A(n_1257),
.B(n_778),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1187),
.Y(n_1467)
);

XOR2x2_ASAP7_75t_L g1468 ( 
.A(n_1250),
.B(n_795),
.Y(n_1468)
);

INVxp33_ASAP7_75t_L g1469 ( 
.A(n_1257),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1248),
.B(n_970),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1171),
.A2(n_1121),
.B(n_1118),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1194),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1194),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1369),
.B(n_1248),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1447),
.B(n_1202),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1273),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1445),
.B(n_1261),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1272),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1452),
.B(n_1202),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1393),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1445),
.B(n_1205),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1278),
.B(n_1134),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1276),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1461),
.A2(n_1171),
.B(n_1219),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1275),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1299),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1410),
.A2(n_1188),
.B(n_1161),
.C(n_1168),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1452),
.B(n_1202),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1442),
.B(n_1444),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_L g1490 ( 
.A(n_1271),
.B(n_692),
.C(n_690),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1433),
.B(n_1470),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1277),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1414),
.B(n_1134),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1406),
.B(n_1202),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1414),
.B(n_1458),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1454),
.B(n_1154),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1402),
.B(n_1134),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1406),
.B(n_1202),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1307),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1433),
.B(n_1205),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1461),
.A2(n_1233),
.B(n_1219),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1402),
.B(n_1455),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1312),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1372),
.B(n_1206),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1455),
.B(n_1262),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1280),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1440),
.B(n_735),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1287),
.A2(n_1160),
.B1(n_1233),
.B2(n_1219),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1438),
.A2(n_1160),
.B1(n_1178),
.B2(n_1219),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_1326),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1281),
.Y(n_1511)
);

INVx2_ASAP7_75t_SL g1512 ( 
.A(n_1290),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1390),
.B(n_1267),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1468),
.A2(n_1178),
.B1(n_1233),
.B2(n_1219),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1292),
.B(n_1202),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1376),
.B(n_1178),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1411),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1437),
.B(n_1313),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1313),
.B(n_1206),
.Y(n_1519)
);

NOR2xp67_ASAP7_75t_L g1520 ( 
.A(n_1298),
.B(n_1258),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1373),
.B(n_1207),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1300),
.B(n_1207),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1301),
.B(n_1210),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1466),
.A2(n_1413),
.B1(n_1274),
.B2(n_1418),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1303),
.B(n_1210),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1304),
.B(n_1150),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1283),
.B(n_1150),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1286),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1288),
.B(n_1153),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1298),
.B(n_1178),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1291),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1293),
.B(n_1153),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1296),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1272),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1401),
.Y(n_1535)
);

AND2x6_ASAP7_75t_L g1536 ( 
.A(n_1311),
.B(n_1178),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1316),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1317),
.B(n_1155),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1319),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1459),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1309),
.B(n_1155),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1272),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1321),
.B(n_1156),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1314),
.B(n_1233),
.Y(n_1544)
);

NAND2x1_ASAP7_75t_L g1545 ( 
.A(n_1285),
.B(n_1253),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1351),
.B(n_1266),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1322),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1432),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1361),
.B(n_857),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1323),
.B(n_1156),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1464),
.B(n_1233),
.Y(n_1551)
);

AOI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1346),
.A2(n_1195),
.B(n_1258),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1361),
.B(n_1339),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1290),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1295),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1336),
.B(n_1253),
.Y(n_1557)
);

AND2x4_ASAP7_75t_SL g1558 ( 
.A(n_1336),
.B(n_1253),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1395),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1397),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1398),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1399),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1332),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1310),
.B(n_1164),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1438),
.A2(n_858),
.B1(n_1166),
.B2(n_1164),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1400),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1427),
.B(n_1428),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_L g1568 ( 
.A(n_1392),
.B(n_1439),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1306),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1427),
.B(n_1166),
.Y(n_1570)
);

NAND2xp33_ASAP7_75t_SL g1571 ( 
.A(n_1340),
.B(n_1253),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1449),
.B(n_1266),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1449),
.B(n_1269),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1374),
.A2(n_860),
.B1(n_829),
.B2(n_1269),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1381),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1405),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1324),
.B(n_1231),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1377),
.B(n_1231),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1350),
.B(n_1231),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1279),
.A2(n_1235),
.B1(n_1198),
.B2(n_1246),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1378),
.B(n_1246),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1428),
.B(n_1441),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1284),
.B(n_1246),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1407),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1320),
.B(n_693),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1284),
.B(n_1127),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1392),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1385),
.A2(n_1129),
.B1(n_1122),
.B2(n_1112),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1337),
.B(n_1127),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1308),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1337),
.B(n_1127),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1382),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1469),
.A2(n_1121),
.B(n_1118),
.C(n_1122),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1368),
.A2(n_1121),
.B(n_1118),
.C(n_1129),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1379),
.B(n_1048),
.Y(n_1595)
);

O2A1O1Ixp5_ASAP7_75t_L g1596 ( 
.A1(n_1471),
.A2(n_1111),
.B(n_1117),
.C(n_1112),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1387),
.A2(n_1021),
.B1(n_1130),
.B2(n_1117),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1383),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1408),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1420),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1302),
.B(n_1130),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1348),
.B(n_952),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1441),
.B(n_1105),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1409),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_L g1605 ( 
.A(n_1392),
.B(n_1111),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1439),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1343),
.A2(n_1120),
.B(n_1130),
.C(n_716),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1421),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1422),
.A2(n_1021),
.B1(n_1120),
.B2(n_1105),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1412),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1343),
.A2(n_633),
.B1(n_634),
.B2(n_631),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1325),
.B(n_1105),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1325),
.B(n_1105),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1389),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1333),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1335),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1334),
.A2(n_846),
.B1(n_752),
.B2(n_788),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1448),
.B(n_1457),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1305),
.B(n_694),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1342),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1344),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1415),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1347),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1349),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1315),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1331),
.B(n_1124),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1424),
.A2(n_1021),
.B1(n_757),
.B2(n_785),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1331),
.B(n_1124),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1354),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1396),
.B(n_735),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1416),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1419),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_1294),
.Y(n_1633)
);

NOR3xp33_ASAP7_75t_L g1634 ( 
.A(n_1425),
.B(n_957),
.C(n_953),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1384),
.B(n_1124),
.Y(n_1635)
);

BUFx5_ASAP7_75t_L g1636 ( 
.A(n_1285),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1355),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_SL g1638 ( 
.A1(n_1375),
.A2(n_1404),
.B1(n_1318),
.B2(n_1380),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1375),
.B(n_1426),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1384),
.B(n_1058),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1297),
.Y(n_1641)
);

OR2x6_ASAP7_75t_L g1642 ( 
.A(n_1375),
.B(n_751),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1353),
.B(n_735),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1388),
.B(n_1058),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1439),
.B(n_1058),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1429),
.A2(n_1091),
.B1(n_1062),
.B2(n_1063),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1356),
.B(n_752),
.Y(n_1648)
);

O2A1O1Ixp33_ASAP7_75t_L g1649 ( 
.A1(n_1357),
.A2(n_731),
.B(n_738),
.C(n_703),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1430),
.A2(n_1058),
.B1(n_1063),
.B2(n_1062),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1338),
.B(n_1341),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1345),
.B(n_1062),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1431),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1282),
.B(n_785),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1285),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1388),
.B(n_1062),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1358),
.B(n_1062),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1352),
.B(n_1062),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1359),
.A2(n_634),
.B1(n_635),
.B2(n_633),
.Y(n_1659)
);

INVx5_ASAP7_75t_L g1660 ( 
.A(n_1285),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1360),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1434),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1362),
.B(n_696),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1364),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1365),
.A2(n_644),
.B1(n_647),
.B2(n_642),
.C(n_635),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1366),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1367),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1435),
.Y(n_1668)
);

AOI22x1_ASAP7_75t_L g1669 ( 
.A1(n_1471),
.A2(n_1077),
.B1(n_1085),
.B2(n_1063),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1436),
.Y(n_1670)
);

BUFx8_ASAP7_75t_L g1671 ( 
.A(n_1446),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1363),
.B(n_1063),
.Y(n_1672)
);

AO22x1_ASAP7_75t_L g1673 ( 
.A1(n_1315),
.A2(n_647),
.B1(n_648),
.B2(n_642),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_SL g1674 ( 
.A(n_1370),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1318),
.A2(n_854),
.B1(n_855),
.B2(n_789),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1371),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1394),
.B(n_698),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1473),
.B(n_1443),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1380),
.B(n_1063),
.Y(n_1679)
);

OR2x6_ASAP7_75t_L g1680 ( 
.A(n_1282),
.B(n_1423),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1329),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1289),
.B(n_1063),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1450),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1451),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1495),
.B(n_1502),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1483),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1484),
.A2(n_1330),
.B(n_1423),
.Y(n_1687)
);

A2O1A1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1489),
.A2(n_1330),
.B(n_1346),
.C(n_1289),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1474),
.A2(n_1456),
.B1(n_1460),
.B2(n_1453),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1559),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1479),
.A2(n_1456),
.B(n_1403),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1488),
.A2(n_1403),
.B(n_1462),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1549),
.B(n_1463),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1567),
.A2(n_1467),
.B(n_1465),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1492),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1567),
.A2(n_1472),
.B1(n_854),
.B2(n_855),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1560),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1582),
.A2(n_1018),
.B(n_1077),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1582),
.A2(n_1018),
.B(n_1077),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1505),
.B(n_1329),
.Y(n_1700)
);

AO21x1_ASAP7_75t_L g1701 ( 
.A1(n_1515),
.A2(n_758),
.B(n_748),
.Y(n_1701)
);

O2A1O1Ixp5_ASAP7_75t_L g1702 ( 
.A1(n_1530),
.A2(n_859),
.B(n_861),
.C(n_789),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1477),
.A2(n_1018),
.B(n_1077),
.Y(n_1703)
);

BUFx8_ASAP7_75t_L g1704 ( 
.A(n_1674),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1491),
.B(n_1329),
.Y(n_1705)
);

BUFx3_ASAP7_75t_L g1706 ( 
.A(n_1548),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1639),
.B(n_1329),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1639),
.B(n_1417),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1491),
.B(n_1417),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1482),
.B(n_1417),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1660),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1506),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1553),
.B(n_699),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1501),
.A2(n_1018),
.B(n_1077),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1590),
.B(n_1417),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1513),
.B(n_760),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1487),
.A2(n_1085),
.B(n_1077),
.Y(n_1717)
);

NOR2x1p5_ASAP7_75t_SL g1718 ( 
.A(n_1636),
.B(n_1552),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1660),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1497),
.B(n_644),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1493),
.B(n_762),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1660),
.A2(n_1091),
.B(n_1085),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1660),
.A2(n_1091),
.B(n_1085),
.Y(n_1723)
);

NOR3xp33_ASAP7_75t_L g1724 ( 
.A(n_1585),
.B(n_961),
.C(n_958),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1680),
.A2(n_1091),
.B(n_1085),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1682),
.A2(n_1596),
.B(n_1594),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1680),
.A2(n_1091),
.B(n_1085),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1680),
.A2(n_1125),
.B(n_1091),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1507),
.B(n_963),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1511),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1518),
.B(n_767),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1509),
.A2(n_1125),
.B(n_1096),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1546),
.B(n_770),
.Y(n_1733)
);

OAI321xp33_ASAP7_75t_L g1734 ( 
.A1(n_1524),
.A2(n_786),
.A3(n_781),
.B1(n_794),
.B2(n_792),
.C(n_783),
.Y(n_1734)
);

NAND2x1p5_ASAP7_75t_L g1735 ( 
.A(n_1655),
.B(n_1125),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1579),
.B(n_798),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1509),
.A2(n_1125),
.B(n_1096),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1577),
.B(n_799),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1480),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1516),
.A2(n_1125),
.B(n_1096),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1625),
.A2(n_1125),
.B(n_1096),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1496),
.B(n_804),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1510),
.B(n_648),
.Y(n_1743)
);

INVx4_ASAP7_75t_L g1744 ( 
.A(n_1606),
.Y(n_1744)
);

O2A1O1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1610),
.A2(n_823),
.B(n_828),
.C(n_806),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1512),
.B(n_649),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1490),
.A2(n_836),
.B(n_837),
.C(n_835),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1570),
.A2(n_1041),
.B(n_1039),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1555),
.B(n_1677),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1528),
.Y(n_1750)
);

O2A1O1Ixp33_ASAP7_75t_SL g1751 ( 
.A1(n_1607),
.A2(n_840),
.B(n_841),
.C(n_838),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1569),
.B(n_700),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1499),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1555),
.B(n_849),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1682),
.A2(n_966),
.B(n_965),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1561),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1531),
.B(n_1533),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1570),
.A2(n_1041),
.B(n_1039),
.Y(n_1758)
);

OAI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1626),
.A2(n_972),
.B(n_971),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1640),
.A2(n_1041),
.B(n_1039),
.Y(n_1760)
);

AOI21xp33_ASAP7_75t_L g1761 ( 
.A1(n_1647),
.A2(n_651),
.B(n_649),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1537),
.B(n_973),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1539),
.B(n_974),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1547),
.B(n_702),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1554),
.B(n_651),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1563),
.B(n_704),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1575),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1671),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1592),
.B(n_705),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1640),
.A2(n_1041),
.B(n_1039),
.Y(n_1770)
);

NOR2xp67_ASAP7_75t_SL g1771 ( 
.A(n_1608),
.B(n_654),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1644),
.A2(n_1041),
.B(n_1039),
.Y(n_1772)
);

NOR3xp33_ASAP7_75t_L g1773 ( 
.A(n_1619),
.B(n_825),
.C(n_655),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1562),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1514),
.A2(n_655),
.B1(n_658),
.B2(n_654),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1566),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1598),
.B(n_706),
.Y(n_1777)
);

NOR2xp67_ASAP7_75t_L g1778 ( 
.A(n_1600),
.B(n_602),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1614),
.A2(n_861),
.B1(n_859),
.B2(n_659),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1576),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1519),
.B(n_707),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1684),
.Y(n_1782)
);

INVx6_ASAP7_75t_L g1783 ( 
.A(n_1671),
.Y(n_1783)
);

AOI21xp33_ASAP7_75t_L g1784 ( 
.A1(n_1630),
.A2(n_1611),
.B(n_1663),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1556),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1644),
.A2(n_994),
.B(n_981),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1643),
.B(n_709),
.Y(n_1787)
);

OAI22x1_ASAP7_75t_L g1788 ( 
.A1(n_1588),
.A2(n_1618),
.B1(n_1583),
.B2(n_1591),
.Y(n_1788)
);

OR2x6_ASAP7_75t_SL g1789 ( 
.A(n_1622),
.B(n_658),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1500),
.A2(n_661),
.B1(n_662),
.B2(n_659),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1565),
.A2(n_788),
.B1(n_818),
.B2(n_752),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1617),
.B(n_661),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1648),
.B(n_788),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1681),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1656),
.A2(n_994),
.B(n_981),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1656),
.A2(n_994),
.B(n_981),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1584),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1626),
.A2(n_714),
.B(n_712),
.Y(n_1798)
);

OAI21xp33_ASAP7_75t_L g1799 ( 
.A1(n_1602),
.A2(n_665),
.B(n_662),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1500),
.B(n_715),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1545),
.A2(n_994),
.B(n_981),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1551),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1615),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1568),
.A2(n_994),
.B(n_981),
.Y(n_1804)
);

NOR2xp67_ASAP7_75t_L g1805 ( 
.A(n_1641),
.B(n_603),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1628),
.A2(n_1036),
.B(n_1028),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1661),
.B(n_717),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1664),
.B(n_718),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1666),
.B(n_1520),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1633),
.A2(n_719),
.B1(n_722),
.B2(n_721),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1616),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1638),
.B(n_665),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1599),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1565),
.B(n_723),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1481),
.B(n_726),
.Y(n_1815)
);

AO21x1_ASAP7_75t_L g1816 ( 
.A1(n_1586),
.A2(n_2),
.B(n_1),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1481),
.B(n_727),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1649),
.A2(n_825),
.B(n_827),
.C(n_749),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1572),
.B(n_728),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1557),
.B(n_1665),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1551),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1673),
.B(n_818),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1551),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1573),
.B(n_729),
.Y(n_1824)
);

AOI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1628),
.A2(n_1036),
.B(n_1028),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1517),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1678),
.B(n_732),
.Y(n_1827)
);

O2A1O1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1589),
.A2(n_846),
.B(n_818),
.C(n_740),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1620),
.B(n_739),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1674),
.Y(n_1830)
);

AOI21x1_ASAP7_75t_L g1831 ( 
.A1(n_1635),
.A2(n_1033),
.B(n_1027),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1621),
.B(n_742),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1635),
.A2(n_1036),
.B(n_1028),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1508),
.A2(n_1036),
.B(n_1028),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1604),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1571),
.A2(n_744),
.B1(n_746),
.B2(n_743),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1603),
.A2(n_1036),
.B(n_1028),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1603),
.A2(n_754),
.B(n_753),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1612),
.A2(n_978),
.B(n_1013),
.Y(n_1839)
);

NOR3xp33_ASAP7_75t_L g1840 ( 
.A(n_1659),
.B(n_867),
.C(n_845),
.Y(n_1840)
);

NAND2x1p5_ASAP7_75t_L g1841 ( 
.A(n_1655),
.B(n_978),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1634),
.A2(n_846),
.B1(n_756),
.B2(n_765),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1612),
.A2(n_1013),
.B(n_1033),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1631),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1623),
.B(n_763),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1624),
.B(n_766),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1613),
.A2(n_1013),
.B(n_1033),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1613),
.A2(n_1669),
.B(n_1605),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1476),
.B(n_749),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1606),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1558),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1629),
.Y(n_1852)
);

OAI21xp33_ASAP7_75t_L g1853 ( 
.A1(n_1597),
.A2(n_1642),
.B(n_831),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1475),
.A2(n_1498),
.B(n_1494),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1679),
.A2(n_1013),
.B(n_1033),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1580),
.A2(n_1013),
.B(n_1033),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1593),
.A2(n_605),
.B(n_604),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1637),
.B(n_769),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1606),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1632),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1544),
.B(n_607),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1654),
.A2(n_609),
.B(n_608),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1667),
.B(n_771),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1642),
.B(n_1485),
.Y(n_1864)
);

BUFx3_ASAP7_75t_L g1865 ( 
.A(n_1642),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1676),
.B(n_773),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1486),
.B(n_774),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1478),
.Y(n_1868)
);

AND2x2_ASAP7_75t_SL g1869 ( 
.A(n_1653),
.B(n_1662),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1544),
.A2(n_831),
.B1(n_832),
.B2(n_827),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1654),
.A2(n_611),
.B(n_610),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1654),
.A2(n_1527),
.B(n_1504),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1683),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1504),
.A2(n_613),
.B(n_612),
.Y(n_1874)
);

AOI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1527),
.A2(n_1532),
.B(n_1529),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1529),
.A2(n_615),
.B(n_614),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1532),
.A2(n_618),
.B(n_616),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1668),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1670),
.A2(n_839),
.B(n_842),
.C(n_832),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1538),
.A2(n_777),
.B(n_776),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1535),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1544),
.A2(n_842),
.B1(n_843),
.B2(n_839),
.Y(n_1882)
);

NAND2x1p5_ASAP7_75t_L g1883 ( 
.A(n_1478),
.B(n_619),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1757),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1685),
.A2(n_1601),
.B1(n_1650),
.B2(n_1646),
.Y(n_1885)
);

BUFx6f_ASAP7_75t_L g1886 ( 
.A(n_1850),
.Y(n_1886)
);

AOI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1687),
.A2(n_1543),
.B(n_1538),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1729),
.B(n_1693),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1739),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1690),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1784),
.B(n_1749),
.Y(n_1891)
);

NOR2x1p5_ASAP7_75t_L g1892 ( 
.A(n_1706),
.B(n_1503),
.Y(n_1892)
);

INVx5_ASAP7_75t_L g1893 ( 
.A(n_1711),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1787),
.B(n_1540),
.Y(n_1894)
);

NAND2x1p5_ASAP7_75t_L g1895 ( 
.A(n_1711),
.B(n_1542),
.Y(n_1895)
);

AO21x1_ASAP7_75t_L g1896 ( 
.A1(n_1696),
.A2(n_1675),
.B(n_1574),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1815),
.B(n_1574),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1869),
.A2(n_1550),
.B1(n_1564),
.B2(n_1543),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1719),
.Y(n_1899)
);

O2A1O1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1761),
.A2(n_1675),
.B(n_1651),
.C(n_1595),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_SL g1901 ( 
.A1(n_1816),
.A2(n_1564),
.B(n_1550),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1812),
.B(n_1534),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1720),
.B(n_1534),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1697),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1773),
.B(n_1636),
.Y(n_1905)
);

OAI21xp33_ASAP7_75t_L g1906 ( 
.A1(n_1791),
.A2(n_845),
.B(n_843),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1817),
.B(n_1521),
.Y(n_1907)
);

NOR2xp67_ASAP7_75t_L g1908 ( 
.A(n_1719),
.B(n_1542),
.Y(n_1908)
);

NAND2x1p5_ASAP7_75t_L g1909 ( 
.A(n_1744),
.B(n_1587),
.Y(n_1909)
);

AOI33xp33_ASAP7_75t_L g1910 ( 
.A1(n_1842),
.A2(n_864),
.A3(n_852),
.B1(n_865),
.B2(n_863),
.B3(n_851),
.Y(n_1910)
);

BUFx12f_ASAP7_75t_L g1911 ( 
.A(n_1704),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1707),
.B(n_1587),
.Y(n_1912)
);

INVx1_ASAP7_75t_SL g1913 ( 
.A(n_1785),
.Y(n_1913)
);

O2A1O1Ixp33_ASAP7_75t_L g1914 ( 
.A1(n_1792),
.A2(n_1523),
.B(n_1525),
.C(n_1522),
.Y(n_1914)
);

OR2x6_ASAP7_75t_SL g1915 ( 
.A(n_1870),
.B(n_851),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1814),
.A2(n_1541),
.B1(n_1526),
.B2(n_1581),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1826),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_L g1918 ( 
.A(n_1778),
.B(n_1578),
.Y(n_1918)
);

CKINVDCx20_ASAP7_75t_R g1919 ( 
.A(n_1704),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1753),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1734),
.B(n_1636),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1840),
.A2(n_1536),
.B1(n_863),
.B2(n_864),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1820),
.A2(n_780),
.B1(n_787),
.B2(n_779),
.Y(n_1923)
);

BUFx4f_ASAP7_75t_L g1924 ( 
.A(n_1783),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1827),
.B(n_793),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1688),
.A2(n_1848),
.B(n_1691),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1875),
.A2(n_1645),
.B(n_1657),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1721),
.B(n_852),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1734),
.B(n_1636),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1800),
.B(n_865),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1700),
.A2(n_1609),
.B1(n_1657),
.B2(n_1627),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1713),
.A2(n_1851),
.B1(n_1710),
.B2(n_1709),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1809),
.B(n_1788),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1716),
.B(n_866),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1805),
.B(n_1636),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1872),
.A2(n_1658),
.B(n_1652),
.Y(n_1936)
);

A2O1A1Ixp33_ASAP7_75t_L g1937 ( 
.A1(n_1828),
.A2(n_1672),
.B(n_867),
.C(n_868),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1692),
.A2(n_1694),
.B(n_1726),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1726),
.A2(n_1636),
.B(n_1536),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_R g1940 ( 
.A(n_1794),
.B(n_1536),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1810),
.B(n_800),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1707),
.Y(n_1942)
);

O2A1O1Ixp5_ASAP7_75t_SL g1943 ( 
.A1(n_1696),
.A2(n_868),
.B(n_869),
.C(n_866),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1819),
.B(n_803),
.Y(n_1944)
);

AOI21x1_ASAP7_75t_L g1945 ( 
.A1(n_1831),
.A2(n_1536),
.B(n_621),
.Y(n_1945)
);

AOI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1732),
.A2(n_1536),
.B(n_624),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1756),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1737),
.A2(n_620),
.B(n_805),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1742),
.B(n_1824),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1793),
.B(n_807),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1880),
.B(n_869),
.Y(n_1951)
);

NAND2x1p5_ASAP7_75t_L g1952 ( 
.A(n_1744),
.B(n_0),
.Y(n_1952)
);

OAI21xp33_ASAP7_75t_L g1953 ( 
.A1(n_1736),
.A2(n_871),
.B(n_870),
.Y(n_1953)
);

INVx5_ASAP7_75t_L g1954 ( 
.A(n_1850),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1880),
.B(n_870),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1774),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1725),
.A2(n_1728),
.B(n_1727),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1781),
.B(n_871),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1738),
.B(n_872),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1864),
.B(n_809),
.Y(n_1960)
);

OAI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1851),
.A2(n_872),
.B1(n_811),
.B2(n_812),
.Y(n_1961)
);

NAND2xp33_ASAP7_75t_L g1962 ( 
.A(n_1853),
.B(n_810),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1754),
.B(n_813),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1799),
.B(n_814),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1686),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1717),
.A2(n_1689),
.B(n_1714),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1733),
.B(n_817),
.Y(n_1967)
);

OAI22x1_ASAP7_75t_L g1968 ( 
.A1(n_1822),
.A2(n_821),
.B1(n_822),
.B2(n_819),
.Y(n_1968)
);

NOR2x1_ASAP7_75t_L g1969 ( 
.A(n_1802),
.B(n_824),
.Y(n_1969)
);

BUFx12f_ASAP7_75t_L g1970 ( 
.A(n_1783),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1731),
.B(n_1798),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1722),
.A2(n_873),
.B(n_2),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1798),
.B(n_3),
.Y(n_1973)
);

NAND2x1p5_ASAP7_75t_L g1974 ( 
.A(n_1708),
.B(n_3),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_SL g1975 ( 
.A(n_1830),
.B(n_4),
.Y(n_1975)
);

A2O1A1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1838),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1838),
.B(n_7),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1695),
.Y(n_1978)
);

AOI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1723),
.A2(n_8),
.B(n_9),
.Y(n_1979)
);

AO32x2_ASAP7_75t_L g1980 ( 
.A1(n_1779),
.A2(n_1870),
.A3(n_1790),
.B1(n_1775),
.B2(n_1882),
.Y(n_1980)
);

AOI21xp33_ASAP7_75t_L g1981 ( 
.A1(n_1705),
.A2(n_8),
.B(n_10),
.Y(n_1981)
);

NAND2x1p5_ASAP7_75t_L g1982 ( 
.A(n_1708),
.B(n_10),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1746),
.B(n_11),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1765),
.B(n_11),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1703),
.A2(n_1699),
.B(n_1698),
.Y(n_1985)
);

BUFx8_ASAP7_75t_SL g1986 ( 
.A(n_1768),
.Y(n_1986)
);

INVx4_ASAP7_75t_L g1987 ( 
.A(n_1850),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1854),
.A2(n_12),
.B(n_13),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1752),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1807),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1990)
);

INVx4_ASAP7_75t_L g1991 ( 
.A(n_1859),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1790),
.B(n_16),
.Y(n_1992)
);

AOI22xp5_ASAP7_75t_L g1993 ( 
.A1(n_1724),
.A2(n_1743),
.B1(n_1779),
.B2(n_1818),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1868),
.Y(n_1994)
);

A2O1A1Ixp33_ASAP7_75t_L g1995 ( 
.A1(n_1857),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_1995)
);

O2A1O1Ixp33_ASAP7_75t_L g1996 ( 
.A1(n_1747),
.A2(n_591),
.B(n_592),
.C(n_590),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1762),
.B(n_17),
.Y(n_1997)
);

O2A1O1Ixp33_ASAP7_75t_L g1998 ( 
.A1(n_1879),
.A2(n_593),
.B(n_594),
.C(n_592),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1741),
.A2(n_18),
.B(n_19),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1763),
.B(n_20),
.Y(n_2000)
);

OR2x6_ASAP7_75t_L g2001 ( 
.A(n_1861),
.B(n_21),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1856),
.A2(n_1876),
.B(n_1874),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1865),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1849),
.B(n_26),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1776),
.B(n_26),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1877),
.A2(n_27),
.B(n_29),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1780),
.B(n_29),
.Y(n_2007)
);

OAI22x1_ASAP7_75t_L g2008 ( 
.A1(n_1861),
.A2(n_1803),
.B1(n_1811),
.B2(n_1782),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1808),
.B(n_30),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1797),
.B(n_30),
.Y(n_2010)
);

AOI221xp5_ASAP7_75t_L g2011 ( 
.A1(n_1745),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.C(n_34),
.Y(n_2011)
);

O2A1O1Ixp5_ASAP7_75t_L g2012 ( 
.A1(n_1701),
.A2(n_1702),
.B(n_1755),
.C(n_1759),
.Y(n_2012)
);

OAI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1852),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1813),
.B(n_34),
.Y(n_2014)
);

BUFx4f_ASAP7_75t_L g2015 ( 
.A(n_1859),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1712),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1755),
.A2(n_1834),
.B(n_1740),
.Y(n_2017)
);

AOI22x1_ASAP7_75t_SL g2018 ( 
.A1(n_1802),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_SL g2019 ( 
.A(n_1859),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1759),
.A2(n_38),
.B(n_39),
.Y(n_2020)
);

A2O1A1Ixp33_ASAP7_75t_L g2021 ( 
.A1(n_1862),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1730),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1871),
.A2(n_1847),
.B(n_1843),
.Y(n_2023)
);

AO22x1_ASAP7_75t_L g2024 ( 
.A1(n_1715),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_2024)
);

A2O1A1Ixp33_ASAP7_75t_L g2025 ( 
.A1(n_1836),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2025)
);

AOI21xp5_ASAP7_75t_L g2026 ( 
.A1(n_1839),
.A2(n_44),
.B(n_45),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1750),
.Y(n_2027)
);

AND2x2_ASAP7_75t_SL g2028 ( 
.A(n_1821),
.B(n_1823),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1835),
.B(n_45),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1829),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2030)
);

AOI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1748),
.A2(n_47),
.B(n_48),
.Y(n_2031)
);

NOR2x1_ASAP7_75t_L g2032 ( 
.A(n_1821),
.B(n_585),
.Y(n_2032)
);

INVx4_ASAP7_75t_L g2033 ( 
.A(n_1794),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1823),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1715),
.B(n_49),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1844),
.B(n_1860),
.Y(n_2036)
);

NOR2xp67_ASAP7_75t_SL g2037 ( 
.A(n_1832),
.B(n_50),
.Y(n_2037)
);

AOI22xp33_ASAP7_75t_L g2038 ( 
.A1(n_1845),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1758),
.A2(n_1825),
.B(n_1806),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1878),
.B(n_51),
.Y(n_2040)
);

AOI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_1846),
.A2(n_1863),
.B1(n_1866),
.B2(n_1858),
.Y(n_2041)
);

INVx3_ASAP7_75t_L g2042 ( 
.A(n_1883),
.Y(n_2042)
);

NOR2x1_ASAP7_75t_L g2043 ( 
.A(n_1873),
.B(n_589),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1767),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1883),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1881),
.B(n_54),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_SL g2047 ( 
.A1(n_1764),
.A2(n_64),
.B1(n_72),
.B2(n_56),
.Y(n_2047)
);

INVxp67_ASAP7_75t_L g2048 ( 
.A(n_1867),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1766),
.B(n_57),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1868),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1833),
.A2(n_57),
.B(n_58),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1769),
.B(n_58),
.Y(n_2052)
);

AOI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_1751),
.A2(n_59),
.B(n_60),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1777),
.B(n_1789),
.Y(n_2054)
);

OR2x6_ASAP7_75t_SL g2055 ( 
.A(n_1771),
.B(n_599),
.Y(n_2055)
);

AND2x2_ASAP7_75t_SL g2056 ( 
.A(n_1718),
.B(n_598),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1735),
.B(n_1841),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1735),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1841),
.Y(n_2059)
);

INVx1_ASAP7_75t_SL g2060 ( 
.A(n_1855),
.Y(n_2060)
);

INVx3_ASAP7_75t_L g2061 ( 
.A(n_2033),
.Y(n_2061)
);

BUFx2_ASAP7_75t_L g2062 ( 
.A(n_1917),
.Y(n_2062)
);

AOI21xp5_ASAP7_75t_L g2063 ( 
.A1(n_2002),
.A2(n_1772),
.B(n_1770),
.Y(n_2063)
);

NAND3x1_ASAP7_75t_L g2064 ( 
.A(n_1891),
.B(n_61),
.C(n_62),
.Y(n_2064)
);

AOI21x1_ASAP7_75t_L g2065 ( 
.A1(n_1945),
.A2(n_1760),
.B(n_1786),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1938),
.A2(n_1837),
.B(n_1796),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1965),
.Y(n_2067)
);

AOI21xp33_ASAP7_75t_L g2068 ( 
.A1(n_1971),
.A2(n_1795),
.B(n_1801),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_1957),
.A2(n_1804),
.B(n_62),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_SL g2070 ( 
.A1(n_2020),
.A2(n_63),
.B(n_65),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_SL g2071 ( 
.A1(n_2001),
.A2(n_595),
.B(n_584),
.Y(n_2071)
);

AOI21x1_ASAP7_75t_L g2072 ( 
.A1(n_1939),
.A2(n_65),
.B(n_66),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_2033),
.Y(n_2073)
);

CKINVDCx11_ASAP7_75t_R g2074 ( 
.A(n_1911),
.Y(n_2074)
);

INVx3_ASAP7_75t_L g2075 ( 
.A(n_1942),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_2034),
.B(n_66),
.Y(n_2076)
);

BUFx10_ASAP7_75t_L g2077 ( 
.A(n_1894),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_2039),
.A2(n_67),
.B(n_68),
.Y(n_2078)
);

AO31x2_ASAP7_75t_L g2079 ( 
.A1(n_1966),
.A2(n_2017),
.A3(n_1985),
.B(n_1926),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1888),
.B(n_67),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1949),
.B(n_68),
.Y(n_2081)
);

NAND2x1p5_ASAP7_75t_L g2082 ( 
.A(n_1954),
.B(n_69),
.Y(n_2082)
);

NAND2x1p5_ASAP7_75t_L g2083 ( 
.A(n_1954),
.B(n_69),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1942),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1884),
.B(n_70),
.Y(n_2085)
);

OAI21x1_ASAP7_75t_L g2086 ( 
.A1(n_2023),
.A2(n_1887),
.B(n_1927),
.Y(n_2086)
);

AOI21x1_ASAP7_75t_L g2087 ( 
.A1(n_1921),
.A2(n_70),
.B(n_71),
.Y(n_2087)
);

A2O1A1Ixp33_ASAP7_75t_L g2088 ( 
.A1(n_1993),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_2088)
);

OAI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_1925),
.A2(n_74),
.B(n_75),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1993),
.A2(n_77),
.B(n_74),
.C(n_76),
.Y(n_2090)
);

OAI21x1_ASAP7_75t_L g2091 ( 
.A1(n_1936),
.A2(n_76),
.B(n_77),
.Y(n_2091)
);

NOR2xp67_ASAP7_75t_SL g2092 ( 
.A(n_1970),
.B(n_78),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1907),
.B(n_78),
.Y(n_2093)
);

OAI21x1_ASAP7_75t_L g2094 ( 
.A1(n_1946),
.A2(n_79),
.B(n_80),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1897),
.B(n_1932),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1978),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_1948),
.A2(n_1929),
.B(n_1935),
.Y(n_2097)
);

OAI21xp33_ASAP7_75t_L g2098 ( 
.A1(n_1923),
.A2(n_79),
.B(n_81),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1889),
.B(n_81),
.Y(n_2099)
);

OAI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_2012),
.A2(n_586),
.B(n_585),
.Y(n_2100)
);

OAI21x1_ASAP7_75t_L g2101 ( 
.A1(n_1901),
.A2(n_82),
.B(n_83),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2022),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2041),
.B(n_82),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2048),
.B(n_83),
.Y(n_2104)
);

INVx2_ASAP7_75t_SL g2105 ( 
.A(n_1924),
.Y(n_2105)
);

INVx2_ASAP7_75t_SL g2106 ( 
.A(n_1924),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1973),
.B(n_84),
.Y(n_2107)
);

INVx3_ASAP7_75t_L g2108 ( 
.A(n_2034),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_2031),
.A2(n_1999),
.B(n_2006),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_1898),
.A2(n_593),
.B(n_591),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2027),
.Y(n_2111)
);

OAI21x1_ASAP7_75t_L g2112 ( 
.A1(n_2051),
.A2(n_84),
.B(n_85),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2050),
.B(n_85),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1977),
.B(n_86),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_1916),
.A2(n_597),
.B(n_596),
.Y(n_2115)
);

AOI21xp33_ASAP7_75t_L g2116 ( 
.A1(n_1951),
.A2(n_86),
.B(n_87),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1994),
.B(n_1890),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2029),
.B(n_87),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1904),
.B(n_88),
.Y(n_2119)
);

AO31x2_ASAP7_75t_L g2120 ( 
.A1(n_1896),
.A2(n_91),
.A3(n_89),
.B(n_90),
.Y(n_2120)
);

OAI21xp33_ASAP7_75t_L g2121 ( 
.A1(n_1923),
.A2(n_89),
.B(n_90),
.Y(n_2121)
);

OAI21x1_ASAP7_75t_L g2122 ( 
.A1(n_2026),
.A2(n_92),
.B(n_93),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_1886),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1947),
.B(n_1956),
.Y(n_2124)
);

AO21x1_ASAP7_75t_L g2125 ( 
.A1(n_1955),
.A2(n_93),
.B(n_94),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2036),
.B(n_94),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2008),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1913),
.B(n_601),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1912),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_2015),
.Y(n_2130)
);

OAI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_1943),
.A2(n_95),
.B(n_96),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1992),
.B(n_597),
.Y(n_2132)
);

INVx4_ASAP7_75t_L g2133 ( 
.A(n_1954),
.Y(n_2133)
);

AOI221x1_ASAP7_75t_L g2134 ( 
.A1(n_1976),
.A2(n_2025),
.B1(n_2021),
.B2(n_1988),
.C(n_1995),
.Y(n_2134)
);

OAI21x1_ASAP7_75t_L g2135 ( 
.A1(n_1933),
.A2(n_95),
.B(n_97),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1902),
.B(n_596),
.Y(n_2136)
);

OAI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_1972),
.A2(n_97),
.B(n_99),
.Y(n_2137)
);

OAI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1915),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_2138)
);

AOI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_1885),
.A2(n_101),
.B(n_102),
.Y(n_2139)
);

AOI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_1905),
.A2(n_1914),
.B(n_2060),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_2028),
.B(n_102),
.Y(n_2141)
);

AOI211x1_ASAP7_75t_L g2142 ( 
.A1(n_1989),
.A2(n_1990),
.B(n_2024),
.C(n_2016),
.Y(n_2142)
);

OAI21x1_ASAP7_75t_SL g2143 ( 
.A1(n_1998),
.A2(n_103),
.B(n_104),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1997),
.B(n_103),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_2019),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_1918),
.A2(n_105),
.B(n_106),
.Y(n_2146)
);

A2O1A1Ixp33_ASAP7_75t_L g2147 ( 
.A1(n_2009),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2007),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2000),
.B(n_1903),
.Y(n_2149)
);

OAI21x1_ASAP7_75t_L g2150 ( 
.A1(n_2042),
.A2(n_2045),
.B(n_1979),
.Y(n_2150)
);

OAI21x1_ASAP7_75t_L g2151 ( 
.A1(n_2042),
.A2(n_108),
.B(n_109),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2052),
.B(n_595),
.Y(n_2152)
);

OAI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_1900),
.A2(n_109),
.B(n_110),
.Y(n_2153)
);

OAI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_2053),
.A2(n_110),
.B(n_111),
.Y(n_2154)
);

OAI22xp5_ASAP7_75t_L g2155 ( 
.A1(n_2001),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2005),
.B(n_112),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_1941),
.A2(n_117),
.B1(n_114),
.B2(n_115),
.Y(n_2157)
);

OAI21x1_ASAP7_75t_L g2158 ( 
.A1(n_2045),
.A2(n_2057),
.B(n_1931),
.Y(n_2158)
);

AO31x2_ASAP7_75t_L g2159 ( 
.A1(n_2059),
.A2(n_118),
.A3(n_114),
.B(n_117),
.Y(n_2159)
);

BUFx5_ASAP7_75t_L g2160 ( 
.A(n_2056),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2010),
.B(n_118),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2014),
.Y(n_2162)
);

OAI21x1_ASAP7_75t_L g2163 ( 
.A1(n_1899),
.A2(n_1969),
.B(n_1895),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_2054),
.B(n_1944),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1962),
.A2(n_1893),
.B(n_2001),
.Y(n_2165)
);

BUFx3_ASAP7_75t_L g2166 ( 
.A(n_1920),
.Y(n_2166)
);

AND2x2_ASAP7_75t_SL g2167 ( 
.A(n_2011),
.B(n_594),
.Y(n_2167)
);

O2A1O1Ixp5_ASAP7_75t_L g2168 ( 
.A1(n_2037),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2035),
.B(n_119),
.Y(n_2169)
);

INVx4_ASAP7_75t_L g2170 ( 
.A(n_2015),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2040),
.B(n_1928),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2046),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_1893),
.A2(n_121),
.B(n_122),
.Y(n_2173)
);

OAI21x1_ASAP7_75t_L g2174 ( 
.A1(n_1899),
.A2(n_122),
.B(n_123),
.Y(n_2174)
);

NAND3x1_ASAP7_75t_L g2175 ( 
.A(n_2032),
.B(n_2043),
.C(n_1984),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_1893),
.A2(n_123),
.B(n_125),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2035),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2049),
.B(n_126),
.Y(n_2178)
);

HB1xp67_ASAP7_75t_L g2179 ( 
.A(n_1892),
.Y(n_2179)
);

OAI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_1937),
.A2(n_126),
.B(n_127),
.Y(n_2180)
);

INVx1_ASAP7_75t_SL g2181 ( 
.A(n_1960),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1912),
.B(n_128),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1886),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_2130),
.Y(n_2184)
);

OAI221xp5_ASAP7_75t_L g2185 ( 
.A1(n_2089),
.A2(n_1906),
.B1(n_1964),
.B2(n_2047),
.C(n_1953),
.Y(n_2185)
);

HB1xp67_ASAP7_75t_L g2186 ( 
.A(n_2127),
.Y(n_2186)
);

AOI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_2098),
.A2(n_1983),
.B1(n_2018),
.B2(n_1975),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2067),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2096),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_2117),
.Y(n_2190)
);

AOI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_2100),
.A2(n_1996),
.B(n_1981),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_2108),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2100),
.A2(n_1930),
.B(n_1963),
.Y(n_2193)
);

AOI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_2063),
.A2(n_1958),
.B(n_1967),
.Y(n_2194)
);

INVx1_ASAP7_75t_SL g2195 ( 
.A(n_2077),
.Y(n_2195)
);

OR2x6_ASAP7_75t_L g2196 ( 
.A(n_2165),
.B(n_1974),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_2167),
.A2(n_2030),
.B1(n_2038),
.B2(n_1922),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2095),
.B(n_2148),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_2164),
.B(n_2055),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2181),
.B(n_2004),
.Y(n_2200)
);

AOI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_2066),
.A2(n_1959),
.B(n_1908),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_SL g2202 ( 
.A(n_2077),
.B(n_1968),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2162),
.B(n_1934),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2149),
.B(n_1910),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2102),
.B(n_1953),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2111),
.B(n_1987),
.Y(n_2206)
);

OAI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2157),
.A2(n_2064),
.B1(n_2090),
.B2(n_2088),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2175),
.A2(n_2003),
.B1(n_1982),
.B2(n_1952),
.Y(n_2208)
);

A2O1A1Ixp33_ASAP7_75t_L g2209 ( 
.A1(n_2098),
.A2(n_1906),
.B(n_2058),
.C(n_2044),
.Y(n_2209)
);

INVx1_ASAP7_75t_SL g2210 ( 
.A(n_2166),
.Y(n_2210)
);

O2A1O1Ixp33_ASAP7_75t_SL g2211 ( 
.A1(n_2147),
.A2(n_2013),
.B(n_1919),
.C(n_1961),
.Y(n_2211)
);

INVx3_ASAP7_75t_L g2212 ( 
.A(n_2108),
.Y(n_2212)
);

OAI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_2121),
.A2(n_1950),
.B1(n_1908),
.B2(n_1909),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_2074),
.Y(n_2214)
);

AOI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_2153),
.A2(n_1940),
.B(n_1980),
.Y(n_2215)
);

AOI21xp33_ASAP7_75t_SL g2216 ( 
.A1(n_2138),
.A2(n_1986),
.B(n_128),
.Y(n_2216)
);

BUFx3_ASAP7_75t_L g2217 ( 
.A(n_2062),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_2160),
.B(n_1886),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2159),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2121),
.A2(n_1980),
.B1(n_1991),
.B2(n_1987),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_2181),
.B(n_2179),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2160),
.B(n_1991),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_2061),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2124),
.Y(n_2224)
);

OAI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_2103),
.A2(n_1980),
.B1(n_131),
.B2(n_129),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_2061),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_2075),
.B(n_129),
.Y(n_2227)
);

NOR2x1_ASAP7_75t_SL g2228 ( 
.A(n_2133),
.B(n_130),
.Y(n_2228)
);

INVx2_ASAP7_75t_SL g2229 ( 
.A(n_2123),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2159),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2159),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2172),
.B(n_130),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2120),
.Y(n_2233)
);

CKINVDCx5p33_ASAP7_75t_R g2234 ( 
.A(n_2105),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_2145),
.Y(n_2235)
);

INVx3_ASAP7_75t_SL g2236 ( 
.A(n_2106),
.Y(n_2236)
);

O2A1O1Ixp33_ASAP7_75t_L g2237 ( 
.A1(n_2153),
.A2(n_2154),
.B(n_2137),
.C(n_2139),
.Y(n_2237)
);

AOI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_2140),
.A2(n_131),
.B(n_132),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2177),
.B(n_132),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_2160),
.A2(n_2137),
.B1(n_2180),
.B2(n_2116),
.Y(n_2240)
);

OAI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_2142),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_2086),
.A2(n_135),
.B(n_136),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2182),
.B(n_136),
.Y(n_2243)
);

NOR2xp67_ASAP7_75t_L g2244 ( 
.A(n_2097),
.B(n_137),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2075),
.B(n_137),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_R g2246 ( 
.A(n_2130),
.B(n_138),
.Y(n_2246)
);

BUFx3_ASAP7_75t_L g2247 ( 
.A(n_2123),
.Y(n_2247)
);

AOI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2154),
.A2(n_2109),
.B(n_2134),
.Y(n_2248)
);

AND2x4_ASAP7_75t_L g2249 ( 
.A(n_2084),
.B(n_138),
.Y(n_2249)
);

NOR2xp67_ASAP7_75t_L g2250 ( 
.A(n_2073),
.B(n_139),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_2068),
.A2(n_139),
.B(n_140),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_2073),
.Y(n_2252)
);

INVx3_ASAP7_75t_L g2253 ( 
.A(n_2133),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_2130),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2129),
.B(n_589),
.Y(n_2255)
);

AND2x4_ASAP7_75t_L g2256 ( 
.A(n_2084),
.B(n_141),
.Y(n_2256)
);

INVx5_ASAP7_75t_L g2257 ( 
.A(n_2076),
.Y(n_2257)
);

OAI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_2142),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_2163),
.Y(n_2259)
);

INVxp67_ASAP7_75t_L g2260 ( 
.A(n_2183),
.Y(n_2260)
);

AOI22xp33_ASAP7_75t_SL g2261 ( 
.A1(n_2207),
.A2(n_2160),
.B1(n_2180),
.B2(n_2143),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2190),
.B(n_2186),
.Y(n_2262)
);

INVx2_ASAP7_75t_SL g2263 ( 
.A(n_2217),
.Y(n_2263)
);

INVx1_ASAP7_75t_SL g2264 ( 
.A(n_2195),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2200),
.B(n_2160),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2188),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2189),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2187),
.A2(n_2185),
.B1(n_2240),
.B2(n_2209),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2219),
.Y(n_2269)
);

AOI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_2197),
.A2(n_2155),
.B1(n_2115),
.B2(n_2114),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2224),
.Y(n_2271)
);

AOI22xp33_ASAP7_75t_L g2272 ( 
.A1(n_2193),
.A2(n_2107),
.B1(n_2070),
.B2(n_2125),
.Y(n_2272)
);

AOI22xp5_ASAP7_75t_SL g2273 ( 
.A1(n_2199),
.A2(n_2145),
.B1(n_2110),
.B2(n_2136),
.Y(n_2273)
);

INVx6_ASAP7_75t_L g2274 ( 
.A(n_2257),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_2187),
.A2(n_2132),
.B1(n_2141),
.B2(n_2152),
.Y(n_2275)
);

BUFx12f_ASAP7_75t_L g2276 ( 
.A(n_2214),
.Y(n_2276)
);

BUFx12f_ASAP7_75t_L g2277 ( 
.A(n_2234),
.Y(n_2277)
);

BUFx5_ASAP7_75t_L g2278 ( 
.A(n_2230),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2259),
.Y(n_2279)
);

BUFx2_ASAP7_75t_SL g2280 ( 
.A(n_2257),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_2210),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_2260),
.Y(n_2282)
);

BUFx2_ASAP7_75t_L g2283 ( 
.A(n_2192),
.Y(n_2283)
);

INVx5_ASAP7_75t_L g2284 ( 
.A(n_2196),
.Y(n_2284)
);

CKINVDCx11_ASAP7_75t_R g2285 ( 
.A(n_2236),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2231),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2233),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2259),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2198),
.Y(n_2289)
);

AOI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2208),
.A2(n_2092),
.B1(n_2171),
.B2(n_2146),
.Y(n_2290)
);

AOI22xp33_ASAP7_75t_L g2291 ( 
.A1(n_2191),
.A2(n_2131),
.B1(n_2178),
.B2(n_2144),
.Y(n_2291)
);

AOI22xp33_ASAP7_75t_L g2292 ( 
.A1(n_2241),
.A2(n_2131),
.B1(n_2161),
.B2(n_2156),
.Y(n_2292)
);

BUFx10_ASAP7_75t_L g2293 ( 
.A(n_2227),
.Y(n_2293)
);

INVx6_ASAP7_75t_L g2294 ( 
.A(n_2257),
.Y(n_2294)
);

CKINVDCx11_ASAP7_75t_R g2295 ( 
.A(n_2235),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_2246),
.Y(n_2296)
);

OAI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2237),
.A2(n_2071),
.B1(n_2083),
.B2(n_2082),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2221),
.B(n_2080),
.Y(n_2298)
);

CKINVDCx20_ASAP7_75t_R g2299 ( 
.A(n_2247),
.Y(n_2299)
);

AOI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_2258),
.A2(n_2081),
.B1(n_2093),
.B2(n_2104),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2203),
.B(n_2099),
.Y(n_2301)
);

AOI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_2225),
.A2(n_2176),
.B1(n_2173),
.B2(n_2112),
.Y(n_2302)
);

CKINVDCx6p67_ASAP7_75t_R g2303 ( 
.A(n_2184),
.Y(n_2303)
);

AOI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_2215),
.A2(n_2122),
.B1(n_2118),
.B2(n_2113),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2212),
.Y(n_2305)
);

CKINVDCx20_ASAP7_75t_R g2306 ( 
.A(n_2184),
.Y(n_2306)
);

CKINVDCx11_ASAP7_75t_R g2307 ( 
.A(n_2184),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2212),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2206),
.B(n_2113),
.Y(n_2309)
);

BUFx12f_ASAP7_75t_L g2310 ( 
.A(n_2227),
.Y(n_2310)
);

BUFx2_ASAP7_75t_SL g2311 ( 
.A(n_2229),
.Y(n_2311)
);

O2A1O1Ixp33_ASAP7_75t_L g2312 ( 
.A1(n_2268),
.A2(n_2216),
.B(n_2211),
.C(n_2238),
.Y(n_2312)
);

OR2x2_ASAP7_75t_L g2313 ( 
.A(n_2262),
.B(n_2079),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2289),
.B(n_2282),
.Y(n_2314)
);

AOI21x1_ASAP7_75t_SL g2315 ( 
.A1(n_2301),
.A2(n_2204),
.B(n_2232),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2283),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2265),
.B(n_2223),
.Y(n_2317)
);

O2A1O1Ixp5_ASAP7_75t_L g2318 ( 
.A1(n_2297),
.A2(n_2248),
.B(n_2202),
.C(n_2222),
.Y(n_2318)
);

O2A1O1Ixp33_ASAP7_75t_L g2319 ( 
.A1(n_2270),
.A2(n_2213),
.B(n_2194),
.C(n_2168),
.Y(n_2319)
);

OAI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2270),
.A2(n_2220),
.B1(n_2244),
.B2(n_2251),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2279),
.B(n_2223),
.Y(n_2321)
);

OAI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2275),
.A2(n_2261),
.B1(n_2300),
.B2(n_2292),
.Y(n_2322)
);

BUFx8_ASAP7_75t_SL g2323 ( 
.A(n_2276),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2287),
.Y(n_2324)
);

O2A1O1Ixp33_ASAP7_75t_L g2325 ( 
.A1(n_2291),
.A2(n_2205),
.B(n_2242),
.C(n_2218),
.Y(n_2325)
);

AOI21x1_ASAP7_75t_SL g2326 ( 
.A1(n_2298),
.A2(n_2206),
.B(n_2128),
.Y(n_2326)
);

A2O1A1Ixp33_ASAP7_75t_L g2327 ( 
.A1(n_2273),
.A2(n_2244),
.B(n_2201),
.C(n_2250),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2279),
.B(n_2226),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2269),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2271),
.B(n_2266),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2286),
.Y(n_2331)
);

OR2x2_ASAP7_75t_L g2332 ( 
.A(n_2288),
.B(n_2079),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2271),
.B(n_2267),
.Y(n_2333)
);

A2O1A1Ixp33_ASAP7_75t_L g2334 ( 
.A1(n_2290),
.A2(n_2250),
.B(n_2220),
.C(n_2135),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_2285),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2288),
.Y(n_2336)
);

AOI21xp5_ASAP7_75t_L g2337 ( 
.A1(n_2291),
.A2(n_2196),
.B(n_2094),
.Y(n_2337)
);

AOI21xp5_ASAP7_75t_SL g2338 ( 
.A1(n_2296),
.A2(n_2196),
.B(n_2228),
.Y(n_2338)
);

AOI22xp33_ASAP7_75t_L g2339 ( 
.A1(n_2322),
.A2(n_2302),
.B1(n_2292),
.B2(n_2272),
.Y(n_2339)
);

AOI21xp5_ASAP7_75t_L g2340 ( 
.A1(n_2322),
.A2(n_2319),
.B(n_2327),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2331),
.Y(n_2341)
);

CKINVDCx8_ASAP7_75t_R g2342 ( 
.A(n_2335),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2317),
.B(n_2263),
.Y(n_2343)
);

OR2x6_ASAP7_75t_L g2344 ( 
.A(n_2338),
.B(n_2280),
.Y(n_2344)
);

INVxp33_ASAP7_75t_SL g2345 ( 
.A(n_2316),
.Y(n_2345)
);

INVx4_ASAP7_75t_L g2346 ( 
.A(n_2335),
.Y(n_2346)
);

HB1xp67_ASAP7_75t_L g2347 ( 
.A(n_2313),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2331),
.Y(n_2348)
);

CKINVDCx11_ASAP7_75t_R g2349 ( 
.A(n_2335),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2341),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2346),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2344),
.B(n_2317),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2348),
.Y(n_2353)
);

HB1xp67_ASAP7_75t_L g2354 ( 
.A(n_2347),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2345),
.Y(n_2355)
);

AO21x2_ASAP7_75t_L g2356 ( 
.A1(n_2340),
.A2(n_2337),
.B(n_2338),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2344),
.B(n_2313),
.Y(n_2357)
);

NOR2xp33_ASAP7_75t_L g2358 ( 
.A(n_2346),
.B(n_2335),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2350),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2355),
.B(n_2351),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2350),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2356),
.B(n_2344),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2353),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2354),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2353),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2356),
.B(n_2344),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2354),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2352),
.B(n_2346),
.Y(n_2368)
);

AOI22xp33_ASAP7_75t_L g2369 ( 
.A1(n_2362),
.A2(n_2339),
.B1(n_2320),
.B2(n_2300),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2368),
.B(n_2358),
.Y(n_2370)
);

OAI33xp33_ASAP7_75t_L g2371 ( 
.A1(n_2367),
.A2(n_2357),
.A3(n_2320),
.B1(n_2312),
.B2(n_2314),
.B3(n_2325),
.Y(n_2371)
);

OAI211xp5_ASAP7_75t_L g2372 ( 
.A1(n_2362),
.A2(n_2342),
.B(n_2358),
.C(n_2349),
.Y(n_2372)
);

AOI22xp33_ASAP7_75t_L g2373 ( 
.A1(n_2366),
.A2(n_2275),
.B1(n_2349),
.B2(n_2272),
.Y(n_2373)
);

AOI222xp33_ASAP7_75t_SL g2374 ( 
.A1(n_2364),
.A2(n_2345),
.B1(n_2264),
.B2(n_2315),
.C1(n_2335),
.C2(n_2323),
.Y(n_2374)
);

OAI211xp5_ASAP7_75t_SL g2375 ( 
.A1(n_2360),
.A2(n_2359),
.B(n_2361),
.C(n_2318),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2368),
.Y(n_2376)
);

AOI222xp33_ASAP7_75t_L g2377 ( 
.A1(n_2366),
.A2(n_2334),
.B1(n_2302),
.B2(n_2304),
.C1(n_2295),
.C2(n_2243),
.Y(n_2377)
);

OAI31xp33_ASAP7_75t_L g2378 ( 
.A1(n_2361),
.A2(n_2304),
.A3(n_2281),
.B(n_2343),
.Y(n_2378)
);

OAI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_2363),
.A2(n_2284),
.B1(n_2294),
.B2(n_2274),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2363),
.B(n_2321),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2370),
.B(n_2365),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2376),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2372),
.B(n_2365),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2369),
.B(n_2330),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2380),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2375),
.Y(n_2386)
);

INVx1_ASAP7_75t_SL g2387 ( 
.A(n_2379),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2369),
.B(n_2333),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2373),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2382),
.B(n_2373),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2381),
.Y(n_2391)
);

OR2x2_ASAP7_75t_L g2392 ( 
.A(n_2388),
.B(n_2378),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2388),
.B(n_2371),
.Y(n_2393)
);

OAI21xp33_ASAP7_75t_SL g2394 ( 
.A1(n_2393),
.A2(n_2386),
.B(n_2389),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2391),
.B(n_2381),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2390),
.Y(n_2396)
);

NOR2xp67_ASAP7_75t_L g2397 ( 
.A(n_2392),
.B(n_2383),
.Y(n_2397)
);

OAI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2397),
.A2(n_2384),
.B1(n_2387),
.B2(n_2383),
.Y(n_2398)
);

INVx1_ASAP7_75t_SL g2399 ( 
.A(n_2395),
.Y(n_2399)
);

AOI32xp33_ASAP7_75t_L g2400 ( 
.A1(n_2394),
.A2(n_2385),
.A3(n_2374),
.B1(n_2377),
.B2(n_2169),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_2395),
.B(n_2299),
.Y(n_2401)
);

AOI211xp5_ASAP7_75t_L g2402 ( 
.A1(n_2396),
.A2(n_2249),
.B(n_2256),
.C(n_2245),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2395),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2403),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2399),
.B(n_2295),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_SL g2406 ( 
.A(n_2398),
.B(n_2276),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_2401),
.Y(n_2407)
);

INVx1_ASAP7_75t_SL g2408 ( 
.A(n_2400),
.Y(n_2408)
);

AOI22xp33_ASAP7_75t_L g2409 ( 
.A1(n_2402),
.A2(n_2294),
.B1(n_2274),
.B2(n_2284),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2401),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2399),
.B(n_2285),
.Y(n_2411)
);

BUFx2_ASAP7_75t_L g2412 ( 
.A(n_2401),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2399),
.B(n_2085),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2406),
.A2(n_2277),
.B1(n_2307),
.B2(n_2294),
.Y(n_2414)
);

INVxp67_ASAP7_75t_SL g2415 ( 
.A(n_2405),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2408),
.A2(n_2277),
.B1(n_2307),
.B2(n_2274),
.Y(n_2416)
);

INVxp33_ASAP7_75t_L g2417 ( 
.A(n_2411),
.Y(n_2417)
);

OAI32xp33_ASAP7_75t_L g2418 ( 
.A1(n_2404),
.A2(n_2170),
.A3(n_2306),
.B1(n_2126),
.B2(n_2239),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_2412),
.A2(n_2119),
.B(n_2245),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2410),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2407),
.B(n_2311),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2413),
.B(n_2310),
.Y(n_2422)
);

OAI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2409),
.A2(n_2284),
.B1(n_2310),
.B2(n_2303),
.Y(n_2423)
);

OAI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_2411),
.A2(n_2256),
.B(n_2249),
.Y(n_2424)
);

OAI22xp33_ASAP7_75t_L g2425 ( 
.A1(n_2406),
.A2(n_2284),
.B1(n_2254),
.B2(n_2170),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2411),
.B(n_2293),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2420),
.B(n_2336),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2415),
.Y(n_2428)
);

NAND3x2_ASAP7_75t_L g2429 ( 
.A(n_2421),
.B(n_2076),
.C(n_2255),
.Y(n_2429)
);

AOI22xp33_ASAP7_75t_L g2430 ( 
.A1(n_2417),
.A2(n_2426),
.B1(n_2422),
.B2(n_2423),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2416),
.B(n_2336),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2419),
.B(n_2321),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2418),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_2425),
.A2(n_2254),
.B1(n_2174),
.B2(n_2151),
.Y(n_2434)
);

OAI32xp33_ASAP7_75t_L g2435 ( 
.A1(n_2424),
.A2(n_2253),
.A3(n_2332),
.B1(n_2308),
.B2(n_2305),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2414),
.B(n_2293),
.Y(n_2436)
);

INVx1_ASAP7_75t_SL g2437 ( 
.A(n_2421),
.Y(n_2437)
);

OAI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2416),
.A2(n_2091),
.B(n_2101),
.Y(n_2438)
);

CKINVDCx5p33_ASAP7_75t_R g2439 ( 
.A(n_2420),
.Y(n_2439)
);

OAI322xp33_ASAP7_75t_L g2440 ( 
.A1(n_2416),
.A2(n_2332),
.A3(n_148),
.B1(n_145),
.B2(n_147),
.C1(n_143),
.C2(n_144),
.Y(n_2440)
);

NOR2xp33_ASAP7_75t_L g2441 ( 
.A(n_2417),
.B(n_144),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2437),
.B(n_2439),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2441),
.B(n_2324),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2428),
.Y(n_2444)
);

HB1xp67_ASAP7_75t_L g2445 ( 
.A(n_2436),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2433),
.B(n_2324),
.Y(n_2446)
);

HB1xp67_ASAP7_75t_SL g2447 ( 
.A(n_2430),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2431),
.B(n_2432),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2427),
.B(n_2328),
.Y(n_2449)
);

INVx1_ASAP7_75t_SL g2450 ( 
.A(n_2440),
.Y(n_2450)
);

BUFx2_ASAP7_75t_L g2451 ( 
.A(n_2429),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_2438),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2435),
.B(n_2434),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2434),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2437),
.B(n_2328),
.Y(n_2455)
);

OAI221xp5_ASAP7_75t_SL g2456 ( 
.A1(n_2450),
.A2(n_2253),
.B1(n_2326),
.B2(n_2329),
.C(n_147),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2450),
.B(n_145),
.Y(n_2457)
);

O2A1O1Ixp5_ASAP7_75t_L g2458 ( 
.A1(n_2442),
.A2(n_2072),
.B(n_2329),
.C(n_150),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2455),
.B(n_146),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_SL g2460 ( 
.A(n_2445),
.B(n_2254),
.Y(n_2460)
);

NOR2x1_ASAP7_75t_L g2461 ( 
.A(n_2444),
.B(n_149),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2447),
.Y(n_2462)
);

NOR2x1_ASAP7_75t_L g2463 ( 
.A(n_2451),
.B(n_2454),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2446),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_2453),
.B(n_2226),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2448),
.Y(n_2466)
);

NOR3xp33_ASAP7_75t_L g2467 ( 
.A(n_2452),
.B(n_150),
.C(n_151),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2449),
.B(n_152),
.Y(n_2468)
);

AOI221xp5_ASAP7_75t_L g2469 ( 
.A1(n_2443),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.C(n_155),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2450),
.B(n_153),
.Y(n_2470)
);

NAND3xp33_ASAP7_75t_L g2471 ( 
.A(n_2445),
.B(n_154),
.C(n_155),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2455),
.B(n_2309),
.Y(n_2472)
);

AOI21xp5_ASAP7_75t_L g2473 ( 
.A1(n_2442),
.A2(n_2078),
.B(n_156),
.Y(n_2473)
);

NAND3xp33_ASAP7_75t_SL g2474 ( 
.A(n_2450),
.B(n_157),
.C(n_158),
.Y(n_2474)
);

NAND3xp33_ASAP7_75t_L g2475 ( 
.A(n_2445),
.B(n_157),
.C(n_159),
.Y(n_2475)
);

NOR3x1_ASAP7_75t_L g2476 ( 
.A(n_2451),
.B(n_159),
.C(n_160),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2455),
.Y(n_2477)
);

NAND4xp25_ASAP7_75t_L g2478 ( 
.A(n_2476),
.B(n_163),
.C(n_160),
.D(n_161),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2474),
.B(n_161),
.Y(n_2479)
);

NAND3xp33_ASAP7_75t_L g2480 ( 
.A(n_2461),
.B(n_164),
.C(n_165),
.Y(n_2480)
);

AOI21xp5_ASAP7_75t_L g2481 ( 
.A1(n_2457),
.A2(n_164),
.B(n_165),
.Y(n_2481)
);

NOR3xp33_ASAP7_75t_L g2482 ( 
.A(n_2462),
.B(n_166),
.C(n_167),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2470),
.Y(n_2483)
);

NOR4xp25_ASAP7_75t_L g2484 ( 
.A(n_2466),
.B(n_2477),
.C(n_2464),
.D(n_2465),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2459),
.Y(n_2485)
);

OR2x2_ASAP7_75t_L g2486 ( 
.A(n_2468),
.B(n_166),
.Y(n_2486)
);

NOR3xp33_ASAP7_75t_L g2487 ( 
.A(n_2463),
.B(n_167),
.C(n_168),
.Y(n_2487)
);

AOI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_2471),
.A2(n_168),
.B(n_169),
.Y(n_2488)
);

NAND4xp25_ASAP7_75t_L g2489 ( 
.A(n_2460),
.B(n_171),
.C(n_169),
.D(n_170),
.Y(n_2489)
);

OAI211xp5_ASAP7_75t_L g2490 ( 
.A1(n_2475),
.A2(n_173),
.B(n_170),
.C(n_171),
.Y(n_2490)
);

NOR3x1_ASAP7_75t_L g2491 ( 
.A(n_2467),
.B(n_173),
.C(n_174),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2472),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2469),
.Y(n_2493)
);

AND4x1_ASAP7_75t_L g2494 ( 
.A(n_2458),
.B(n_176),
.C(n_174),
.D(n_175),
.Y(n_2494)
);

NAND3xp33_ASAP7_75t_SL g2495 ( 
.A(n_2473),
.B(n_175),
.C(n_176),
.Y(n_2495)
);

OAI211xp5_ASAP7_75t_L g2496 ( 
.A1(n_2456),
.A2(n_179),
.B(n_177),
.C(n_178),
.Y(n_2496)
);

NAND4xp75_ASAP7_75t_L g2497 ( 
.A(n_2476),
.B(n_180),
.C(n_177),
.D(n_179),
.Y(n_2497)
);

OR3x1_ASAP7_75t_L g2498 ( 
.A(n_2474),
.B(n_180),
.C(n_181),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_L g2499 ( 
.A(n_2474),
.B(n_181),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2472),
.B(n_182),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2472),
.B(n_184),
.Y(n_2501)
);

INVxp67_ASAP7_75t_SL g2502 ( 
.A(n_2461),
.Y(n_2502)
);

AOI211xp5_ASAP7_75t_L g2503 ( 
.A1(n_2474),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_2503)
);

BUFx4f_ASAP7_75t_SL g2504 ( 
.A(n_2462),
.Y(n_2504)
);

INVxp67_ASAP7_75t_L g2505 ( 
.A(n_2460),
.Y(n_2505)
);

AOI221xp5_ASAP7_75t_L g2506 ( 
.A1(n_2474),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_2506)
);

INVx2_ASAP7_75t_SL g2507 ( 
.A(n_2461),
.Y(n_2507)
);

OR2x2_ASAP7_75t_L g2508 ( 
.A(n_2457),
.B(n_187),
.Y(n_2508)
);

NOR4xp25_ASAP7_75t_L g2509 ( 
.A(n_2474),
.B(n_190),
.C(n_188),
.D(n_189),
.Y(n_2509)
);

AOI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2462),
.A2(n_2252),
.B1(n_2278),
.B2(n_2069),
.Y(n_2510)
);

INVx1_ASAP7_75t_SL g2511 ( 
.A(n_2461),
.Y(n_2511)
);

NOR4xp25_ASAP7_75t_SL g2512 ( 
.A(n_2462),
.B(n_194),
.C(n_191),
.D(n_193),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2461),
.Y(n_2513)
);

INVx2_ASAP7_75t_SL g2514 ( 
.A(n_2461),
.Y(n_2514)
);

NAND3xp33_ASAP7_75t_L g2515 ( 
.A(n_2503),
.B(n_2487),
.C(n_2506),
.Y(n_2515)
);

OAI221xp5_ASAP7_75t_L g2516 ( 
.A1(n_2509),
.A2(n_194),
.B1(n_191),
.B2(n_193),
.C(n_195),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2500),
.B(n_2507),
.Y(n_2517)
);

AOI22xp5_ASAP7_75t_L g2518 ( 
.A1(n_2504),
.A2(n_2252),
.B1(n_2278),
.B2(n_2158),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2498),
.Y(n_2519)
);

NOR3xp33_ASAP7_75t_L g2520 ( 
.A(n_2485),
.B(n_195),
.C(n_196),
.Y(n_2520)
);

NAND3xp33_ASAP7_75t_SL g2521 ( 
.A(n_2512),
.B(n_196),
.C(n_197),
.Y(n_2521)
);

NOR2x1_ASAP7_75t_L g2522 ( 
.A(n_2480),
.B(n_197),
.Y(n_2522)
);

OAI21xp33_ASAP7_75t_L g2523 ( 
.A1(n_2484),
.A2(n_2087),
.B(n_198),
.Y(n_2523)
);

O2A1O1Ixp33_ASAP7_75t_L g2524 ( 
.A1(n_2514),
.A2(n_201),
.B(n_199),
.C(n_200),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2479),
.B(n_199),
.Y(n_2525)
);

NOR4xp75_ASAP7_75t_L g2526 ( 
.A(n_2497),
.B(n_203),
.C(n_200),
.D(n_202),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2499),
.B(n_203),
.Y(n_2527)
);

NAND3xp33_ASAP7_75t_SL g2528 ( 
.A(n_2511),
.B(n_204),
.C(n_206),
.Y(n_2528)
);

AOI221xp5_ASAP7_75t_L g2529 ( 
.A1(n_2505),
.A2(n_2502),
.B1(n_2513),
.B2(n_2496),
.C(n_2495),
.Y(n_2529)
);

AOI211xp5_ASAP7_75t_L g2530 ( 
.A1(n_2490),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_2530)
);

NAND4xp25_ASAP7_75t_L g2531 ( 
.A(n_2492),
.B(n_210),
.C(n_207),
.D(n_209),
.Y(n_2531)
);

O2A1O1Ixp33_ASAP7_75t_L g2532 ( 
.A1(n_2501),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_2532)
);

AOI22xp33_ASAP7_75t_L g2533 ( 
.A1(n_2483),
.A2(n_2278),
.B1(n_2150),
.B2(n_213),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2482),
.B(n_211),
.Y(n_2534)
);

NAND3xp33_ASAP7_75t_L g2535 ( 
.A(n_2478),
.B(n_212),
.C(n_213),
.Y(n_2535)
);

XNOR2xp5_ASAP7_75t_L g2536 ( 
.A(n_2494),
.B(n_212),
.Y(n_2536)
);

AOI211xp5_ASAP7_75t_L g2537 ( 
.A1(n_2488),
.A2(n_217),
.B(n_214),
.C(n_216),
.Y(n_2537)
);

OAI21xp33_ASAP7_75t_SL g2538 ( 
.A1(n_2493),
.A2(n_216),
.B(n_217),
.Y(n_2538)
);

AOI211xp5_ASAP7_75t_L g2539 ( 
.A1(n_2489),
.A2(n_221),
.B(n_218),
.C(n_220),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2491),
.B(n_218),
.Y(n_2540)
);

NAND4xp75_ASAP7_75t_L g2541 ( 
.A(n_2481),
.B(n_224),
.C(n_222),
.D(n_223),
.Y(n_2541)
);

AND3x1_ASAP7_75t_L g2542 ( 
.A(n_2485),
.B(n_2508),
.C(n_2486),
.Y(n_2542)
);

NAND3x1_ASAP7_75t_L g2543 ( 
.A(n_2510),
.B(n_222),
.C(n_224),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_SL g2544 ( 
.A(n_2497),
.B(n_225),
.Y(n_2544)
);

AOI211xp5_ASAP7_75t_L g2545 ( 
.A1(n_2509),
.A2(n_228),
.B(n_225),
.C(n_227),
.Y(n_2545)
);

NAND4xp75_ASAP7_75t_L g2546 ( 
.A(n_2491),
.B(n_229),
.C(n_227),
.D(n_228),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2500),
.B(n_229),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2500),
.B(n_230),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2500),
.B(n_230),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2502),
.A2(n_231),
.B(n_232),
.Y(n_2550)
);

NOR3xp33_ASAP7_75t_SL g2551 ( 
.A(n_2496),
.B(n_231),
.C(n_232),
.Y(n_2551)
);

NOR3xp33_ASAP7_75t_L g2552 ( 
.A(n_2485),
.B(n_233),
.C(n_234),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2546),
.Y(n_2553)
);

NAND3xp33_ASAP7_75t_L g2554 ( 
.A(n_2537),
.B(n_234),
.C(n_235),
.Y(n_2554)
);

NAND4xp75_ASAP7_75t_L g2555 ( 
.A(n_2529),
.B(n_237),
.C(n_235),
.D(n_236),
.Y(n_2555)
);

AOI221x1_ASAP7_75t_L g2556 ( 
.A1(n_2525),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.C(n_239),
.Y(n_2556)
);

AOI21xp5_ASAP7_75t_L g2557 ( 
.A1(n_2517),
.A2(n_239),
.B(n_240),
.Y(n_2557)
);

OAI211xp5_ASAP7_75t_SL g2558 ( 
.A1(n_2551),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2540),
.B(n_241),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2535),
.A2(n_2065),
.B1(n_245),
.B2(n_243),
.Y(n_2560)
);

NOR3xp33_ASAP7_75t_L g2561 ( 
.A(n_2527),
.B(n_243),
.C(n_244),
.Y(n_2561)
);

NAND4xp75_ASAP7_75t_L g2562 ( 
.A(n_2538),
.B(n_247),
.C(n_244),
.D(n_246),
.Y(n_2562)
);

NAND3xp33_ASAP7_75t_L g2563 ( 
.A(n_2545),
.B(n_2530),
.C(n_2544),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2536),
.B(n_247),
.Y(n_2564)
);

NOR2x1_ASAP7_75t_L g2565 ( 
.A(n_2521),
.B(n_248),
.Y(n_2565)
);

OAI21xp33_ASAP7_75t_L g2566 ( 
.A1(n_2519),
.A2(n_249),
.B(n_250),
.Y(n_2566)
);

AOI211xp5_ASAP7_75t_SL g2567 ( 
.A1(n_2516),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_2567)
);

OAI211xp5_ASAP7_75t_L g2568 ( 
.A1(n_2539),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_2568)
);

NAND3xp33_ASAP7_75t_L g2569 ( 
.A(n_2524),
.B(n_254),
.C(n_255),
.Y(n_2569)
);

AOI211xp5_ASAP7_75t_L g2570 ( 
.A1(n_2528),
.A2(n_2515),
.B(n_2532),
.C(n_2534),
.Y(n_2570)
);

NOR3xp33_ASAP7_75t_L g2571 ( 
.A(n_2547),
.B(n_254),
.C(n_255),
.Y(n_2571)
);

AOI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2548),
.A2(n_256),
.B(n_257),
.Y(n_2572)
);

AOI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2542),
.A2(n_2278),
.B1(n_261),
.B2(n_256),
.Y(n_2573)
);

OAI221xp5_ASAP7_75t_L g2574 ( 
.A1(n_2523),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.C(n_263),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2549),
.Y(n_2575)
);

NOR2xp33_ASAP7_75t_L g2576 ( 
.A(n_2531),
.B(n_262),
.Y(n_2576)
);

AOI221xp5_ASAP7_75t_L g2577 ( 
.A1(n_2550),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_266),
.Y(n_2577)
);

NAND5xp2_ASAP7_75t_L g2578 ( 
.A(n_2520),
.B(n_266),
.C(n_264),
.D(n_265),
.E(n_267),
.Y(n_2578)
);

OAI211xp5_ASAP7_75t_L g2579 ( 
.A1(n_2522),
.A2(n_270),
.B(n_268),
.C(n_269),
.Y(n_2579)
);

NOR3xp33_ASAP7_75t_L g2580 ( 
.A(n_2541),
.B(n_268),
.C(n_269),
.Y(n_2580)
);

OAI221xp5_ASAP7_75t_L g2581 ( 
.A1(n_2552),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.C(n_273),
.Y(n_2581)
);

NAND3xp33_ASAP7_75t_L g2582 ( 
.A(n_2533),
.B(n_272),
.C(n_274),
.Y(n_2582)
);

AND3x4_ASAP7_75t_L g2583 ( 
.A(n_2526),
.B(n_274),
.C(n_275),
.Y(n_2583)
);

OAI211xp5_ASAP7_75t_L g2584 ( 
.A1(n_2518),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_2584)
);

AOI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_2543),
.A2(n_276),
.B(n_277),
.Y(n_2585)
);

AOI221x1_ASAP7_75t_L g2586 ( 
.A1(n_2525),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.C(n_281),
.Y(n_2586)
);

OAI21xp5_ASAP7_75t_SL g2587 ( 
.A1(n_2536),
.A2(n_278),
.B(n_280),
.Y(n_2587)
);

NAND4xp25_ASAP7_75t_SL g2588 ( 
.A(n_2529),
.B(n_283),
.C(n_281),
.D(n_282),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2536),
.Y(n_2589)
);

AOI221xp5_ASAP7_75t_L g2590 ( 
.A1(n_2521),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.C(n_285),
.Y(n_2590)
);

NAND2x1p5_ASAP7_75t_L g2591 ( 
.A(n_2542),
.B(n_284),
.Y(n_2591)
);

NAND3xp33_ASAP7_75t_SL g2592 ( 
.A(n_2545),
.B(n_285),
.C(n_286),
.Y(n_2592)
);

INVx3_ASAP7_75t_SL g2593 ( 
.A(n_2540),
.Y(n_2593)
);

OAI211xp5_ASAP7_75t_L g2594 ( 
.A1(n_2538),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_2594)
);

AOI211xp5_ASAP7_75t_L g2595 ( 
.A1(n_2521),
.A2(n_290),
.B(n_287),
.C(n_289),
.Y(n_2595)
);

AOI211xp5_ASAP7_75t_L g2596 ( 
.A1(n_2521),
.A2(n_292),
.B(n_290),
.C(n_291),
.Y(n_2596)
);

A2O1A1Ixp33_ASAP7_75t_L g2597 ( 
.A1(n_2524),
.A2(n_294),
.B(n_291),
.C(n_293),
.Y(n_2597)
);

AOI211xp5_ASAP7_75t_L g2598 ( 
.A1(n_2521),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_SL g2599 ( 
.A(n_2545),
.B(n_295),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2536),
.Y(n_2600)
);

NOR4xp25_ASAP7_75t_L g2601 ( 
.A(n_2521),
.B(n_299),
.C(n_296),
.D(n_297),
.Y(n_2601)
);

AOI221xp5_ASAP7_75t_L g2602 ( 
.A1(n_2521),
.A2(n_301),
.B1(n_297),
.B2(n_300),
.C(n_302),
.Y(n_2602)
);

AOI221xp5_ASAP7_75t_SL g2603 ( 
.A1(n_2529),
.A2(n_303),
.B1(n_300),
.B2(n_302),
.C(n_304),
.Y(n_2603)
);

NOR5xp2_ASAP7_75t_L g2604 ( 
.A(n_2516),
.B(n_306),
.C(n_303),
.D(n_305),
.E(n_307),
.Y(n_2604)
);

AOI211xp5_ASAP7_75t_L g2605 ( 
.A1(n_2521),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_2605)
);

NAND4xp25_ASAP7_75t_L g2606 ( 
.A(n_2529),
.B(n_311),
.C(n_309),
.D(n_310),
.Y(n_2606)
);

AOI221xp5_ASAP7_75t_L g2607 ( 
.A1(n_2521),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.C(n_316),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2536),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2540),
.B(n_312),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2540),
.B(n_314),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2536),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2540),
.B(n_316),
.Y(n_2612)
);

NOR4xp75_ASAP7_75t_L g2613 ( 
.A(n_2521),
.B(n_320),
.C(n_317),
.D(n_318),
.Y(n_2613)
);

AOI211xp5_ASAP7_75t_L g2614 ( 
.A1(n_2521),
.A2(n_321),
.B(n_317),
.C(n_320),
.Y(n_2614)
);

OAI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2573),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_2615)
);

BUFx2_ASAP7_75t_L g2616 ( 
.A(n_2591),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2612),
.B(n_322),
.Y(n_2617)
);

AOI211xp5_ASAP7_75t_L g2618 ( 
.A1(n_2601),
.A2(n_325),
.B(n_323),
.C(n_324),
.Y(n_2618)
);

OAI222xp33_ASAP7_75t_L g2619 ( 
.A1(n_2565),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.C1(n_329),
.C2(n_330),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_L g2620 ( 
.A(n_2606),
.B(n_326),
.Y(n_2620)
);

AND2x4_ASAP7_75t_L g2621 ( 
.A(n_2613),
.B(n_327),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2593),
.B(n_328),
.Y(n_2622)
);

NAND3xp33_ASAP7_75t_L g2623 ( 
.A(n_2595),
.B(n_329),
.C(n_330),
.Y(n_2623)
);

OA21x2_ASAP7_75t_L g2624 ( 
.A1(n_2589),
.A2(n_331),
.B(n_332),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2562),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2566),
.B(n_332),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_R g2627 ( 
.A(n_2588),
.B(n_333),
.Y(n_2627)
);

HB1xp67_ASAP7_75t_L g2628 ( 
.A(n_2583),
.Y(n_2628)
);

A2O1A1Ixp33_ASAP7_75t_SL g2629 ( 
.A1(n_2600),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_2629)
);

NOR3xp33_ASAP7_75t_L g2630 ( 
.A(n_2564),
.B(n_334),
.C(n_335),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2555),
.Y(n_2631)
);

AOI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2559),
.A2(n_2610),
.B(n_2609),
.Y(n_2632)
);

OR2x2_ASAP7_75t_L g2633 ( 
.A(n_2578),
.B(n_336),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2580),
.A2(n_2278),
.B1(n_338),
.B2(n_336),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2566),
.B(n_337),
.Y(n_2635)
);

NOR3xp33_ASAP7_75t_L g2636 ( 
.A(n_2587),
.B(n_338),
.C(n_340),
.Y(n_2636)
);

AOI211xp5_ASAP7_75t_L g2637 ( 
.A1(n_2574),
.A2(n_342),
.B(n_340),
.C(n_341),
.Y(n_2637)
);

OAI221xp5_ASAP7_75t_L g2638 ( 
.A1(n_2590),
.A2(n_345),
.B1(n_341),
.B2(n_344),
.C(n_346),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2553),
.B(n_344),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2603),
.B(n_345),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2594),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2569),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2596),
.B(n_346),
.Y(n_2643)
);

NOR2x1_ASAP7_75t_SL g2644 ( 
.A(n_2579),
.B(n_348),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2598),
.B(n_348),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2576),
.Y(n_2646)
);

NAND3xp33_ASAP7_75t_L g2647 ( 
.A(n_2605),
.B(n_349),
.C(n_350),
.Y(n_2647)
);

OAI211xp5_ASAP7_75t_L g2648 ( 
.A1(n_2602),
.A2(n_353),
.B(n_349),
.C(n_351),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2614),
.B(n_351),
.Y(n_2649)
);

AOI221xp5_ASAP7_75t_L g2650 ( 
.A1(n_2607),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.C(n_356),
.Y(n_2650)
);

AOI221xp5_ASAP7_75t_L g2651 ( 
.A1(n_2558),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.C(n_358),
.Y(n_2651)
);

AOI221xp5_ASAP7_75t_L g2652 ( 
.A1(n_2592),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.C(n_361),
.Y(n_2652)
);

INVx1_ASAP7_75t_SL g2653 ( 
.A(n_2585),
.Y(n_2653)
);

AOI22xp5_ASAP7_75t_SL g2654 ( 
.A1(n_2557),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_2654)
);

AOI321xp33_ASAP7_75t_L g2655 ( 
.A1(n_2570),
.A2(n_362),
.A3(n_363),
.B1(n_364),
.B2(n_365),
.C(n_366),
.Y(n_2655)
);

NOR3xp33_ASAP7_75t_L g2656 ( 
.A(n_2563),
.B(n_364),
.C(n_365),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2567),
.B(n_366),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_R g2658 ( 
.A(n_2608),
.B(n_367),
.Y(n_2658)
);

HB1xp67_ASAP7_75t_L g2659 ( 
.A(n_2556),
.Y(n_2659)
);

HB1xp67_ASAP7_75t_L g2660 ( 
.A(n_2586),
.Y(n_2660)
);

AOI211xp5_ASAP7_75t_L g2661 ( 
.A1(n_2568),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_2661)
);

O2A1O1Ixp33_ASAP7_75t_L g2662 ( 
.A1(n_2597),
.A2(n_370),
.B(n_368),
.C(n_369),
.Y(n_2662)
);

OR2x2_ASAP7_75t_L g2663 ( 
.A(n_2554),
.B(n_370),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2571),
.B(n_371),
.Y(n_2664)
);

OAI222xp33_ASAP7_75t_L g2665 ( 
.A1(n_2599),
.A2(n_2611),
.B1(n_2560),
.B2(n_2575),
.C1(n_2581),
.C2(n_2572),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2582),
.Y(n_2666)
);

NAND2xp33_ASAP7_75t_R g2667 ( 
.A(n_2604),
.B(n_371),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_2577),
.B(n_372),
.Y(n_2668)
);

NOR2x1_ASAP7_75t_L g2669 ( 
.A(n_2584),
.B(n_372),
.Y(n_2669)
);

OAI21xp5_ASAP7_75t_L g2670 ( 
.A1(n_2561),
.A2(n_373),
.B(n_374),
.Y(n_2670)
);

A2O1A1Ixp33_ASAP7_75t_SL g2671 ( 
.A1(n_2589),
.A2(n_377),
.B(n_374),
.C(n_376),
.Y(n_2671)
);

NAND3xp33_ASAP7_75t_SL g2672 ( 
.A(n_2595),
.B(n_377),
.C(n_378),
.Y(n_2672)
);

AOI221xp5_ASAP7_75t_L g2673 ( 
.A1(n_2601),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.C(n_381),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2591),
.Y(n_2674)
);

OAI222xp33_ASAP7_75t_L g2675 ( 
.A1(n_2565),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.C1(n_384),
.C2(n_385),
.Y(n_2675)
);

AOI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2564),
.A2(n_382),
.B(n_383),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2580),
.A2(n_2278),
.B1(n_386),
.B2(n_384),
.Y(n_2677)
);

AND2x2_ASAP7_75t_L g2678 ( 
.A(n_2612),
.B(n_385),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_R g2679 ( 
.A(n_2588),
.B(n_386),
.Y(n_2679)
);

OAI221xp5_ASAP7_75t_L g2680 ( 
.A1(n_2601),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.C(n_390),
.Y(n_2680)
);

NAND4xp75_ASAP7_75t_L g2681 ( 
.A(n_2565),
.B(n_390),
.C(n_388),
.D(n_389),
.Y(n_2681)
);

NAND4xp75_ASAP7_75t_L g2682 ( 
.A(n_2639),
.B(n_2625),
.C(n_2641),
.D(n_2669),
.Y(n_2682)
);

NOR2x1p5_ASAP7_75t_L g2683 ( 
.A(n_2681),
.B(n_391),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2678),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2633),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2621),
.A2(n_2620),
.B1(n_2667),
.B2(n_2636),
.Y(n_2686)
);

HB1xp67_ASAP7_75t_L g2687 ( 
.A(n_2624),
.Y(n_2687)
);

NOR2x1p5_ASAP7_75t_L g2688 ( 
.A(n_2672),
.B(n_391),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2621),
.B(n_392),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2617),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2622),
.B(n_392),
.Y(n_2691)
);

OR2x2_ASAP7_75t_L g2692 ( 
.A(n_2626),
.B(n_393),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2635),
.B(n_394),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2659),
.Y(n_2694)
);

AOI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2656),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_2695)
);

OR2x6_ASAP7_75t_L g2696 ( 
.A(n_2674),
.B(n_396),
.Y(n_2696)
);

NAND4xp75_ASAP7_75t_L g2697 ( 
.A(n_2642),
.B(n_399),
.C(n_397),
.D(n_398),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2660),
.Y(n_2698)
);

NOR2x1p5_ASAP7_75t_L g2699 ( 
.A(n_2657),
.B(n_398),
.Y(n_2699)
);

NOR4xp75_ASAP7_75t_L g2700 ( 
.A(n_2640),
.B(n_2668),
.C(n_2645),
.D(n_2649),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2644),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2624),
.Y(n_2702)
);

OAI221xp5_ASAP7_75t_L g2703 ( 
.A1(n_2673),
.A2(n_2671),
.B1(n_2629),
.B2(n_2677),
.C(n_2634),
.Y(n_2703)
);

AND2x4_ASAP7_75t_L g2704 ( 
.A(n_2616),
.B(n_399),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2628),
.Y(n_2705)
);

NOR2xp33_ASAP7_75t_L g2706 ( 
.A(n_2680),
.B(n_400),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2654),
.Y(n_2707)
);

AO22x2_ASAP7_75t_L g2708 ( 
.A1(n_2653),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_2708)
);

AOI22xp5_ASAP7_75t_L g2709 ( 
.A1(n_2630),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_2709)
);

INVx1_ASAP7_75t_SL g2710 ( 
.A(n_2658),
.Y(n_2710)
);

NOR2xp33_ASAP7_75t_L g2711 ( 
.A(n_2619),
.B(n_404),
.Y(n_2711)
);

NOR2x1_ASAP7_75t_L g2712 ( 
.A(n_2675),
.B(n_405),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2643),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2663),
.Y(n_2714)
);

NAND4xp75_ASAP7_75t_L g2715 ( 
.A(n_2676),
.B(n_408),
.C(n_406),
.D(n_407),
.Y(n_2715)
);

NOR2x1p5_ASAP7_75t_L g2716 ( 
.A(n_2631),
.B(n_407),
.Y(n_2716)
);

NOR2x1_ASAP7_75t_L g2717 ( 
.A(n_2631),
.B(n_408),
.Y(n_2717)
);

NOR2x1_ASAP7_75t_L g2718 ( 
.A(n_2623),
.B(n_409),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2664),
.Y(n_2719)
);

AND3x4_ASAP7_75t_L g2720 ( 
.A(n_2666),
.B(n_410),
.C(n_411),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2647),
.Y(n_2721)
);

AOI22xp5_ASAP7_75t_L g2722 ( 
.A1(n_2651),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_2722)
);

NOR2x1_ASAP7_75t_L g2723 ( 
.A(n_2670),
.B(n_412),
.Y(n_2723)
);

XOR2xp5_ASAP7_75t_L g2724 ( 
.A(n_2615),
.B(n_413),
.Y(n_2724)
);

INVx3_ASAP7_75t_L g2725 ( 
.A(n_2646),
.Y(n_2725)
);

AOI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2648),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2662),
.Y(n_2727)
);

NAND2x1p5_ASAP7_75t_L g2728 ( 
.A(n_2632),
.B(n_415),
.Y(n_2728)
);

NAND4xp75_ASAP7_75t_L g2729 ( 
.A(n_2652),
.B(n_418),
.C(n_416),
.D(n_417),
.Y(n_2729)
);

INVxp67_ASAP7_75t_L g2730 ( 
.A(n_2638),
.Y(n_2730)
);

NOR2x1_ASAP7_75t_L g2731 ( 
.A(n_2665),
.B(n_417),
.Y(n_2731)
);

AOI22xp5_ASAP7_75t_SL g2732 ( 
.A1(n_2655),
.A2(n_2618),
.B1(n_2679),
.B2(n_2627),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2661),
.Y(n_2733)
);

INVxp33_ASAP7_75t_SL g2734 ( 
.A(n_2650),
.Y(n_2734)
);

AOI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2637),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2639),
.B(n_419),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2633),
.B(n_420),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2678),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2678),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2624),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2678),
.Y(n_2741)
);

NOR2x1_ASAP7_75t_L g2742 ( 
.A(n_2681),
.B(n_421),
.Y(n_2742)
);

AOI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2621),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2736),
.B(n_423),
.Y(n_2744)
);

AOI211xp5_ASAP7_75t_L g2745 ( 
.A1(n_2711),
.A2(n_426),
.B(n_424),
.C(n_425),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2689),
.B(n_424),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2687),
.Y(n_2747)
);

OR3x1_ASAP7_75t_L g2748 ( 
.A(n_2706),
.B(n_425),
.C(n_426),
.Y(n_2748)
);

NOR4xp25_ASAP7_75t_L g2749 ( 
.A(n_2694),
.B(n_429),
.C(n_427),
.D(n_428),
.Y(n_2749)
);

AOI211xp5_ASAP7_75t_L g2750 ( 
.A1(n_2703),
.A2(n_430),
.B(n_427),
.C(n_429),
.Y(n_2750)
);

AOI221xp5_ASAP7_75t_L g2751 ( 
.A1(n_2698),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.C(n_433),
.Y(n_2751)
);

AO211x2_ASAP7_75t_L g2752 ( 
.A1(n_2701),
.A2(n_431),
.B(n_432),
.C(n_433),
.Y(n_2752)
);

NAND4xp25_ASAP7_75t_L g2753 ( 
.A(n_2686),
.B(n_434),
.C(n_435),
.D(n_436),
.Y(n_2753)
);

OAI221xp5_ASAP7_75t_L g2754 ( 
.A1(n_2726),
.A2(n_434),
.B1(n_435),
.B2(n_437),
.C(n_438),
.Y(n_2754)
);

NAND3xp33_ASAP7_75t_L g2755 ( 
.A(n_2743),
.B(n_437),
.C(n_438),
.Y(n_2755)
);

NOR3xp33_ASAP7_75t_L g2756 ( 
.A(n_2705),
.B(n_439),
.C(n_440),
.Y(n_2756)
);

NAND5xp2_ASAP7_75t_L g2757 ( 
.A(n_2684),
.B(n_2738),
.C(n_2741),
.D(n_2739),
.E(n_2685),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2708),
.Y(n_2758)
);

NOR5xp2_ASAP7_75t_L g2759 ( 
.A(n_2730),
.B(n_439),
.C(n_440),
.D(n_441),
.E(n_442),
.Y(n_2759)
);

NAND4xp25_ASAP7_75t_L g2760 ( 
.A(n_2722),
.B(n_443),
.C(n_444),
.D(n_445),
.Y(n_2760)
);

NOR5xp2_ASAP7_75t_L g2761 ( 
.A(n_2702),
.B(n_443),
.C(n_444),
.D(n_445),
.E(n_446),
.Y(n_2761)
);

AOI21xp5_ASAP7_75t_L g2762 ( 
.A1(n_2740),
.A2(n_446),
.B(n_447),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2708),
.Y(n_2763)
);

AOI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2734),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.Y(n_2764)
);

NOR3xp33_ASAP7_75t_L g2765 ( 
.A(n_2682),
.B(n_450),
.C(n_452),
.Y(n_2765)
);

XNOR2xp5_ASAP7_75t_L g2766 ( 
.A(n_2720),
.B(n_452),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2728),
.Y(n_2767)
);

NAND3xp33_ASAP7_75t_SL g2768 ( 
.A(n_2710),
.B(n_453),
.C(n_454),
.Y(n_2768)
);

AOI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2707),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2696),
.Y(n_2770)
);

NOR4xp75_ASAP7_75t_L g2771 ( 
.A(n_2729),
.B(n_455),
.C(n_456),
.D(n_457),
.Y(n_2771)
);

XOR2xp5_ASAP7_75t_L g2772 ( 
.A(n_2732),
.B(n_457),
.Y(n_2772)
);

AO22x2_ASAP7_75t_L g2773 ( 
.A1(n_2737),
.A2(n_458),
.B1(n_459),
.B2(n_460),
.Y(n_2773)
);

AND2x4_ASAP7_75t_L g2774 ( 
.A(n_2716),
.B(n_460),
.Y(n_2774)
);

AND2x4_ASAP7_75t_L g2775 ( 
.A(n_2717),
.B(n_461),
.Y(n_2775)
);

NOR3xp33_ASAP7_75t_SL g2776 ( 
.A(n_2727),
.B(n_461),
.C(n_463),
.Y(n_2776)
);

NAND2x1p5_ASAP7_75t_L g2777 ( 
.A(n_2731),
.B(n_463),
.Y(n_2777)
);

NAND5xp2_ASAP7_75t_L g2778 ( 
.A(n_2733),
.B(n_464),
.C(n_465),
.D(n_467),
.E(n_468),
.Y(n_2778)
);

NAND5xp2_ASAP7_75t_L g2779 ( 
.A(n_2721),
.B(n_2714),
.C(n_2690),
.D(n_2713),
.E(n_2719),
.Y(n_2779)
);

OR2x2_ASAP7_75t_L g2780 ( 
.A(n_2691),
.B(n_2692),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2696),
.Y(n_2781)
);

NAND3xp33_ASAP7_75t_SL g2782 ( 
.A(n_2700),
.B(n_465),
.C(n_467),
.Y(n_2782)
);

HB1xp67_ASAP7_75t_L g2783 ( 
.A(n_2697),
.Y(n_2783)
);

NOR3xp33_ASAP7_75t_L g2784 ( 
.A(n_2725),
.B(n_469),
.C(n_470),
.Y(n_2784)
);

NOR3xp33_ASAP7_75t_L g2785 ( 
.A(n_2693),
.B(n_469),
.C(n_470),
.Y(n_2785)
);

NOR3xp33_ASAP7_75t_L g2786 ( 
.A(n_2723),
.B(n_471),
.C(n_472),
.Y(n_2786)
);

NOR3xp33_ASAP7_75t_L g2787 ( 
.A(n_2742),
.B(n_472),
.C(n_473),
.Y(n_2787)
);

CKINVDCx5p33_ASAP7_75t_R g2788 ( 
.A(n_2770),
.Y(n_2788)
);

INVxp33_ASAP7_75t_SL g2789 ( 
.A(n_2772),
.Y(n_2789)
);

CKINVDCx5p33_ASAP7_75t_R g2790 ( 
.A(n_2783),
.Y(n_2790)
);

BUFx2_ASAP7_75t_L g2791 ( 
.A(n_2775),
.Y(n_2791)
);

INVx3_ASAP7_75t_SL g2792 ( 
.A(n_2781),
.Y(n_2792)
);

BUFx2_ASAP7_75t_L g2793 ( 
.A(n_2775),
.Y(n_2793)
);

OAI21xp33_ASAP7_75t_L g2794 ( 
.A1(n_2757),
.A2(n_2735),
.B(n_2712),
.Y(n_2794)
);

CKINVDCx16_ASAP7_75t_R g2795 ( 
.A(n_2774),
.Y(n_2795)
);

CKINVDCx16_ASAP7_75t_R g2796 ( 
.A(n_2774),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2771),
.B(n_2683),
.Y(n_2797)
);

NAND2xp33_ASAP7_75t_R g2798 ( 
.A(n_2776),
.B(n_2704),
.Y(n_2798)
);

NOR2x1_ASAP7_75t_L g2799 ( 
.A(n_2758),
.B(n_2699),
.Y(n_2799)
);

INVx2_ASAP7_75t_SL g2800 ( 
.A(n_2752),
.Y(n_2800)
);

NOR2x1_ASAP7_75t_L g2801 ( 
.A(n_2763),
.B(n_2715),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2744),
.Y(n_2802)
);

AND3x4_ASAP7_75t_L g2803 ( 
.A(n_2787),
.B(n_2718),
.C(n_2724),
.Y(n_2803)
);

CKINVDCx5p33_ASAP7_75t_R g2804 ( 
.A(n_2767),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2780),
.Y(n_2805)
);

BUFx2_ASAP7_75t_L g2806 ( 
.A(n_2773),
.Y(n_2806)
);

BUFx2_ASAP7_75t_L g2807 ( 
.A(n_2773),
.Y(n_2807)
);

CKINVDCx16_ASAP7_75t_R g2808 ( 
.A(n_2766),
.Y(n_2808)
);

HB1xp67_ASAP7_75t_L g2809 ( 
.A(n_2777),
.Y(n_2809)
);

INVx1_ASAP7_75t_SL g2810 ( 
.A(n_2748),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2746),
.Y(n_2811)
);

AOI221xp5_ASAP7_75t_L g2812 ( 
.A1(n_2782),
.A2(n_2695),
.B1(n_2709),
.B2(n_2688),
.C(n_477),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2765),
.Y(n_2813)
);

BUFx2_ASAP7_75t_L g2814 ( 
.A(n_2753),
.Y(n_2814)
);

CKINVDCx16_ASAP7_75t_R g2815 ( 
.A(n_2747),
.Y(n_2815)
);

CKINVDCx5p33_ASAP7_75t_R g2816 ( 
.A(n_2768),
.Y(n_2816)
);

OAI221xp5_ASAP7_75t_L g2817 ( 
.A1(n_2745),
.A2(n_474),
.B1(n_475),
.B2(n_476),
.C(n_477),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2755),
.Y(n_2818)
);

BUFx2_ASAP7_75t_L g2819 ( 
.A(n_2760),
.Y(n_2819)
);

CKINVDCx5p33_ASAP7_75t_R g2820 ( 
.A(n_2779),
.Y(n_2820)
);

OAI211xp5_ASAP7_75t_L g2821 ( 
.A1(n_2749),
.A2(n_475),
.B(n_476),
.C(n_478),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_2764),
.Y(n_2822)
);

AOI322xp5_ASAP7_75t_L g2823 ( 
.A1(n_2801),
.A2(n_2786),
.A3(n_2785),
.B1(n_2756),
.B2(n_2784),
.C1(n_2751),
.C2(n_2769),
.Y(n_2823)
);

AOI322xp5_ASAP7_75t_L g2824 ( 
.A1(n_2800),
.A2(n_2759),
.A3(n_2761),
.B1(n_2754),
.B2(n_2778),
.C1(n_2750),
.C2(n_2762),
.Y(n_2824)
);

INVx6_ASAP7_75t_L g2825 ( 
.A(n_2795),
.Y(n_2825)
);

NOR3xp33_ASAP7_75t_L g2826 ( 
.A(n_2815),
.B(n_478),
.C(n_479),
.Y(n_2826)
);

AND2x4_ASAP7_75t_L g2827 ( 
.A(n_2799),
.B(n_480),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2806),
.Y(n_2828)
);

NOR3xp33_ASAP7_75t_L g2829 ( 
.A(n_2796),
.B(n_481),
.C(n_482),
.Y(n_2829)
);

OAI211xp5_ASAP7_75t_SL g2830 ( 
.A1(n_2794),
.A2(n_481),
.B(n_482),
.C(n_483),
.Y(n_2830)
);

AOI322xp5_ASAP7_75t_L g2831 ( 
.A1(n_2810),
.A2(n_484),
.A3(n_485),
.B1(n_486),
.B2(n_487),
.C1(n_488),
.C2(n_489),
.Y(n_2831)
);

NAND3xp33_ASAP7_75t_SL g2832 ( 
.A(n_2820),
.B(n_2788),
.C(n_2816),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2807),
.Y(n_2833)
);

BUFx2_ASAP7_75t_L g2834 ( 
.A(n_2791),
.Y(n_2834)
);

OAI322xp33_ASAP7_75t_L g2835 ( 
.A1(n_2813),
.A2(n_484),
.A3(n_485),
.B1(n_486),
.B2(n_487),
.C1(n_488),
.C2(n_490),
.Y(n_2835)
);

NAND3xp33_ASAP7_75t_SL g2836 ( 
.A(n_2790),
.B(n_490),
.C(n_491),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2804),
.A2(n_492),
.B1(n_493),
.B2(n_494),
.Y(n_2837)
);

AOI322xp5_ASAP7_75t_L g2838 ( 
.A1(n_2812),
.A2(n_492),
.A3(n_494),
.B1(n_495),
.B2(n_496),
.C1(n_497),
.C2(n_498),
.Y(n_2838)
);

NOR2xp67_ASAP7_75t_L g2839 ( 
.A(n_2821),
.B(n_495),
.Y(n_2839)
);

OAI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_2817),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_2840)
);

OAI211xp5_ASAP7_75t_SL g2841 ( 
.A1(n_2818),
.A2(n_499),
.B(n_500),
.C(n_501),
.Y(n_2841)
);

AOI322xp5_ASAP7_75t_L g2842 ( 
.A1(n_2797),
.A2(n_499),
.A3(n_500),
.B1(n_501),
.B2(n_502),
.C1(n_503),
.C2(n_504),
.Y(n_2842)
);

NOR2x1_ASAP7_75t_L g2843 ( 
.A(n_2793),
.B(n_502),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2797),
.Y(n_2844)
);

OAI211xp5_ASAP7_75t_L g2845 ( 
.A1(n_2809),
.A2(n_2814),
.B(n_2819),
.C(n_2805),
.Y(n_2845)
);

AOI221xp5_ASAP7_75t_L g2846 ( 
.A1(n_2789),
.A2(n_503),
.B1(n_504),
.B2(n_505),
.C(n_506),
.Y(n_2846)
);

OAI221xp5_ASAP7_75t_L g2847 ( 
.A1(n_2792),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.C(n_508),
.Y(n_2847)
);

AOI322xp5_ASAP7_75t_L g2848 ( 
.A1(n_2808),
.A2(n_507),
.A3(n_508),
.B1(n_509),
.B2(n_510),
.C1(n_511),
.C2(n_512),
.Y(n_2848)
);

AOI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2825),
.A2(n_2803),
.B1(n_2798),
.B2(n_2822),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2843),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2827),
.Y(n_2851)
);

OAI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2825),
.A2(n_2802),
.B1(n_2811),
.B2(n_511),
.Y(n_2852)
);

OAI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2833),
.A2(n_509),
.B1(n_510),
.B2(n_512),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2834),
.Y(n_2854)
);

OAI22x1_ASAP7_75t_L g2855 ( 
.A1(n_2828),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.Y(n_2855)
);

AO22x2_ASAP7_75t_L g2856 ( 
.A1(n_2844),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.Y(n_2856)
);

OAI22xp5_ASAP7_75t_SL g2857 ( 
.A1(n_2840),
.A2(n_516),
.B1(n_517),
.B2(n_518),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2832),
.A2(n_517),
.B1(n_519),
.B2(n_520),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2836),
.A2(n_520),
.B1(n_521),
.B2(n_522),
.Y(n_2859)
);

AOI22x1_ASAP7_75t_L g2860 ( 
.A1(n_2845),
.A2(n_522),
.B1(n_523),
.B2(n_524),
.Y(n_2860)
);

INVxp67_ASAP7_75t_L g2861 ( 
.A(n_2839),
.Y(n_2861)
);

OAI22xp5_ASAP7_75t_SL g2862 ( 
.A1(n_2847),
.A2(n_524),
.B1(n_525),
.B2(n_526),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2830),
.Y(n_2863)
);

OR3x1_ASAP7_75t_L g2864 ( 
.A(n_2854),
.B(n_2841),
.C(n_2823),
.Y(n_2864)
);

AOI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2862),
.A2(n_2826),
.B1(n_2829),
.B2(n_2846),
.Y(n_2865)
);

NAND4xp25_ASAP7_75t_L g2866 ( 
.A(n_2849),
.B(n_2824),
.C(n_2838),
.D(n_2837),
.Y(n_2866)
);

OAI221xp5_ASAP7_75t_L g2867 ( 
.A1(n_2859),
.A2(n_2831),
.B1(n_2842),
.B2(n_2848),
.C(n_2835),
.Y(n_2867)
);

NAND5xp2_ASAP7_75t_L g2868 ( 
.A(n_2863),
.B(n_525),
.C(n_526),
.D(n_527),
.E(n_528),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2852),
.Y(n_2869)
);

AOI221xp5_ASAP7_75t_L g2870 ( 
.A1(n_2861),
.A2(n_527),
.B1(n_528),
.B2(n_529),
.C(n_530),
.Y(n_2870)
);

OAI221xp5_ASAP7_75t_L g2871 ( 
.A1(n_2860),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.C(n_532),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2856),
.Y(n_2872)
);

OAI22xp5_ASAP7_75t_L g2873 ( 
.A1(n_2858),
.A2(n_532),
.B1(n_533),
.B2(n_534),
.Y(n_2873)
);

HB1xp67_ASAP7_75t_L g2874 ( 
.A(n_2872),
.Y(n_2874)
);

AOI221xp5_ASAP7_75t_L g2875 ( 
.A1(n_2867),
.A2(n_2850),
.B1(n_2857),
.B2(n_2851),
.C(n_2855),
.Y(n_2875)
);

OAI31xp33_ASAP7_75t_L g2876 ( 
.A1(n_2871),
.A2(n_2853),
.A3(n_2856),
.B(n_535),
.Y(n_2876)
);

OA21x2_ASAP7_75t_L g2877 ( 
.A1(n_2866),
.A2(n_533),
.B(n_534),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2873),
.B(n_536),
.Y(n_2878)
);

OAI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2865),
.A2(n_536),
.B(n_537),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2870),
.B(n_537),
.Y(n_2880)
);

AOI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_2869),
.A2(n_538),
.B(n_539),
.Y(n_2881)
);

OAI22x1_ASAP7_75t_L g2882 ( 
.A1(n_2874),
.A2(n_2864),
.B1(n_2868),
.B2(n_541),
.Y(n_2882)
);

AOI21xp5_ASAP7_75t_L g2883 ( 
.A1(n_2875),
.A2(n_539),
.B(n_540),
.Y(n_2883)
);

OAI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2878),
.A2(n_2880),
.B(n_2876),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2877),
.Y(n_2885)
);

AOI222xp33_ASAP7_75t_L g2886 ( 
.A1(n_2879),
.A2(n_540),
.B1(n_542),
.B2(n_543),
.C1(n_544),
.C2(n_545),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2881),
.Y(n_2887)
);

AOI211x1_ASAP7_75t_SL g2888 ( 
.A1(n_2880),
.A2(n_544),
.B(n_545),
.C(n_546),
.Y(n_2888)
);

OAI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2883),
.A2(n_546),
.B(n_547),
.Y(n_2889)
);

OAI21xp5_ASAP7_75t_SL g2890 ( 
.A1(n_2888),
.A2(n_548),
.B(n_549),
.Y(n_2890)
);

OAI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2884),
.A2(n_548),
.B(n_550),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2890),
.A2(n_2885),
.B(n_2887),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2889),
.A2(n_2882),
.B1(n_2886),
.B2(n_553),
.Y(n_2893)
);

AOI22xp33_ASAP7_75t_L g2894 ( 
.A1(n_2891),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2891),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_L g2896 ( 
.A1(n_2894),
.A2(n_551),
.B1(n_554),
.B2(n_555),
.Y(n_2896)
);

AO22x2_ASAP7_75t_L g2897 ( 
.A1(n_2893),
.A2(n_554),
.B1(n_557),
.B2(n_558),
.Y(n_2897)
);

OR2x6_ASAP7_75t_L g2898 ( 
.A(n_2896),
.B(n_2892),
.Y(n_2898)
);

OR2x2_ASAP7_75t_L g2899 ( 
.A(n_2897),
.B(n_2895),
.Y(n_2899)
);

CKINVDCx20_ASAP7_75t_R g2900 ( 
.A(n_2899),
.Y(n_2900)
);

AOI22xp5_ASAP7_75t_L g2901 ( 
.A1(n_2900),
.A2(n_2898),
.B1(n_559),
.B2(n_560),
.Y(n_2901)
);

XNOR2xp5_ASAP7_75t_L g2902 ( 
.A(n_2901),
.B(n_557),
.Y(n_2902)
);

AOI211xp5_ASAP7_75t_L g2903 ( 
.A1(n_2902),
.A2(n_559),
.B(n_560),
.C(n_561),
.Y(n_2903)
);


endmodule