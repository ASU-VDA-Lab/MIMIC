module fake_jpeg_22434_n_31 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_13),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_16),
.A2(n_8),
.B1(n_13),
.B2(n_9),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_10),
.C(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_18),
.B(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_19),
.C(n_18),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_24),
.C(n_8),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_12),
.C(n_17),
.Y(n_24)
);

AOI21x1_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B(n_12),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_12),
.B1(n_14),
.B2(n_2),
.Y(n_26)
);

OAI21x1_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_12),
.B(n_1),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_0),
.C(n_4),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_5),
.C(n_6),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_6),
.Y(n_31)
);


endmodule