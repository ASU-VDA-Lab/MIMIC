module real_jpeg_12664_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_3),
.A2(n_33),
.B1(n_55),
.B2(n_56),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_4),
.A2(n_36),
.B1(n_43),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_48),
.B1(n_55),
.B2(n_56),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_48),
.Y(n_193)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_55),
.B1(n_56),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_84),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_6),
.A2(n_36),
.B1(n_43),
.B2(n_84),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_7),
.A2(n_36),
.B1(n_43),
.B2(n_67),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_67),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_36),
.B1(n_43),
.B2(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_55),
.B1(n_56),
.B2(n_69),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_69),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_11),
.B(n_90),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_11),
.B(n_26),
.C(n_79),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_11),
.A2(n_41),
.B1(n_55),
.B2(n_56),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_93),
.B1(n_97),
.B2(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_11),
.B(n_58),
.Y(n_210)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_13),
.A2(n_36),
.B1(n_43),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_13),
.A2(n_55),
.B1(n_56),
.B2(n_60),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_60),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_14),
.A2(n_31),
.B1(n_55),
.B2(n_56),
.Y(n_101)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_104),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.C(n_91),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_20),
.B(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_45),
.B1(n_70),
.B2(n_71),
.Y(n_20)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_22),
.A2(n_23),
.B1(n_34),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_23)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_24),
.B(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_24),
.A2(n_96),
.B(n_123),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_24),
.A2(n_28),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_25),
.A2(n_26),
.B1(n_77),
.B2(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_25),
.B(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_28),
.B(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_30),
.A2(n_97),
.B(n_120),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_34),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B(n_37),
.C(n_42),
.Y(n_34)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_44),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_64)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_43),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g158 ( 
.A(n_36),
.B(n_41),
.CON(n_158),
.SN(n_158)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_36),
.B(n_53),
.C(n_56),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_37),
.A2(n_66),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.CON(n_37),
.SN(n_37)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_43),
.C(n_44),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_41),
.B(n_97),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_41),
.B(n_100),
.Y(n_201)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_61),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_61),
.C(n_70),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_49),
.B1(n_54),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_49),
.A2(n_54),
.B1(n_87),
.B2(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_50),
.A2(n_59),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_50),
.A2(n_58),
.B1(n_142),
.B2(n_158),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_52),
.A2(n_55),
.B(n_158),
.C(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_56),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_55),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_64),
.B1(n_68),
.B2(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_91),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_85),
.C(n_88),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_73),
.A2(n_74),
.B1(n_85),
.B2(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_81),
.B(n_82),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_75),
.A2(n_100),
.B1(n_101),
.B2(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_75),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_75),
.A2(n_100),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_75),
.A2(n_100),
.B1(n_163),
.B2(n_188),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_SL g79 ( 
.A(n_77),
.Y(n_79)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_80),
.B(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_80),
.A2(n_103),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_80),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_99),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B(n_95),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_93),
.A2(n_97),
.B1(n_191),
.B2(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_93),
.A2(n_122),
.B(n_193),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_124),
.B2(n_125),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_228),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_148),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_146),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_133),
.B(n_146),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_139),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_134),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_145),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_222),
.B(n_227),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_177),
.B(n_221),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_165),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_151),
.B(n_165),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_160),
.C(n_161),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_152),
.A2(n_153),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_161),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_164),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_171),
.C(n_175),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_169)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_215),
.B(n_220),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_205),
.B(n_214),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_194),
.B(n_204),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_189),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_200),
.B(n_203),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_207),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_219)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_219),
.Y(n_220)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_226),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);


endmodule