module real_jpeg_5255_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_0),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_0),
.Y(n_211)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_0),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_0),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

INVx8_ASAP7_75t_L g414 ( 
.A(n_0),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_1),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_1),
.A2(n_148),
.B1(n_196),
.B2(n_265),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_1),
.A2(n_68),
.B1(n_265),
.B2(n_386),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_L g442 ( 
.A1(n_1),
.A2(n_265),
.B1(n_322),
.B2(n_443),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_2),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_2),
.Y(n_331)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_2),
.Y(n_346)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_2),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_2),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_3),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_3),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_87),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_3),
.A2(n_87),
.B1(n_115),
.B2(n_176),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_3),
.A2(n_87),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_4),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_5),
.A2(n_52),
.B1(n_300),
.B2(n_303),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_5),
.A2(n_52),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_5),
.A2(n_52),
.B1(n_269),
.B2(n_388),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_148),
.B1(n_150),
.B2(n_152),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_6),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_6),
.B(n_112),
.C(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_6),
.B(n_73),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_6),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_6),
.B(n_157),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_6),
.B(n_92),
.Y(n_253)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_7),
.Y(n_520)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_10),
.A2(n_95),
.B1(n_101),
.B2(n_123),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_10),
.A2(n_95),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_10),
.A2(n_95),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_11),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_11),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_11),
.A2(n_197),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_11),
.A2(n_92),
.B1(n_197),
.B2(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_11),
.A2(n_48),
.B1(n_197),
.B2(n_350),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_12),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_13),
.A2(n_101),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_13),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_13),
.A2(n_156),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_13),
.A2(n_156),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_13),
.A2(n_156),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_15),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_15),
.A2(n_175),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_15),
.A2(n_175),
.B1(n_291),
.B2(n_356),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_15),
.A2(n_51),
.B1(n_175),
.B2(n_394),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_16),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_17),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_17),
.A2(n_60),
.B1(n_163),
.B2(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_17),
.A2(n_60),
.B1(n_123),
.B2(n_380),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_17),
.A2(n_60),
.B1(n_270),
.B2(n_429),
.Y(n_428)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_518),
.B(n_521),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_137),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_135),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_131),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_23),
.B(n_131),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_124),
.C(n_128),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_24),
.A2(n_25),
.B1(n_514),
.B2(n_515),
.Y(n_513)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_61),
.C(n_96),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_26),
.B(n_506),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_27),
.A2(n_53),
.B1(n_55),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_27),
.A2(n_53),
.B1(n_125),
.B2(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_27),
.A2(n_348),
.B(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_27),
.A2(n_37),
.B1(n_393),
.B2(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_27),
.A2(n_47),
.B1(n_53),
.B2(n_491),
.Y(n_490)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_28),
.A2(n_344),
.B(n_347),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_28),
.B(n_349),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_35),
.Y(n_352)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_37),
.B(n_152),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_38),
.A2(n_316),
.A3(n_319),
.B1(n_323),
.B2(n_328),
.Y(n_315)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_41),
.Y(n_271)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_42),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_42),
.Y(n_259)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_45),
.Y(n_386)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_53),
.A2(n_417),
.B(n_445),
.Y(n_455)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_54),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_54),
.B(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_61),
.A2(n_96),
.B1(n_97),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_61),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_62),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_62),
.A2(n_88),
.B1(n_290),
.B2(n_355),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_62),
.A2(n_88),
.B1(n_385),
.B2(n_387),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_62),
.A2(n_81),
.B1(n_88),
.B2(n_495),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_73),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_63)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_64),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_67),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_72),
.Y(n_251)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_72),
.Y(n_318)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_72),
.Y(n_327)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_72),
.Y(n_391)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_72),
.Y(n_430)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

AOI22x1_ASAP7_75t_L g418 ( 
.A1(n_73),
.A2(n_129),
.B1(n_295),
.B2(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_73),
.A2(n_129),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_73)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_75),
.Y(n_273)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_76),
.Y(n_382)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_77),
.Y(n_199)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_77),
.Y(n_378)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_88),
.B(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_88),
.A2(n_290),
.B(n_294),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_93),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_96),
.A2(n_97),
.B1(n_493),
.B2(n_494),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_96),
.B(n_490),
.C(n_493),
.Y(n_501)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_111),
.B(n_122),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_147),
.B(n_153),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_98),
.A2(n_194),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_98),
.A2(n_153),
.B(n_244),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_98),
.A2(n_243),
.B1(n_360),
.B2(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_99),
.B(n_154),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_99),
.A2(n_157),
.B1(n_374),
.B2(n_379),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_99),
.A2(n_157),
.B1(n_379),
.B2(n_399),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_99),
.A2(n_157),
.B1(n_399),
.B2(n_433),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_111),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_106),
.B2(n_108),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx5_ASAP7_75t_SL g247 ( 
.A(n_108),
.Y(n_247)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_111),
.A2(n_194),
.B(n_200),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_111),
.A2(n_200),
.B(n_360),
.Y(n_359)
);

AOI22x1_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_122),
.Y(n_433)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_123),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_124),
.B(n_128),
.Y(n_515)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_129),
.A2(n_250),
.B(n_254),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_129),
.B(n_295),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_129),
.A2(n_254),
.B(n_458),
.Y(n_457)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_512),
.B(n_517),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_484),
.B(n_509),
.Y(n_138)
);

OAI311xp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_363),
.A3(n_460),
.B1(n_478),
.C1(n_483),
.Y(n_139)
);

AOI21x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_309),
.B(n_362),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_281),
.B(n_308),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_237),
.B(n_280),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_203),
.B(n_236),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_168),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_145),
.B(n_168),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_158),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_146),
.A2(n_158),
.B1(n_159),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_150),
.B(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_150),
.Y(n_401)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g400 ( 
.A(n_151),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_152),
.A2(n_178),
.B(n_183),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_SL g250 ( 
.A1(n_152),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_152),
.B(n_329),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_SL g344 ( 
.A1(n_152),
.A2(n_328),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_191),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_169),
.B(n_192),
.C(n_202),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_178),
.B(n_183),
.Y(n_169)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_173),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

BUFx8_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_178),
.A2(n_209),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_178),
.A2(n_232),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_178),
.A2(n_370),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_185),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_179),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_179),
.A2(n_263),
.B1(n_299),
.B2(n_305),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_179),
.A2(n_336),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_181),
.Y(n_266)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_188),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_189),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_201),
.B2(n_202),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_227),
.B(n_235),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_213),
.B(n_226),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_225),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_225),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_222),
.B(n_224),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_216),
.Y(n_372)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_262),
.B(n_267),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_233),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_239),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_260),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_248),
.B2(n_249),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_248),
.C(n_260),
.Y(n_282)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI32xp33_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_269),
.A3(n_272),
.B1(n_274),
.B2(n_278),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_273),
.Y(n_375)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_282),
.B(n_283),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_288),
.B2(n_307),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_287),
.C(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_296),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_297),
.C(n_298),
.Y(n_338)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_305),
.Y(n_403)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_310),
.B(n_311),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_341),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_312)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_332),
.B2(n_333),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_315),
.B(n_332),
.Y(n_456)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_338),
.B(n_339),
.C(n_341),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_353),
.B2(n_361),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_342),
.B(n_354),
.C(n_359),
.Y(n_469)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_353),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_359),
.Y(n_353)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_355),
.Y(n_458)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_SL g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_446),
.Y(n_363)
);

A2O1A1Ixp33_ASAP7_75t_SL g478 ( 
.A1(n_364),
.A2(n_446),
.B(n_479),
.C(n_482),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_420),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_365),
.B(n_420),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_396),
.C(n_405),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g459 ( 
.A(n_366),
.B(n_396),
.CI(n_405),
.CON(n_459),
.SN(n_459)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_383),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_384),
.C(n_392),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_373),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_368),
.B(n_373),
.Y(n_452)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx6_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_392),
.Y(n_383)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

INVx5_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_402),
.B2(n_404),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_402),
.Y(n_437)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_402),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_402),
.A2(n_404),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_402),
.A2(n_437),
.B(n_440),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_415),
.C(n_418),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_407),
.B(n_409),
.Y(n_468)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx8_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_415),
.A2(n_416),
.B1(n_418),
.B2(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_418),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_421),
.B(n_424),
.C(n_435),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_435),
.B2(n_436),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_431),
.B(n_434),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_432),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_428),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g486 ( 
.A(n_434),
.B(n_487),
.CI(n_488),
.CON(n_486),
.SN(n_486)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_434),
.B(n_487),
.C(n_488),
.Y(n_508)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_445),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_442),
.Y(n_491)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_459),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_459),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_452),
.C(n_453),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_448),
.A2(n_449),
.B1(n_452),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_452),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.C(n_457),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_454),
.A2(n_455),
.B1(n_457),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_459),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_473),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_462),
.A2(n_480),
.B(n_481),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_470),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_470),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_467),
.C(n_469),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_476),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_467),
.A2(n_468),
.B1(n_469),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_469),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_474),
.B(n_475),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_498),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_486),
.B(n_497),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_497),
.Y(n_510)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_486),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_489),
.A2(n_490),
.B1(n_492),
.B2(n_496),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_489),
.A2(n_490),
.B1(n_504),
.B2(n_505),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_489),
.B(n_500),
.C(n_504),
.Y(n_516)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_492),
.Y(n_496)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_498),
.A2(n_510),
.B(n_511),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_508),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_508),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_513),
.B(n_516),
.Y(n_517)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx13_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_520),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_524),
.Y(n_521)
);

BUFx12f_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);


endmodule