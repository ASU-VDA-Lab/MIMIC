module fake_jpeg_20098_n_106 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_4),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_27),
.B(n_20),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_4),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_12),
.B1(n_15),
.B2(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_13),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_35),
.B(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_12),
.B1(n_21),
.B2(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_41),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_25),
.Y(n_39)
);

OAI21x1_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_43),
.B(n_45),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_34),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_18),
.B1(n_15),
.B2(n_25),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_17),
.B1(n_32),
.B2(n_14),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_26),
.B1(n_24),
.B2(n_20),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_34),
.B1(n_32),
.B2(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_51),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_53),
.B1(n_56),
.B2(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_36),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_45),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_17),
.B1(n_11),
.B2(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_71),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_39),
.B(n_37),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_65),
.B(n_68),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_39),
.C(n_37),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_60),
.B1(n_56),
.B2(n_55),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_R g67 ( 
.A(n_57),
.B(n_39),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_45),
.C(n_42),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_50),
.B1(n_60),
.B2(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_79),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_58),
.B(n_53),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_64),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_78),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_63),
.C(n_70),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_11),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_61),
.C(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_92),
.B1(n_11),
.B2(n_19),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_87),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_83),
.B1(n_82),
.B2(n_11),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_2),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_6),
.C1(n_7),
.C2(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_3),
.Y(n_99)
);

NOR2xp67_ASAP7_75t_SL g97 ( 
.A(n_94),
.B(n_1),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_94),
.B(n_93),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_6),
.C(n_7),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_0),
.A3(n_3),
.B1(n_6),
.B2(n_7),
.C1(n_100),
.C2(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_105),
.Y(n_106)
);


endmodule