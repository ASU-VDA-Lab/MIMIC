module fake_jpeg_18086_n_167 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_9),
.B(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_38),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_18),
.B1(n_26),
.B2(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_15),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_17),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_37),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_30),
.B1(n_24),
.B2(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_22),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_48),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_26),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_61),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_26),
.B1(n_22),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_52),
.B1(n_67),
.B2(n_20),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_27),
.B1(n_25),
.B2(n_16),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_54),
.A2(n_45),
.B1(n_47),
.B2(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_25),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_30),
.C(n_16),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_16),
.C(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_68),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_93),
.B1(n_62),
.B2(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_77),
.B(n_92),
.Y(n_112)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_6),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_45),
.B1(n_32),
.B2(n_21),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_32),
.B(n_37),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_91),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_3),
.B(n_5),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_13),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_51),
.B1(n_61),
.B2(n_46),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_13),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_98),
.B1(n_99),
.B2(n_108),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_74),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_50),
.B1(n_62),
.B2(n_55),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_7),
.C(n_11),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_106),
.C(n_110),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_7),
.C(n_3),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_6),
.B1(n_88),
.B2(n_83),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_71),
.CI(n_86),
.CON(n_122),
.SN(n_122)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_69),
.Y(n_110)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_91),
.B(n_75),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_82),
.B(n_79),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_119),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_118),
.C(n_108),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_124),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_122),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_97),
.B(n_89),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_103),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_111),
.B(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_132),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_122),
.B1(n_119),
.B2(n_90),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_99),
.B1(n_125),
.B2(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_136),
.B(n_137),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_106),
.C(n_105),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_138),
.B(n_120),
.C(n_113),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_118),
.C(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_140),
.B(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_70),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_113),
.C(n_98),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_132),
.B(n_129),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_140),
.Y(n_157)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_135),
.A3(n_81),
.B1(n_94),
.B2(n_102),
.C(n_127),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_147),
.C(n_146),
.Y(n_156)
);

AOI31xp33_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_159),
.A3(n_117),
.B(n_78),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

OAI211xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_152),
.B(n_153),
.C(n_101),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_76),
.C(n_73),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_76),
.C(n_72),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_166),
.CI(n_158),
.CON(n_167),
.SN(n_167)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_72),
.C(n_153),
.Y(n_166)
);


endmodule