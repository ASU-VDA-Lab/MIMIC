module real_aes_491_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_789, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_789;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g172 ( .A(n_0), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_1), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_2), .B(n_178), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_3), .B(n_175), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_4), .A2(n_43), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_4), .Y(n_448) );
INVx1_ASAP7_75t_L g138 ( .A(n_5), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_6), .B(n_178), .Y(n_200) );
NAND2xp33_ASAP7_75t_SL g158 ( .A(n_7), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g129 ( .A(n_8), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_9), .Y(n_114) );
AND2x2_ASAP7_75t_L g198 ( .A(n_10), .B(n_181), .Y(n_198) );
AND2x2_ASAP7_75t_L g504 ( .A(n_11), .B(n_154), .Y(n_504) );
AND2x2_ASAP7_75t_L g555 ( .A(n_12), .B(n_209), .Y(n_555) );
INVx2_ASAP7_75t_L g132 ( .A(n_13), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_14), .B(n_175), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_15), .Y(n_115) );
AOI221x1_ASAP7_75t_L g150 ( .A1(n_16), .A2(n_151), .B1(n_153), .B2(n_154), .C(n_157), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_17), .B(n_178), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_18), .B(n_178), .Y(n_560) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_19), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g461 ( .A(n_19), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_20), .A2(n_92), .B1(n_133), .B2(n_178), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_21), .A2(n_153), .B(n_202), .Y(n_201) );
AOI221xp5_ASAP7_75t_SL g245 ( .A1(n_22), .A2(n_35), .B1(n_153), .B2(n_178), .C(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_23), .B(n_173), .Y(n_203) );
OR2x2_ASAP7_75t_L g131 ( .A(n_24), .B(n_91), .Y(n_131) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_24), .A2(n_91), .B(n_132), .Y(n_156) );
INVxp67_ASAP7_75t_L g149 ( .A(n_25), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_26), .B(n_175), .Y(n_240) );
AND2x2_ASAP7_75t_L g192 ( .A(n_27), .B(n_180), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_28), .A2(n_153), .B(n_171), .Y(n_170) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_29), .A2(n_154), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_30), .B(n_175), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_31), .A2(n_153), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_32), .B(n_175), .Y(n_536) );
AND2x2_ASAP7_75t_L g140 ( .A(n_33), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g144 ( .A(n_33), .Y(n_144) );
AND2x2_ASAP7_75t_L g159 ( .A(n_33), .B(n_138), .Y(n_159) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_34), .B(n_113), .C(n_115), .Y(n_112) );
OR2x6_ASAP7_75t_L g459 ( .A(n_34), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_36), .B(n_178), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_37), .A2(n_84), .B1(n_142), .B2(n_153), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_38), .B(n_175), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_39), .A2(n_48), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_39), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_40), .B(n_178), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_41), .B(n_173), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_42), .A2(n_153), .B(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_43), .Y(n_449) );
AND2x2_ASAP7_75t_L g179 ( .A(n_44), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_45), .B(n_173), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_46), .B(n_180), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_47), .B(n_178), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_48), .Y(n_780) );
INVx1_ASAP7_75t_L g136 ( .A(n_49), .Y(n_136) );
INVx1_ASAP7_75t_L g163 ( .A(n_49), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_50), .B(n_175), .Y(n_502) );
AND2x2_ASAP7_75t_L g514 ( .A(n_51), .B(n_180), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_52), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_53), .B(n_178), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_54), .B(n_173), .Y(n_501) );
INVxp33_ASAP7_75t_L g786 ( .A(n_55), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_56), .B(n_173), .Y(n_535) );
AND2x2_ASAP7_75t_L g221 ( .A(n_57), .B(n_180), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_58), .B(n_178), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_59), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_60), .B(n_178), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_61), .A2(n_153), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_62), .B(n_173), .Y(n_219) );
AND2x2_ASAP7_75t_SL g241 ( .A(n_63), .B(n_181), .Y(n_241) );
XNOR2xp5_ASAP7_75t_L g778 ( .A(n_64), .B(n_779), .Y(n_778) );
XNOR2x1_ASAP7_75t_SL g118 ( .A(n_65), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g566 ( .A(n_65), .B(n_181), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_66), .A2(n_153), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_67), .B(n_175), .Y(n_204) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_68), .B(n_209), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_69), .B(n_173), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_70), .B(n_173), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_71), .A2(n_94), .B1(n_142), .B2(n_153), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_72), .B(n_467), .Y(n_466) );
XNOR2xp5_ASAP7_75t_L g777 ( .A(n_73), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_74), .B(n_175), .Y(n_563) );
INVx1_ASAP7_75t_L g141 ( .A(n_75), .Y(n_141) );
INVx1_ASAP7_75t_L g165 ( .A(n_75), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_76), .B(n_173), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_77), .A2(n_153), .B(n_518), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_78), .A2(n_153), .B(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_79), .A2(n_153), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g538 ( .A(n_80), .B(n_181), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_81), .B(n_180), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_82), .A2(n_86), .B1(n_133), .B2(n_178), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_83), .B(n_178), .Y(n_220) );
INVx1_ASAP7_75t_L g111 ( .A(n_85), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_87), .B(n_173), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_88), .B(n_173), .Y(n_248) );
AND2x2_ASAP7_75t_L g495 ( .A(n_89), .B(n_209), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_90), .A2(n_153), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_93), .B(n_175), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_95), .A2(n_153), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_96), .B(n_175), .Y(n_493) );
OAI22x1_ASAP7_75t_R g445 ( .A1(n_97), .A2(n_446), .B1(n_447), .B2(n_450), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_97), .Y(n_450) );
INVxp67_ASAP7_75t_L g152 ( .A(n_98), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_99), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_100), .B(n_175), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_101), .A2(n_153), .B(n_238), .Y(n_237) );
BUFx2_ASAP7_75t_L g565 ( .A(n_102), .Y(n_565) );
BUFx2_ASAP7_75t_L g452 ( .A(n_103), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_116), .B(n_785), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g787 ( .A(n_108), .Y(n_787) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_112), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_111), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_115), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g470 ( .A(n_115), .B(n_459), .Y(n_470) );
AND2x6_ASAP7_75t_SL g478 ( .A(n_115), .B(n_459), .Y(n_478) );
OR2x6_ASAP7_75t_SL g482 ( .A(n_115), .B(n_458), .Y(n_482) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_463), .Y(n_116) );
AOI22x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_451), .B1(n_454), .B2(n_462), .Y(n_117) );
OAI22x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B1(n_444), .B2(n_445), .Y(n_119) );
OAI22x1_ASAP7_75t_L g783 ( .A1(n_120), .A2(n_477), .B1(n_480), .B2(n_784), .Y(n_783) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OA22x2_ASAP7_75t_L g476 ( .A1(n_121), .A2(n_477), .B1(n_479), .B2(n_483), .Y(n_476) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_321), .Y(n_121) );
NOR4xp25_ASAP7_75t_L g122 ( .A(n_123), .B(n_264), .C(n_303), .D(n_310), .Y(n_122) );
OAI221xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_182), .B1(n_222), .B2(n_231), .C(n_250), .Y(n_123) );
OR2x2_ASAP7_75t_L g394 ( .A(n_124), .B(n_256), .Y(n_394) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g309 ( .A(n_125), .B(n_234), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_125), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_125), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_166), .Y(n_125) );
AND2x4_ASAP7_75t_SL g233 ( .A(n_126), .B(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g255 ( .A(n_126), .Y(n_255) );
AND2x2_ASAP7_75t_L g290 ( .A(n_126), .B(n_263), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_126), .B(n_167), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_126), .B(n_257), .Y(n_342) );
OR2x2_ASAP7_75t_L g420 ( .A(n_126), .B(n_234), .Y(n_420) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_150), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_133), .B1(n_142), .B2(n_148), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_130), .B(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_130), .B(n_152), .Y(n_151) );
NOR3xp33_ASAP7_75t_L g157 ( .A(n_130), .B(n_158), .C(n_160), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_130), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_130), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_130), .A2(n_525), .B(n_526), .Y(n_524) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_131), .B(n_132), .Y(n_181) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_139), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g147 ( .A(n_136), .B(n_138), .Y(n_147) );
AND2x4_ASAP7_75t_L g175 ( .A(n_136), .B(n_164), .Y(n_175) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x6_ASAP7_75t_L g153 ( .A(n_140), .B(n_147), .Y(n_153) );
INVx2_ASAP7_75t_L g146 ( .A(n_141), .Y(n_146) );
AND2x6_ASAP7_75t_L g173 ( .A(n_141), .B(n_162), .Y(n_173) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_147), .Y(n_142) );
NOR2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g531 ( .A(n_154), .Y(n_531) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21x1_ASAP7_75t_L g168 ( .A1(n_155), .A2(n_169), .B(n_179), .Y(n_168) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_155), .A2(n_498), .B(n_504), .Y(n_497) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx4f_ASAP7_75t_L g209 ( .A(n_156), .Y(n_209) );
INVx5_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
AND2x4_ASAP7_75t_L g178 ( .A(n_159), .B(n_161), .Y(n_178) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g242 ( .A(n_167), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_167), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g268 ( .A(n_167), .Y(n_268) );
OR2x2_ASAP7_75t_L g273 ( .A(n_167), .B(n_257), .Y(n_273) );
AND2x2_ASAP7_75t_L g286 ( .A(n_167), .B(n_244), .Y(n_286) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_167), .Y(n_289) );
INVx1_ASAP7_75t_L g301 ( .A(n_167), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_167), .B(n_255), .Y(n_366) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_177), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .B(n_176), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_173), .B(n_565), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_176), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_176), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_176), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_176), .A2(n_239), .B(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_176), .A2(n_247), .B(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_176), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_176), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_176), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_176), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_176), .A2(n_535), .B(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_176), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_176), .A2(n_563), .B(n_564), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_180), .Y(n_191) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_180), .A2(n_245), .B(n_249), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_180), .A2(n_490), .B(n_491), .Y(n_489) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_180), .A2(n_508), .B(n_509), .Y(n_507) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_183), .B(n_193), .Y(n_182) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g230 ( .A(n_184), .B(n_214), .Y(n_230) );
AND2x4_ASAP7_75t_L g260 ( .A(n_184), .B(n_197), .Y(n_260) );
INVx2_ASAP7_75t_L g294 ( .A(n_184), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_184), .B(n_214), .Y(n_352) );
AND2x2_ASAP7_75t_L g399 ( .A(n_184), .B(n_228), .Y(n_399) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_191), .B(n_192), .Y(n_184) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_185), .A2(n_191), .B(n_192), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_190), .Y(n_185) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_191), .A2(n_215), .B(n_221), .Y(n_214) );
AOI21x1_ASAP7_75t_L g548 ( .A1(n_191), .A2(n_549), .B(n_555), .Y(n_548) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_193), .A2(n_259), .B1(n_302), .B2(n_362), .C1(n_388), .C2(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_205), .Y(n_194) );
AND2x2_ASAP7_75t_L g306 ( .A(n_195), .B(n_226), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_195), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g435 ( .A(n_195), .B(n_275), .Y(n_435) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_196), .A2(n_266), .B(n_270), .Y(n_265) );
AND2x2_ASAP7_75t_L g346 ( .A(n_196), .B(n_229), .Y(n_346) );
OR2x2_ASAP7_75t_L g371 ( .A(n_196), .B(n_230), .Y(n_371) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx5_ASAP7_75t_L g225 ( .A(n_197), .Y(n_225) );
AND2x2_ASAP7_75t_L g312 ( .A(n_197), .B(n_294), .Y(n_312) );
AND2x2_ASAP7_75t_L g338 ( .A(n_197), .B(n_214), .Y(n_338) );
OR2x2_ASAP7_75t_L g341 ( .A(n_197), .B(n_228), .Y(n_341) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_197), .Y(n_359) );
AND2x4_ASAP7_75t_SL g416 ( .A(n_197), .B(n_293), .Y(n_416) );
OR2x2_ASAP7_75t_L g425 ( .A(n_197), .B(n_252), .Y(n_425) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
AOI221xp5_ASAP7_75t_SL g376 ( .A1(n_205), .A2(n_260), .B1(n_377), .B2(n_379), .C(n_380), .Y(n_376) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_214), .Y(n_205) );
OR2x2_ASAP7_75t_L g315 ( .A(n_206), .B(n_285), .Y(n_315) );
OR2x2_ASAP7_75t_L g325 ( .A(n_206), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g351 ( .A(n_206), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g357 ( .A(n_206), .B(n_276), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_206), .B(n_340), .Y(n_369) );
INVx2_ASAP7_75t_L g382 ( .A(n_206), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_206), .B(n_260), .Y(n_403) );
AND2x2_ASAP7_75t_L g407 ( .A(n_206), .B(n_229), .Y(n_407) );
AND2x2_ASAP7_75t_L g415 ( .A(n_206), .B(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g228 ( .A(n_207), .Y(n_228) );
AOI21x1_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_210), .B(n_213), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_209), .A2(n_236), .B(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_209), .A2(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_214), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g259 ( .A(n_214), .B(n_228), .Y(n_259) );
INVx2_ASAP7_75t_L g276 ( .A(n_214), .Y(n_276) );
AND2x4_ASAP7_75t_L g293 ( .A(n_214), .B(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_214), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_220), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_226), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g405 ( .A(n_224), .B(n_227), .Y(n_405) );
AND2x4_ASAP7_75t_L g251 ( .A(n_225), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g292 ( .A(n_225), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g319 ( .A(n_225), .B(n_259), .Y(n_319) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
AND2x2_ASAP7_75t_L g423 ( .A(n_227), .B(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g275 ( .A(n_228), .B(n_276), .Y(n_275) );
OAI21xp5_ASAP7_75t_SL g295 ( .A1(n_229), .A2(n_296), .B(n_302), .Y(n_295) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_242), .Y(n_232) );
INVx1_ASAP7_75t_SL g349 ( .A(n_233), .Y(n_349) );
AND2x2_ASAP7_75t_L g379 ( .A(n_233), .B(n_289), .Y(n_379) );
AND2x4_ASAP7_75t_L g390 ( .A(n_233), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g256 ( .A(n_234), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g263 ( .A(n_234), .Y(n_263) );
AND2x4_ASAP7_75t_L g269 ( .A(n_234), .B(n_255), .Y(n_269) );
INVx2_ASAP7_75t_L g280 ( .A(n_234), .Y(n_280) );
INVx1_ASAP7_75t_L g329 ( .A(n_234), .Y(n_329) );
OR2x2_ASAP7_75t_L g350 ( .A(n_234), .B(n_334), .Y(n_350) );
OR2x2_ASAP7_75t_L g364 ( .A(n_234), .B(n_244), .Y(n_364) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_234), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_234), .B(n_286), .Y(n_436) );
OR2x6_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
INVx1_ASAP7_75t_L g281 ( .A(n_242), .Y(n_281) );
AND2x2_ASAP7_75t_L g414 ( .A(n_242), .B(n_280), .Y(n_414) );
AND2x2_ASAP7_75t_L g439 ( .A(n_242), .B(n_269), .Y(n_439) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g257 ( .A(n_244), .Y(n_257) );
BUFx3_ASAP7_75t_L g299 ( .A(n_244), .Y(n_299) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_244), .Y(n_326) );
INVx1_ASAP7_75t_L g335 ( .A(n_244), .Y(n_335) );
AOI33xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .A3(n_258), .B1(n_259), .B2(n_260), .B3(n_261), .Y(n_250) );
AOI21x1_ASAP7_75t_SL g353 ( .A1(n_251), .A2(n_275), .B(n_337), .Y(n_353) );
INVx2_ASAP7_75t_L g383 ( .A(n_251), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_251), .B(n_382), .Y(n_389) );
AND2x2_ASAP7_75t_L g337 ( .A(n_252), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g300 ( .A(n_255), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g401 ( .A(n_256), .Y(n_401) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_257), .Y(n_391) );
OAI32xp33_ASAP7_75t_L g440 ( .A1(n_258), .A2(n_260), .A3(n_436), .B1(n_441), .B2(n_443), .Y(n_440) );
AND2x2_ASAP7_75t_L g358 ( .A(n_259), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_SL g348 ( .A(n_260), .Y(n_348) );
AND2x2_ASAP7_75t_L g413 ( .A(n_260), .B(n_357), .Y(n_413) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI221xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_274), .B1(n_277), .B2(n_291), .C(n_295), .Y(n_264) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_268), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_269), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_269), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_269), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g318 ( .A(n_273), .Y(n_318) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR3xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_282), .C(n_287), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_279), .A2(n_341), .B1(n_381), .B2(n_384), .Y(n_380) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g284 ( .A(n_280), .Y(n_284) );
NOR2x1p5_ASAP7_75t_L g298 ( .A(n_280), .B(n_299), .Y(n_298) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_280), .Y(n_320) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI322xp33_ASAP7_75t_L g347 ( .A1(n_283), .A2(n_325), .A3(n_348), .B1(n_349), .B2(n_350), .C1(n_351), .C2(n_353), .Y(n_347) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_285), .A2(n_304), .B(n_305), .C(n_307), .Y(n_303) );
OR2x2_ASAP7_75t_L g395 ( .A(n_285), .B(n_349), .Y(n_395) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g302 ( .A(n_286), .B(n_290), .Y(n_302) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g308 ( .A(n_292), .B(n_309), .Y(n_308) );
INVx3_ASAP7_75t_SL g340 ( .A(n_293), .Y(n_340) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_297), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_SL g344 ( .A(n_300), .Y(n_344) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_301), .Y(n_386) );
OR2x6_ASAP7_75t_SL g441 ( .A(n_304), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI211xp5_ASAP7_75t_L g431 ( .A1(n_309), .A2(n_432), .B(n_433), .C(n_440), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_313), .B(n_316), .C(n_320), .Y(n_310) );
OAI211xp5_ASAP7_75t_SL g322 ( .A1(n_311), .A2(n_323), .B(n_330), .C(n_354), .Y(n_322) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
NOR3xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_367), .C(n_411), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_326), .Y(n_418) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
NOR3xp33_ASAP7_75t_SL g330 ( .A(n_331), .B(n_343), .C(n_347), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_336), .B1(n_339), .B2(n_342), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_335), .Y(n_442) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_SL g428 ( .A(n_341), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
OR2x2_ASAP7_75t_L g378 ( .A(n_344), .B(n_364), .Y(n_378) );
OR2x2_ASAP7_75t_L g429 ( .A(n_344), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g427 ( .A(n_352), .Y(n_427) );
OR2x2_ASAP7_75t_L g443 ( .A(n_352), .B(n_382), .Y(n_443) );
OAI21xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B(n_360), .Y(n_354) );
OAI31xp33_ASAP7_75t_L g368 ( .A1(n_355), .A2(n_369), .A3(n_370), .B(n_372), .Y(n_368) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g400 ( .A(n_365), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND4xp25_ASAP7_75t_SL g367 ( .A(n_368), .B(n_376), .C(n_387), .D(n_392), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_375), .Y(n_410) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B1(n_400), .B2(n_402), .C(n_404), .Y(n_392) );
NAND2xp33_ASAP7_75t_SL g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g437 ( .A(n_396), .Y(n_437) );
AND2x2_ASAP7_75t_SL g396 ( .A(n_397), .B(n_399), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_412), .B(n_431), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_415), .B2(n_417), .C(n_421), .Y(n_412) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_426), .B(n_429), .Y(n_421) );
INVxp33_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_437), .B2(n_438), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVxp33_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NOR2x1_ASAP7_75t_R g462 ( .A(n_452), .B(n_457), .Y(n_462) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_452), .Y(n_474) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_454), .B(n_466), .C(n_471), .Y(n_465) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_782), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_777), .Y(n_475) );
CKINVDCx11_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
BUFx4f_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
CKINVDCx11_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_SL g784 ( .A(n_483), .Y(n_784) );
AND2x4_ASAP7_75t_SL g483 ( .A(n_484), .B(n_673), .Y(n_483) );
NOR3xp33_ASAP7_75t_SL g484 ( .A(n_485), .B(n_582), .C(n_614), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_510), .B1(n_539), .B2(n_556), .C(n_567), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_496), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g545 ( .A(n_488), .B(n_497), .Y(n_545) );
INVx4_ASAP7_75t_L g573 ( .A(n_488), .Y(n_573) );
AND2x4_ASAP7_75t_SL g613 ( .A(n_488), .B(n_547), .Y(n_613) );
BUFx2_ASAP7_75t_L g623 ( .A(n_488), .Y(n_623) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_488), .B(n_628), .Y(n_689) );
AND2x2_ASAP7_75t_L g698 ( .A(n_488), .B(n_626), .Y(n_698) );
OR2x2_ASAP7_75t_L g706 ( .A(n_488), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g732 ( .A(n_488), .B(n_571), .Y(n_732) );
AND2x4_ASAP7_75t_L g751 ( .A(n_488), .B(n_752), .Y(n_751) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_495), .Y(n_488) );
INVx2_ASAP7_75t_SL g664 ( .A(n_496), .Y(n_664) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_505), .Y(n_496) );
AND2x2_ASAP7_75t_L g571 ( .A(n_497), .B(n_548), .Y(n_571) );
INVx2_ASAP7_75t_L g598 ( .A(n_497), .Y(n_598) );
INVx2_ASAP7_75t_L g628 ( .A(n_497), .Y(n_628) );
AND2x2_ASAP7_75t_L g642 ( .A(n_497), .B(n_547), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
AND2x2_ASAP7_75t_L g572 ( .A(n_505), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g595 ( .A(n_505), .Y(n_595) );
BUFx3_ASAP7_75t_L g609 ( .A(n_505), .Y(n_609) );
AND2x2_ASAP7_75t_L g638 ( .A(n_505), .B(n_639), .Y(n_638) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
AND2x4_ASAP7_75t_L g543 ( .A(n_506), .B(n_507), .Y(n_543) );
INVx1_ASAP7_75t_L g644 ( .A(n_510), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
OR2x2_ASAP7_75t_L g755 ( .A(n_511), .B(n_556), .Y(n_755) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g611 ( .A(n_512), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_512), .B(n_521), .Y(n_672) );
OR2x2_ASAP7_75t_L g770 ( .A(n_512), .B(n_692), .Y(n_770) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g581 ( .A(n_513), .B(n_557), .Y(n_581) );
OR2x2_ASAP7_75t_SL g591 ( .A(n_513), .B(n_592), .Y(n_591) );
INVx4_ASAP7_75t_L g602 ( .A(n_513), .Y(n_602) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_513), .Y(n_653) );
NAND2x1_ASAP7_75t_L g659 ( .A(n_513), .B(n_558), .Y(n_659) );
AND2x2_ASAP7_75t_L g684 ( .A(n_513), .B(n_523), .Y(n_684) );
OR2x2_ASAP7_75t_L g705 ( .A(n_513), .B(n_588), .Y(n_705) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_L g693 ( .A1(n_521), .A2(n_694), .B(n_697), .C(n_699), .Y(n_693) );
AND2x2_ASAP7_75t_L g766 ( .A(n_521), .B(n_542), .Y(n_766) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_530), .Y(n_521) );
INVx1_ASAP7_75t_L g633 ( .A(n_522), .Y(n_633) );
AND2x2_ASAP7_75t_L g703 ( .A(n_522), .B(n_558), .Y(n_703) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g577 ( .A(n_523), .Y(n_577) );
OR2x2_ASAP7_75t_L g592 ( .A(n_523), .B(n_558), .Y(n_592) );
INVx1_ASAP7_75t_L g608 ( .A(n_523), .Y(n_608) );
AND2x2_ASAP7_75t_L g620 ( .A(n_523), .B(n_530), .Y(n_620) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_523), .Y(n_726) );
NOR2x1_ASAP7_75t_SL g557 ( .A(n_530), .B(n_558), .Y(n_557) );
AO21x1_ASAP7_75t_SL g530 ( .A1(n_531), .A2(n_532), .B(n_538), .Y(n_530) );
AO21x2_ASAP7_75t_L g589 ( .A1(n_531), .A2(n_532), .B(n_538), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_537), .Y(n_532) );
INVxp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .Y(n_540) );
OR2x2_ASAP7_75t_L g690 ( .A(n_541), .B(n_625), .Y(n_690) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_542), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g772 ( .A(n_542), .B(n_669), .Y(n_772) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g617 ( .A(n_543), .B(n_598), .Y(n_617) );
AND2x2_ASAP7_75t_L g713 ( .A(n_543), .B(n_626), .Y(n_713) );
INVx1_ASAP7_75t_L g630 ( .A(n_544), .Y(n_630) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g680 ( .A(n_545), .Y(n_680) );
INVx2_ASAP7_75t_L g647 ( .A(n_546), .Y(n_647) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g597 ( .A(n_547), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g627 ( .A(n_547), .Y(n_627) );
INVx1_ASAP7_75t_L g752 ( .A(n_547), .Y(n_752) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_548), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
OR2x2_ASAP7_75t_L g723 ( .A(n_556), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g578 ( .A(n_558), .Y(n_578) );
OR2x2_ASAP7_75t_L g601 ( .A(n_558), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g612 ( .A(n_558), .B(n_588), .Y(n_612) );
AND2x2_ASAP7_75t_L g686 ( .A(n_558), .B(n_602), .Y(n_686) );
BUFx2_ASAP7_75t_L g769 ( .A(n_558), .Y(n_769) );
OR2x6_ASAP7_75t_L g558 ( .A(n_559), .B(n_566), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_574), .B(n_579), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
AND2x2_ASAP7_75t_L g721 ( .A(n_570), .B(n_643), .Y(n_721) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g580 ( .A(n_571), .B(n_573), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_572), .B(n_642), .Y(n_743) );
INVx1_ASAP7_75t_L g773 ( .A(n_572), .Y(n_773) );
NAND2x1p5_ASAP7_75t_L g669 ( .A(n_573), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_573), .B(n_709), .Y(n_746) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
AND2x4_ASAP7_75t_SL g610 ( .A(n_576), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_576), .B(n_604), .Y(n_757) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_577), .B(n_659), .Y(n_715) );
AND2x2_ASAP7_75t_L g733 ( .A(n_577), .B(n_686), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_578), .B(n_620), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_578), .A2(n_624), .B(n_666), .C(n_671), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_578), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_580), .A2(n_653), .B1(n_761), .B2(n_767), .C(n_771), .Y(n_760) );
INVx1_ASAP7_75t_SL g748 ( .A(n_581), .Y(n_748) );
OAI221xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_593), .B1(n_599), .B2(n_603), .C(n_789), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g658 ( .A(n_587), .Y(n_658) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g632 ( .A(n_588), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g663 ( .A(n_588), .B(n_608), .Y(n_663) );
INVx2_ASAP7_75t_L g696 ( .A(n_588), .Y(n_696) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OAI32xp33_ASAP7_75t_L g747 ( .A1(n_591), .A2(n_638), .A3(n_669), .B1(n_748), .B2(n_749), .Y(n_747) );
OR2x2_ASAP7_75t_L g718 ( .A(n_592), .B(n_705), .Y(n_718) );
INVx1_ASAP7_75t_L g728 ( .A(n_593), .Y(n_728) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx2_ASAP7_75t_L g643 ( .A(n_594), .Y(n_643) );
AND2x2_ASAP7_75t_L g714 ( .A(n_594), .B(n_689), .Y(n_714) );
OR2x2_ASAP7_75t_L g745 ( .A(n_594), .B(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_595), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g639 ( .A(n_598), .Y(n_639) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx2_ASAP7_75t_SL g604 ( .A(n_601), .Y(n_604) );
OR2x2_ASAP7_75t_L g691 ( .A(n_601), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_602), .B(n_620), .Y(n_619) );
NOR2xp67_ASAP7_75t_L g725 ( .A(n_602), .B(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g738 ( .A(n_602), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B(n_610), .C(n_613), .Y(n_603) );
AND2x2_ASAP7_75t_L g753 ( .A(n_605), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g679 ( .A(n_609), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_609), .B(n_613), .Y(n_700) );
AND2x2_ASAP7_75t_L g731 ( .A(n_609), .B(n_732), .Y(n_731) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_611), .A2(n_742), .B(n_744), .C(n_747), .Y(n_741) );
AOI222xp33_ASAP7_75t_L g615 ( .A1(n_612), .A2(n_616), .B1(n_618), .B2(n_621), .C1(n_629), .C2(n_631), .Y(n_615) );
AND2x2_ASAP7_75t_L g683 ( .A(n_612), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g616 ( .A(n_613), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g637 ( .A(n_613), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g614 ( .A(n_615), .B(n_634), .C(n_655), .D(n_665), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_617), .B(n_623), .Y(n_677) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g685 ( .A(n_620), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g692 ( .A(n_620), .Y(n_692) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_622), .A2(n_656), .B(n_660), .C(n_664), .Y(n_655) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_623), .B(n_638), .Y(n_759) );
OR2x2_ASAP7_75t_L g763 ( .A(n_623), .B(n_649), .Y(n_763) );
INVx1_ASAP7_75t_L g736 ( .A(n_624), .Y(n_736) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_SL g670 ( .A(n_627), .Y(n_670) );
INVx1_ASAP7_75t_L g650 ( .A(n_628), .Y(n_650) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_630), .B(n_667), .Y(n_666) );
BUFx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g654 ( .A(n_632), .Y(n_654) );
AOI322xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .A3(n_638), .B1(n_640), .B2(n_644), .C1(n_645), .C2(n_651), .Y(n_634) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_SL g716 ( .A1(n_637), .A2(n_717), .B(n_718), .C(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g739 ( .A(n_638), .Y(n_739) );
NOR2xp67_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g697 ( .A(n_643), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_649), .Y(n_719) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx3_ASAP7_75t_L g662 ( .A(n_659), .Y(n_662) );
OR2x2_ASAP7_75t_L g730 ( .A(n_659), .B(n_692), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_659), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_SL g762 ( .A(n_663), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_664), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND3xp33_ASAP7_75t_SL g767 ( .A(n_672), .B(n_768), .C(n_770), .Y(n_767) );
NOR3xp33_ASAP7_75t_SL g673 ( .A(n_674), .B(n_711), .C(n_740), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_675), .B(n_693), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B(n_681), .C(n_687), .Y(n_675) );
OAI31xp33_ASAP7_75t_L g720 ( .A1(n_676), .A2(n_698), .A3(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx2_ASAP7_75t_L g735 ( .A(n_683), .Y(n_735) );
INVx1_ASAP7_75t_L g710 ( .A(n_685), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g737 ( .A(n_695), .B(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g776 ( .A(n_696), .Y(n_776) );
OAI22xp33_ASAP7_75t_SL g699 ( .A1(n_700), .A2(n_701), .B1(n_706), .B2(n_710), .Y(n_699) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_705), .Y(n_717) );
OR2x2_ASAP7_75t_L g768 ( .A(n_705), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_712), .B(n_720), .C(n_727), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B(n_715), .C(n_716), .Y(n_712) );
INVx2_ASAP7_75t_L g749 ( .A(n_713), .Y(n_749) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_731), .B2(n_733), .C(n_734), .Y(n_727) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_737), .B2(n_739), .Y(n_734) );
NAND3xp33_ASAP7_75t_SL g740 ( .A(n_741), .B(n_750), .C(n_760), .Y(n_740) );
INVxp33_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_753), .B1(n_756), .B2(n_758), .Y(n_750) );
INVx2_ASAP7_75t_L g764 ( .A(n_751), .Y(n_764) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_761) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI22xp33_ASAP7_75t_SL g771 ( .A1(n_770), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp33_ASAP7_75t_SL g782 ( .A(n_777), .B(n_783), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
endmodule