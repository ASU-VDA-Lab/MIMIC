module fake_jpeg_9634_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_34),
.B(n_20),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_16),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_28),
.B1(n_21),
.B2(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_69),
.B1(n_71),
.B2(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_57),
.Y(n_80)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_33),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_26),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_28),
.B1(n_37),
.B2(n_36),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_41),
.B1(n_36),
.B2(n_44),
.Y(n_77)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_28),
.B1(n_33),
.B2(n_30),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_41),
.B1(n_36),
.B2(n_30),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_88),
.B1(n_67),
.B2(n_25),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_91),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_63),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_36),
.B1(n_44),
.B2(n_40),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_35),
.B1(n_42),
.B2(n_39),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_24),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_21),
.B1(n_30),
.B2(n_24),
.Y(n_88)
);

OAI22x1_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_35),
.B1(n_31),
.B2(n_23),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_40),
.B1(n_21),
.B2(n_25),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_32),
.B1(n_18),
.B2(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_61),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_98),
.Y(n_126)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_99),
.A2(n_103),
.B1(n_110),
.B2(n_111),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_105),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_79),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_106),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_59),
.B1(n_52),
.B2(n_63),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_59),
.B1(n_48),
.B2(n_60),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_108),
.B1(n_113),
.B2(n_114),
.Y(n_127)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_80),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_57),
.B(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_81),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_75),
.B(n_86),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_73),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_35),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_54),
.B1(n_46),
.B2(n_56),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_81),
.B1(n_91),
.B2(n_82),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_76),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_142),
.B(n_147),
.Y(n_154)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_79),
.B(n_77),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_39),
.B(n_96),
.Y(n_171)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_89),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_118),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_106),
.B1(n_116),
.B2(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_83),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_108),
.Y(n_144)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_73),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_149),
.A2(n_171),
.B1(n_130),
.B2(n_70),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_115),
.B1(n_112),
.B2(n_81),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_150),
.A2(n_166),
.B1(n_143),
.B2(n_133),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_102),
.B1(n_99),
.B2(n_32),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_151),
.A2(n_153),
.B(n_161),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_84),
.B(n_22),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_156),
.B(n_174),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_84),
.B1(n_46),
.B2(n_107),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_159),
.B1(n_125),
.B2(n_123),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_35),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_172),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_107),
.B1(n_85),
.B2(n_69),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_22),
.B(n_26),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_123),
.A2(n_85),
.B1(n_18),
.B2(n_22),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_18),
.B(n_26),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_135),
.B(n_137),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_16),
.B1(n_17),
.B2(n_29),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_151),
.B1(n_166),
.B2(n_165),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_39),
.C(n_53),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_39),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_126),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_53),
.C(n_96),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_176),
.A2(n_183),
.B(n_188),
.Y(n_208)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_180),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_157),
.B1(n_165),
.B2(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_144),
.B1(n_128),
.B2(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_122),
.B1(n_127),
.B2(n_134),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_137),
.B1(n_163),
.B2(n_132),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_127),
.B1(n_124),
.B2(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_194),
.B(n_195),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_16),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_87),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_200),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_130),
.B(n_16),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_31),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_154),
.A2(n_152),
.B1(n_172),
.B2(n_161),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_155),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_154),
.B(n_158),
.Y(n_205)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_189),
.B(n_192),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_155),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_207),
.C(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_177),
.C(n_201),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_215),
.C(n_219),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_168),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_7),
.B1(n_14),
.B2(n_12),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_29),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_197),
.B1(n_186),
.B2(n_17),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_130),
.C(n_65),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_29),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_17),
.C(n_19),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_241),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_225),
.A2(n_184),
.B1(n_176),
.B2(n_193),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_230),
.B1(n_236),
.B2(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_194),
.B1(n_192),
.B2(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_235),
.B(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_238),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_55),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_206),
.C(n_214),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_212),
.Y(n_240)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_211),
.A2(n_7),
.B1(n_14),
.B2(n_11),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_242),
.A2(n_215),
.B1(n_222),
.B2(n_8),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_203),
.A2(n_223),
.B1(n_217),
.B2(n_208),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_208),
.B(n_0),
.CI(n_1),
.CON(n_244),
.SN(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_245),
.Y(n_259)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_6),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_246),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_209),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_251),
.C(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_210),
.Y(n_251)
);

BUFx12f_ASAP7_75t_SL g256 ( 
.A(n_226),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_244),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_205),
.B(n_202),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_244),
.B(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_207),
.B1(n_2),
.B2(n_3),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_241),
.B1(n_242),
.B2(n_231),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_1),
.C(n_2),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_264),
.C(n_6),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_8),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_265),
.B(n_268),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_230),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_272),
.C(n_279),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_278),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_274),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_275),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_237),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_276),
.A2(n_277),
.B1(n_250),
.B2(n_257),
.Y(n_281)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_8),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_258),
.B(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_249),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_290),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_264),
.C(n_263),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_288),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_252),
.C(n_261),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_252),
.B(n_250),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_10),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_6),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_272),
.B(n_279),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_296),
.B(n_282),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_9),
.Y(n_293)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_9),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_298),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_15),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_302),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_290),
.B(n_283),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_299),
.B(n_294),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_3),
.C(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_283),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_306),
.B(n_307),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_288),
.Y(n_307)
);

OAI311xp33_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_303),
.A3(n_301),
.B1(n_5),
.C1(n_4),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_312),
.B(n_4),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_3),
.C(n_4),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_311),
.B(n_308),
.Y(n_316)
);

O2A1O1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_5),
.B(n_314),
.C(n_309),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_5),
.Y(n_318)
);


endmodule