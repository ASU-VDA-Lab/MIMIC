module fake_jpeg_2479_n_165 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_56),
.Y(n_75)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_45),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_59),
.B1(n_44),
.B2(n_49),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_47),
.B(n_58),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_60),
.B1(n_62),
.B2(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_53),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_62),
.B1(n_59),
.B2(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_51),
.B1(n_56),
.B2(n_47),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_44),
.B1(n_52),
.B2(n_50),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_72),
.B1(n_61),
.B2(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_19),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_3),
.C(n_4),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_113)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_0),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_1),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_91),
.B(n_93),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_23),
.B(n_36),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_20),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_107),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_111),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_108),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_3),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_119),
.B1(n_123),
.B2(n_120),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_40),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_5),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_24),
.B(n_35),
.C(n_32),
.Y(n_123)
);

INVx2_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_126),
.B(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_10),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_120),
.C(n_114),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_99),
.B1(n_104),
.B2(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_99),
.B1(n_13),
.B2(n_12),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_14),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_135),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_118),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_132),
.B1(n_124),
.B2(n_116),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_146),
.B(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_155),
.C(n_158),
.Y(n_161)
);

NOR4xp25_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_144),
.C(n_156),
.D(n_154),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_149),
.B(n_144),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_153),
.B(n_152),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_137),
.Y(n_165)
);


endmodule