module real_jpeg_7124_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_1),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_1),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_1),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_1),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_1),
.B(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_3),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_3),
.B(n_114),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_3),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_4),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_4),
.B(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_4),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_4),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_4),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_4),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_5),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_5),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_5),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_5),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_5),
.B(n_38),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_5),
.B(n_454),
.Y(n_453)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_7),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_7),
.Y(n_343)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_8),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_8),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g436 ( 
.A(n_8),
.Y(n_436)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_10),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_10),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_10),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_11),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_11),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_11),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_11),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_11),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_11),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g421 ( 
.A(n_11),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_12),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_12),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_12),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_12),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_12),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_12),
.B(n_341),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_13),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_14),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_14),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_14),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_14),
.B(n_315),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_14),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_14),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_43),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_15),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_15),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_15),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_15),
.B(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_15),
.B(n_38),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_15),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_15),
.B(n_457),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_442),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_412),
.B(n_441),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_302),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_221),
.B(n_262),
.C(n_263),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_193),
.B(n_220),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_22),
.B(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_154),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_23),
.B(n_154),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_105),
.C(n_137),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_24),
.B(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_72),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_25),
.B(n_73),
.C(n_86),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_48),
.C(n_62),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_26),
.B(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_36),
.B2(n_41),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_28),
.A2(n_29),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_28),
.A2(n_29),
.B1(n_74),
.B2(n_75),
.Y(n_464)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_29),
.B(n_36),
.C(n_42),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_29),
.B(n_202),
.C(n_421),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_50),
.Y(n_49)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_30),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_30),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_35),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_35),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_35),
.Y(n_322)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_35),
.Y(n_351)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_39),
.Y(n_162)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_40),
.Y(n_136)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_40),
.Y(n_207)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g312 ( 
.A(n_47),
.Y(n_312)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_47),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_48),
.A2(n_62),
.B1(n_63),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_48),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.C(n_56),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_49),
.A2(n_56),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_49),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_49),
.A2(n_202),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_49),
.A2(n_202),
.B1(n_421),
.B2(n_424),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_49),
.B(n_126),
.C(n_272),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_50),
.B(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_50),
.Y(n_165)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_51),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_52),
.B(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_54),
.B(n_101),
.Y(n_208)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_56),
.Y(n_203)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_60),
.Y(n_213)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_60),
.Y(n_256)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_61),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_61),
.Y(n_285)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_64),
.A2(n_172),
.B1(n_173),
.B2(n_175),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_64),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_64),
.A2(n_68),
.B1(n_69),
.B2(n_175),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_64),
.B(n_173),
.C(n_176),
.Y(n_260)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_67),
.Y(n_338)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_67),
.Y(n_361)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_71),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_86),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_75),
.B(n_80),
.C(n_84),
.Y(n_192)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_81),
.B(n_126),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_88),
.B(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_87),
.B(n_95),
.C(n_100),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_93),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_98),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_105),
.B(n_137),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_121),
.C(n_123),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_106),
.A2(n_121),
.B1(n_122),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_113),
.C(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_108),
.B(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_108),
.B(n_377),
.Y(n_376)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_111),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_117),
.A2(n_118),
.B1(n_241),
.B2(n_245),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_118),
.B(n_173),
.C(n_242),
.Y(n_297)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_123),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.C(n_133),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_124),
.A2(n_125),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_126),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_126),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_126),
.A2(n_230),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_126),
.B(n_233),
.C(n_239),
.Y(n_277)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_400)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_153),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_140),
.C(n_153),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_147),
.C(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_147),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_147),
.Y(n_287)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_157),
.C(n_180),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_180),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_169),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_159),
.B(n_160),
.C(n_169),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_161),
.Y(n_228)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_162),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_164),
.B(n_166),
.C(n_228),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_176),
.B2(n_179),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_172),
.A2(n_173),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_172),
.A2(n_173),
.B1(n_310),
.B2(n_311),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_173),
.B(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_174),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_176),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_176),
.A2(n_179),
.B1(n_438),
.B2(n_439),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_179),
.B(n_433),
.C(n_438),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_181),
.B(n_183),
.C(n_184),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_189),
.C(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_188),
.Y(n_281)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_218),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_194),
.B(n_218),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.C(n_215),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_195),
.A2(n_196),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_199),
.B(n_215),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.C(n_214),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_200),
.B(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_204),
.B(n_214),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.C(n_209),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_208),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_209),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_210),
.B(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_210),
.B(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_222),
.B(n_264),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_224),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_265),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_224),
.B(n_265),
.Y(n_411)
);

FAx1_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_246),
.CI(n_261),
.CON(n_224),
.SN(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_240),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_227),
.B(n_229),
.C(n_240),
.Y(n_291)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_239),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_236),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_236),
.A2(n_239),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_249),
.C(n_251),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_260),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_259),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_257),
.C(n_260),
.Y(n_294)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_257),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_257),
.A2(n_259),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_259),
.B(n_296),
.C(n_301),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_266),
.B(n_268),
.C(n_289),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_289),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_276),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_269),
.B(n_277),
.C(n_278),
.Y(n_440)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_288),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_280),
.B(n_283),
.C(n_287),
.Y(n_428)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_290),
.B(n_294),
.C(n_295),
.Y(n_415)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

AO22x1_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

OAI31xp33_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_408),
.A3(n_409),
.B(n_411),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_402),
.B(n_407),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_389),
.B(n_401),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_345),
.B(n_388),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_330),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_307),
.B(n_330),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_308),
.B(n_318),
.C(n_327),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_309),
.B(n_314),
.C(n_316),
.Y(n_397)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_327),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.C(n_325),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_319),
.B(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.C(n_344),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_331),
.B(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_333),
.A2(n_334),
.B1(n_344),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_335),
.A2(n_336),
.B1(n_339),
.B2(n_340),
.Y(n_354)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_382),
.B(n_387),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_366),
.B(n_381),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_355),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_355),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_354),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_362),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_357),
.B1(n_362),
.B2(n_363),
.Y(n_379)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_375),
.B(n_380),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_376),
.B(n_379),
.Y(n_380)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_384),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_391),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_395),
.B2(n_396),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_397),
.C(n_398),
.Y(n_406)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_406),
.Y(n_407)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_404),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_414),
.Y(n_441)
);

BUFx24_ASAP7_75t_SL g468 ( 
.A(n_414),
.Y(n_468)
);

FAx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_416),
.CI(n_429),
.CON(n_414),
.SN(n_414)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_416),
.C(n_429),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_425),
.B2(n_426),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_427),
.C(n_428),
.Y(n_448)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_421),
.Y(n_424)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_440),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_432),
.C(n_440),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_437),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_438),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_465),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_444),
.B(n_445),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_460),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_453),
.A2(n_456),
.B1(n_458),
.B2(n_459),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_453),
.Y(n_458)
);

INVx6_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_456),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);


endmodule