module fake_ibex_819_n_219 (n_60, n_49, n_70, n_7, n_20, n_40, n_17, n_66, n_69, n_74, n_75, n_25, n_36, n_58, n_41, n_48, n_43, n_57, n_59, n_18, n_3, n_22, n_28, n_32, n_39, n_53, n_65, n_4, n_73, n_33, n_54, n_5, n_11, n_30, n_6, n_50, n_62, n_71, n_64, n_72, n_55, n_63, n_29, n_68, n_13, n_2, n_8, n_26, n_61, n_35, n_14, n_0, n_67, n_9, n_34, n_12, n_38, n_42, n_15, n_37, n_24, n_52, n_47, n_31, n_44, n_10, n_23, n_21, n_51, n_56, n_27, n_46, n_45, n_19, n_16, n_1, n_219);

input n_60;
input n_49;
input n_70;
input n_7;
input n_20;
input n_40;
input n_17;
input n_66;
input n_69;
input n_74;
input n_75;
input n_25;
input n_36;
input n_58;
input n_41;
input n_48;
input n_43;
input n_57;
input n_59;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_39;
input n_53;
input n_65;
input n_4;
input n_73;
input n_33;
input n_54;
input n_5;
input n_11;
input n_30;
input n_6;
input n_50;
input n_62;
input n_71;
input n_64;
input n_72;
input n_55;
input n_63;
input n_29;
input n_68;
input n_13;
input n_2;
input n_8;
input n_26;
input n_61;
input n_35;
input n_14;
input n_0;
input n_67;
input n_9;
input n_34;
input n_12;
input n_38;
input n_42;
input n_15;
input n_37;
input n_24;
input n_52;
input n_47;
input n_31;
input n_44;
input n_10;
input n_23;
input n_21;
input n_51;
input n_56;
input n_27;
input n_46;
input n_45;
input n_19;
input n_16;
input n_1;

output n_219;

wire n_151;
wire n_147;
wire n_85;
wire n_167;
wire n_128;
wire n_208;
wire n_84;
wire n_171;
wire n_152;
wire n_145;
wire n_103;
wire n_95;
wire n_205;
wire n_204;
wire n_139;
wire n_130;
wire n_129;
wire n_161;
wire n_98;
wire n_143;
wire n_106;
wire n_177;
wire n_203;
wire n_148;
wire n_76;
wire n_118;
wire n_183;
wire n_209;
wire n_164;
wire n_198;
wire n_124;
wire n_193;
wire n_110;
wire n_169;
wire n_108;
wire n_217;
wire n_82;
wire n_165;
wire n_78;
wire n_86;
wire n_87;
wire n_109;
wire n_121;
wire n_127;
wire n_175;
wire n_137;
wire n_125;
wire n_191;
wire n_178;
wire n_153;
wire n_173;
wire n_120;
wire n_93;
wire n_168;
wire n_155;
wire n_162;
wire n_194;
wire n_180;
wire n_122;
wire n_116;
wire n_201;
wire n_134;
wire n_94;
wire n_77;
wire n_112;
wire n_150;
wire n_88;
wire n_133;
wire n_142;
wire n_80;
wire n_215;
wire n_172;
wire n_90;
wire n_176;
wire n_192;
wire n_140;
wire n_216;
wire n_136;
wire n_119;
wire n_100;
wire n_179;
wire n_206;
wire n_166;
wire n_195;
wire n_163;
wire n_212;
wire n_188;
wire n_200;
wire n_114;
wire n_199;
wire n_97;
wire n_102;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_189;
wire n_99;
wire n_135;
wire n_156;
wire n_187;
wire n_126;
wire n_105;
wire n_154;
wire n_182;
wire n_111;
wire n_196;
wire n_104;
wire n_141;
wire n_89;
wire n_83;
wire n_107;
wire n_115;
wire n_149;
wire n_186;
wire n_92;
wire n_170;
wire n_144;
wire n_213;
wire n_101;
wire n_190;
wire n_113;
wire n_138;
wire n_96;
wire n_185;
wire n_117;
wire n_214;
wire n_79;
wire n_81;
wire n_159;
wire n_202;
wire n_158;
wire n_211;
wire n_218;
wire n_132;
wire n_174;
wire n_210;
wire n_157;
wire n_160;
wire n_184;
wire n_146;
wire n_91;
wire n_207;

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_11),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g84 ( 
.A(n_36),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_1),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_14),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_74),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_10),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_70),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_23),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_43),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_44),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_7),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_64),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_50),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_5),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_52),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_37),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_71),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_49),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_25),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_34),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_16),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_53),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_27),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_15),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_12),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_8),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_17),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_40),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_18),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_42),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_22),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_3),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_6),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_87),
.B(n_0),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_0),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_123),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_77),
.B(n_28),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_31),
.B1(n_38),
.B2(n_48),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_80),
.B(n_51),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_102),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_125),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_66),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_108),
.B(n_72),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_91),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_86),
.B(n_73),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_101),
.B(n_106),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_132),
.Y(n_170)
);

AND2x4_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_112),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_79),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_149),
.B(n_76),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_97),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_121),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_113),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_134),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_169),
.B(n_126),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_159),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_81),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_85),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_166),
.B(n_100),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_130),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_98),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_127),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_157),
.B(n_154),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_158),
.B1(n_144),
.B2(n_155),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_142),
.Y(n_192)
);

AO32x2_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_147),
.A3(n_105),
.B1(n_120),
.B2(n_143),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_189),
.B(n_181),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_148),
.B(n_124),
.C(n_90),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_185),
.B(n_184),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_179),
.Y(n_197)
);

AND2x4_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_178),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_196),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_177),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_R g201 ( 
.A(n_193),
.B(n_89),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_175),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_110),
.B1(n_93),
.B2(n_94),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_201),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_131),
.B1(n_95),
.B2(n_99),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

OAI211xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_195),
.B(n_137),
.C(n_139),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_R g213 ( 
.A(n_212),
.B(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_199),
.B1(n_152),
.B2(n_210),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_214),
.A2(n_152),
.B1(n_202),
.B2(n_204),
.Y(n_217)
);

AOI22x1_ASAP7_75t_SL g218 ( 
.A1(n_216),
.A2(n_193),
.B1(n_115),
.B2(n_118),
.Y(n_218)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_217),
.B1(n_172),
.B2(n_174),
.C(n_180),
.Y(n_219)
);


endmodule