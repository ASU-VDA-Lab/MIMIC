module fake_jpeg_3971_n_178 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_9),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_37),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_29),
.B1(n_22),
.B2(n_16),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_44),
.B1(n_27),
.B2(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_29),
.B1(n_16),
.B2(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_57),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_58),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_27),
.B(n_25),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_37),
.B1(n_36),
.B2(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_71),
.B1(n_25),
.B2(n_28),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_73),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_24),
.B(n_35),
.C(n_30),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_35),
.B(n_30),
.C(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_38),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_38),
.B1(n_21),
.B2(n_17),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_39),
.B1(n_49),
.B2(n_26),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_19),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_85),
.B1(n_89),
.B2(n_91),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_50),
.C(n_49),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_59),
.C(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_28),
.Y(n_87)
);

AOI22x1_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_56),
.B1(n_71),
.B2(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_0),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_39),
.B1(n_26),
.B2(n_21),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_65),
.B1(n_72),
.B2(n_58),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_114),
.C(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_54),
.B(n_66),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_93),
.B(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_113),
.B1(n_80),
.B2(n_84),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_57),
.A3(n_26),
.B1(n_21),
.B2(n_18),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_76),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_60),
.B1(n_26),
.B2(n_21),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_92),
.C(n_88),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_123),
.B(n_18),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_105),
.B1(n_106),
.B2(n_111),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_122),
.B1(n_99),
.B2(n_75),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_76),
.B1(n_91),
.B2(n_75),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_76),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_64),
.B1(n_3),
.B2(n_4),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_78),
.A3(n_77),
.B1(n_18),
.B2(n_17),
.Y(n_136)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_112),
.B(n_108),
.C(n_114),
.D(n_101),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_13),
.C(n_3),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_17),
.C(n_64),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_140),
.CI(n_123),
.CON(n_153),
.SN(n_153)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_139),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_103),
.B1(n_99),
.B2(n_104),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_137),
.B(n_142),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_84),
.B1(n_103),
.B2(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_104),
.A3(n_17),
.B1(n_18),
.B2(n_20),
.C(n_13),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_116),
.C(n_115),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_123),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_130),
.C(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_122),
.B1(n_119),
.B2(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_153),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_128),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_6),
.B(n_7),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_152),
.B1(n_7),
.B2(n_8),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_133),
.B1(n_131),
.B2(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_1),
.C(n_5),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_142),
.B(n_136),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_159),
.B(n_160),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_157),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_138),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_161),
.C(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_1),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_165),
.B(n_167),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_149),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_168),
.B(n_7),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_145),
.B1(n_150),
.B2(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_153),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_167),
.B(n_10),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_170),
.B(n_12),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_174),
.C(n_175),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_12),
.Y(n_178)
);


endmodule