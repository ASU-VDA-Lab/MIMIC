module real_jpeg_13638_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_202;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_4),
.A2(n_26),
.B1(n_44),
.B2(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_4),
.A2(n_26),
.B1(n_55),
.B2(n_57),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_4),
.B(n_31),
.C(n_34),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_32),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_4),
.B(n_41),
.C(n_44),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_4),
.B(n_52),
.C(n_57),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_5),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_7),
.A2(n_38),
.B1(n_55),
.B2(n_57),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_14),
.B(n_263),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_10),
.B(n_264),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_11),
.A2(n_47),
.B1(n_55),
.B2(n_57),
.Y(n_84)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_259),
.B(n_261),
.Y(n_14)
);

AO21x1_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_68),
.B(n_258),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_66),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_17),
.B(n_66),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_61),
.C(n_62),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_18),
.A2(n_19),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.C(n_48),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_20),
.A2(n_21),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_20),
.B(n_76),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_20),
.A2(n_21),
.B1(n_89),
.B2(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_20),
.A2(n_21),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI211xp5_ASAP7_75t_SL g158 ( 
.A1(n_20),
.A2(n_85),
.B(n_106),
.C(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_20),
.A2(n_21),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_20),
.A2(n_89),
.B(n_113),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_20),
.A2(n_21),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_20),
.A2(n_21),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_21),
.B(n_77),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_21),
.B(n_49),
.C(n_234),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_21),
.B(n_243),
.C(n_247),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_22),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_24),
.B(n_141),
.Y(n_140)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_26),
.B(n_97),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_26),
.B(n_83),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_27),
.B(n_67),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_34),
.B(n_175),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_36),
.A2(n_48),
.B1(n_49),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_36),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_37),
.A2(n_39),
.B1(n_43),
.B2(n_78),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_43),
.B(n_46),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_39),
.A2(n_43),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OA22x2_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_43),
.Y(n_194)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_44),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_48),
.A2(n_49),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_60),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_59),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_58),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_58),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_55),
.B(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_61),
.B(n_62),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_66),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_66),
.B(n_260),
.Y(n_262)
);

OAI21x1_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_252),
.B(n_257),
.Y(n_68)
);

AOI21x1_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_226),
.B(n_249),
.Y(n_69)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_124),
.B(n_225),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_107),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_72),
.B(n_107),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_88),
.C(n_99),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_88),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_87),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_74),
.A2(n_75),
.B1(n_101),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_74),
.A2(n_75),
.B1(n_138),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_76),
.A2(n_77),
.B1(n_85),
.B2(n_134),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_142),
.C(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_76),
.A2(n_77),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_77),
.B(n_119),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_77),
.B(n_134),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_134),
.B(n_171),
.C(n_176),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_79),
.A2(n_100),
.B(n_105),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_80),
.A2(n_85),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_85),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_85),
.A2(n_102),
.B1(n_134),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_85),
.A2(n_134),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_85),
.A2(n_134),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_85),
.A2(n_134),
.B1(n_188),
.B2(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_85),
.B(n_142),
.C(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_85),
.B(n_178),
.C(n_182),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_98),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_93),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_105),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_105),
.B(n_138),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_123),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_117),
.B2(n_118),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_112),
.B(n_117),
.C(n_123),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_122),
.A2(n_230),
.B1(n_231),
.B2(n_236),
.Y(n_229)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_122),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_144),
.B(n_224),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_128),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_136),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_222)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_136),
.A2(n_137),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_143),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_142),
.A2(n_143),
.B1(n_153),
.B2(n_154),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_173),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_143),
.B1(n_191),
.B2(n_195),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_142),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_142),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_143),
.B(n_204),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_165),
.B(n_218),
.C(n_223),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_147),
.B(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_148),
.A2(n_149),
.B1(n_171),
.B2(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_161),
.C(n_163),
.Y(n_219)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_212),
.B(n_217),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_184),
.B(n_211),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_207),
.B(n_210),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_196),
.B(n_206),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_216),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_220),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_239),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_238),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_237),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_236),
.C(n_237),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_248),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_248),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_247),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_256),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);


endmodule