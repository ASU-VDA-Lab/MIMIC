module fake_jpeg_20425_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_48),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_44)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_48),
.Y(n_88)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_72),
.B(n_78),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_50),
.B(n_38),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_19),
.B(n_18),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_77),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_75),
.B(n_88),
.Y(n_133)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_47),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_20),
.B1(n_32),
.B2(n_27),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_32),
.B1(n_28),
.B2(n_44),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_91),
.B1(n_98),
.B2(n_38),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_92),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_64),
.B(n_40),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_49),
.C(n_46),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_28),
.B1(n_43),
.B2(n_32),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_49),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_28),
.B1(n_27),
.B2(n_31),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_26),
.Y(n_100)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_20),
.B1(n_36),
.B2(n_29),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_43),
.B1(n_31),
.B2(n_27),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_107),
.B1(n_120),
.B2(n_91),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_31),
.B1(n_38),
.B2(n_19),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_112),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_22),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_69),
.B1(n_97),
.B2(n_68),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_42),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_73),
.A2(n_21),
.B1(n_46),
.B2(n_45),
.Y(n_120)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_126),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_20),
.A3(n_19),
.B1(n_45),
.B2(n_42),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_46),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_90),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_21),
.B1(n_36),
.B2(n_29),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_139),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_140),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_80),
.B1(n_92),
.B2(n_89),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_143),
.B1(n_136),
.B2(n_139),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_111),
.A2(n_87),
.B1(n_86),
.B2(n_102),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_144),
.A2(n_157),
.B1(n_160),
.B2(n_162),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_42),
.Y(n_188)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_67),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_158),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_106),
.A2(n_76),
.B1(n_71),
.B2(n_67),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_109),
.B1(n_129),
.B2(n_121),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_69),
.B1(n_99),
.B2(n_70),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_70),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_160),
.A2(n_113),
.B1(n_128),
.B2(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_162),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_171),
.B1(n_176),
.B2(n_146),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_137),
.B1(n_153),
.B2(n_154),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_117),
.B1(n_113),
.B2(n_108),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_26),
.B1(n_22),
.B2(n_30),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_149),
.A2(n_131),
.B(n_112),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_173),
.A2(n_175),
.B(n_178),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_26),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_120),
.B(n_112),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_118),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_180),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_114),
.B(n_29),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_18),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_113),
.B(n_105),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_181),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_113),
.B(n_105),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_185),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_115),
.C(n_110),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_105),
.B(n_81),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_161),
.B(n_155),
.C(n_26),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_188),
.B(n_184),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_192),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_115),
.B1(n_123),
.B2(n_69),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_193),
.B1(n_141),
.B2(n_161),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_36),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_219),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_179),
.B1(n_182),
.B2(n_191),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_211),
.B(n_223),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_161),
.B1(n_18),
.B2(n_13),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_200),
.A2(n_203),
.B1(n_209),
.B2(n_215),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_22),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_163),
.A2(n_35),
.B1(n_25),
.B2(n_30),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_163),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_164),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

AO221x1_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_220),
.B1(n_221),
.B2(n_1),
.C(n_3),
.Y(n_247)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_217),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_165),
.B1(n_183),
.B2(n_189),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_190),
.B(n_11),
.Y(n_216)
);

OA21x2_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_209),
.B(n_186),
.Y(n_241)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_22),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_30),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_164),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_33),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_175),
.B(n_165),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_242),
.B(n_243),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_212),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_188),
.C(n_173),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_240),
.C(n_248),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_234),
.A2(n_199),
.B1(n_204),
.B2(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_181),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_206),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_180),
.C(n_178),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_246),
.C(n_9),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_179),
.B(n_192),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_10),
.B(n_11),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_33),
.B(n_2),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_251),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_9),
.C(n_16),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_35),
.C(n_25),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_251),
.A2(n_200),
.B1(n_203),
.B2(n_222),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_196),
.Y(n_254)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_215),
.CI(n_217),
.CON(n_256),
.SN(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_257),
.Y(n_273)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_260),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_272),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_269),
.B1(n_231),
.B2(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_206),
.Y(n_263)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_243),
.B1(n_199),
.B2(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_225),
.C(n_214),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_236),
.C(n_242),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_244),
.Y(n_289)
);

BUFx12_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_199),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_238),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_228),
.B(n_199),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_274),
.A2(n_278),
.B1(n_229),
.B2(n_265),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_262),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_272),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_270),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_257),
.A2(n_234),
.B1(n_249),
.B2(n_227),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_270),
.B1(n_290),
.B2(n_256),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_248),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_271),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_232),
.C(n_235),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_261),
.C(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_289),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_267),
.A2(n_238),
.B(n_245),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_295),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_274),
.B1(n_273),
.B2(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

XNOR2x1_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_256),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_300),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_305),
.Y(n_308)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_304),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_252),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_282),
.B(n_250),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_285),
.C(n_280),
.Y(n_310)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_310),
.A2(n_316),
.B1(n_301),
.B2(n_311),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_305),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_278),
.B(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_300),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_292),
.A2(n_281),
.B(n_293),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_319),
.B(n_295),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_276),
.B(n_250),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_296),
.Y(n_321)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_314),
.B(n_317),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_326),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_327),
.C(n_328),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_279),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_265),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_333),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_317),
.C(n_35),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_320),
.A2(n_12),
.B(n_14),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_325),
.B1(n_14),
.B2(n_6),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_328),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_336),
.A2(n_338),
.B(n_335),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_332),
.B(n_337),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_334),
.B(n_329),
.Y(n_341)
);

AOI322xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_338),
.A3(n_336),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_25),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_25),
.C(n_35),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_8),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_8),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_4),
.B(n_5),
.Y(n_346)
);


endmodule