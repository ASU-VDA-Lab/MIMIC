module real_jpeg_33214_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_0),
.Y(n_122)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_0),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_0),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_1),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_1),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_1),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_1),
.B(n_178),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_1),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_1),
.B(n_326),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_2),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_2),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_5),
.Y(n_129)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_5),
.Y(n_306)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_6),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_6),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_6),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_6),
.B(n_95),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_6),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_6),
.B(n_223),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_7),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_7),
.B(n_79),
.Y(n_188)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_7),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_8),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_8),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_128),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_8),
.B(n_116),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_8),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_8),
.B(n_77),
.Y(n_364)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_9),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_11),
.Y(n_322)
);

NAND2x1_ASAP7_75t_L g76 ( 
.A(n_12),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_12),
.B(n_35),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_12),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_12),
.B(n_269),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_SL g304 ( 
.A(n_12),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_12),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_13),
.B(n_143),
.Y(n_190)
);

NAND2x1_ASAP7_75t_L g361 ( 
.A(n_13),
.B(n_128),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_14),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_41),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_14),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_14),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_14),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_14),
.B(n_95),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_14),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_15),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_15),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_15),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_15),
.B(n_370),
.Y(n_369)
);

NAND2x1_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_16),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_16),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_16),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_16),
.B(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_16),
.B(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_16),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_16),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_17),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_17),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_17),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_17),
.B(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_347),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_240),
.B(n_345),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_162),
.B(n_213),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_22),
.B(n_162),
.C(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_110),
.C(n_138),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_23),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_71),
.B2(n_72),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_52),
.B2(n_53),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_26),
.Y(n_165)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XOR2x1_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_32),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_33),
.B(n_37),
.C(n_38),
.Y(n_199)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJx2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_44),
.C(n_49),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_39),
.A2(n_40),
.B1(n_49),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_42),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_44),
.B(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_50),
.Y(n_204)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_51),
.Y(n_275)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_53),
.B(n_71),
.C(n_165),
.Y(n_164)
);

XNOR2x1_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_55),
.A2(n_182),
.B(n_184),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_60),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_62),
.B(n_67),
.Y(n_184)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_63),
.B(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_65),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_67),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_87),
.C(n_98),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_73),
.B(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_84),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_76),
.B(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_78),
.A2(n_85),
.B(n_159),
.Y(n_158)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_82),
.A2(n_84),
.B(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_87),
.A2(n_98),
.B1(n_99),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_87),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_233)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_97),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_97),
.Y(n_328)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_106),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_100),
.A2(n_101),
.B1(n_106),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_104),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_105),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_106),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_110),
.B(n_139),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_124),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_111),
.B(n_114),
.Y(n_216)
);

OA21x2_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_120),
.B(n_123),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_120),
.Y(n_123)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_156),
.B1(n_157),
.B2(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_124),
.B(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_132),
.C(n_134),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_125),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_126),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_246)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_129),
.Y(n_254)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_129),
.Y(n_282)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_259)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_155),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_141),
.B(n_150),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_145),
.B1(n_146),
.B2(n_149),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_SL g206 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_388)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_161),
.C(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_160),
.B(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_164),
.B(n_351),
.C(n_352),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_197),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_167),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_180),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_169),
.B(n_181),
.C(n_196),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_171),
.B(n_174),
.C(n_177),
.Y(n_379)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_185),
.B1(n_195),
.B2(n_196),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_188),
.B(n_189),
.C(n_191),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_189),
.A2(n_190),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_194),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_197),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_211),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_209),
.B2(n_210),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_199),
.Y(n_355)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_205),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_202),
.B(n_205),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_202),
.B(n_205),
.Y(n_390)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_209),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_211),
.B(n_355),
.C(n_356),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_238),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_214),
.B(n_238),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.C(n_234),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_235),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.C(n_233),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_233),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.C(n_229),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_222),
.B(n_229),
.Y(n_294)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_225),
.B(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_228),
.Y(n_370)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_262),
.B(n_344),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_260),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g344 ( 
.A(n_242),
.B(n_260),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.C(n_258),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_243),
.B(n_342),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_245),
.B(n_258),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.C(n_251),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_247),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_248),
.B(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

AO22x1_ASAP7_75t_L g284 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_339),
.B(n_343),
.Y(n_262)
);

OAI21x1_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_296),
.B(n_338),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_285),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_265),
.B(n_285),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_278),
.C(n_284),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_266),
.A2(n_267),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_291),
.C(n_292),
.Y(n_290)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_278),
.A2(n_279),
.B1(n_284),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_283),
.Y(n_314)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_284),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_295),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_290),
.C(n_293),
.Y(n_340)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_331),
.B(n_337),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_315),
.B(n_330),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_307),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_299),
.B(n_307),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_304),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_304),
.Y(n_323)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_314),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_313),
.Y(n_308)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_313),
.C(n_314),
.Y(n_332)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_324),
.B(n_329),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_323),
.Y(n_329)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_341),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_391),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_353),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_375),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_365),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_361),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_373),
.Y(n_367)
);

XNOR2x1_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_387),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_389),
.B(n_390),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);


endmodule