module real_jpeg_18229_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_13),
.B1(n_19),
.B2(n_21),
.Y(n_18)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_1),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_2),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_2),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_2),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_3),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_3),
.A2(n_58),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_3),
.A2(n_58),
.B1(n_138),
.B2(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_3),
.A2(n_58),
.B1(n_335),
.B2(n_338),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_137),
.B1(n_138),
.B2(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_4),
.A2(n_137),
.B1(n_212),
.B2(n_217),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_5),
.A2(n_158),
.B1(n_161),
.B2(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_5),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_5),
.A2(n_164),
.B1(n_231),
.B2(n_235),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_6),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_6),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_6),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_7),
.A2(n_171),
.B1(n_174),
.B2(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_7),
.Y(n_177)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_8),
.Y(n_141)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_8),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_8),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_8),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_93),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_9),
.A2(n_104),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_9),
.A2(n_104),
.B1(n_363),
.B2(n_365),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_10),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_10),
.A2(n_131),
.B1(n_181),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_10),
.A2(n_131),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_12),
.A2(n_179),
.A3(n_182),
.B1(n_183),
.B2(n_188),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_12),
.B(n_28),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_12),
.B(n_65),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_12),
.B(n_135),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_12),
.B(n_352),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_12),
.A2(n_53),
.B1(n_98),
.B2(n_184),
.Y(n_371)
);

OAI32xp33_ASAP7_75t_L g373 ( 
.A1(n_12),
.A2(n_374),
.A3(n_377),
.B1(n_380),
.B2(n_381),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_15),
.Y(n_91)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_16),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_16),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_16),
.Y(n_216)
);

BUFx4f_ASAP7_75t_L g350 ( 
.A(n_16),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_258),
.B1(n_413),
.B2(n_414),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_22),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_257),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_221),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_24),
.B(n_221),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_145),
.C(n_194),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_25),
.B(n_409),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_62),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_26),
.B(n_63),
.C(n_108),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_48),
.B1(n_54),
.B2(n_61),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_27),
.Y(n_245)
);

OR2x6_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_28),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_32),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_34),
.Y(n_376)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_42),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_45),
.Y(n_192)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_51),
.A2(n_97),
.B1(n_102),
.B2(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_53),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_53),
.B(n_138),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_SL g279 ( 
.A1(n_53),
.A2(n_274),
.B(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_53),
.A2(n_149),
.B1(n_334),
.B2(n_341),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_53),
.B(n_265),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_54),
.Y(n_244)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_108),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_92),
.B1(n_103),
.B2(n_107),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_64),
.A2(n_92),
.B1(n_107),
.B2(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_64),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_64),
.A2(n_107),
.B1(n_196),
.B2(n_371),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_76),
.Y(n_64)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

AO22x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_74),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_112),
.B1(n_115),
.B2(n_117),
.Y(n_111)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_71),
.Y(n_234)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_83),
.B2(n_88),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_82),
.Y(n_200)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_91),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_91),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_97),
.B1(n_98),
.B2(n_102),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_97),
.A2(n_102),
.B1(n_311),
.B2(n_313),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_97),
.A2(n_102),
.B1(n_321),
.B2(n_325),
.Y(n_320)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_103),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_L g253 ( 
.A(n_107),
.B(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_127),
.B(n_134),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_109),
.A2(n_120),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_110),
.B(n_136),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_110),
.A2(n_135),
.B1(n_279),
.B2(n_284),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_110),
.A2(n_135),
.B1(n_284),
.B2(n_310),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_110),
.A2(n_403),
.B(n_404),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_121),
.B1(n_124),
.B2(n_126),
.Y(n_120)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_118),
.Y(n_286)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_119),
.Y(n_268)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_120),
.B(n_129),
.Y(n_404)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_122),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_124),
.Y(n_290)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_125),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_125),
.Y(n_326)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_125),
.Y(n_337)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_126),
.Y(n_276)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_133),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_135),
.B(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_145),
.A2(n_146),
.B1(n_194),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_178),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_147),
.B(n_178),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_157),
.B1(n_165),
.B2(n_170),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_148),
.A2(n_170),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_148),
.A2(n_319),
.B1(n_327),
.B2(n_328),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_148),
.A2(n_225),
.B(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_149),
.B(n_211),
.Y(n_210)
);

AOI21x1_ASAP7_75t_L g288 ( 
.A1(n_149),
.A2(n_289),
.B(n_296),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_149),
.A2(n_320),
.B1(n_334),
.B2(n_339),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_150),
.Y(n_338)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_152),
.Y(n_324)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_155),
.Y(n_300)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_156),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_206),
.B(n_210),
.Y(n_205)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_194),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_203),
.C(n_205),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_195),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_205),
.Y(n_399)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_209),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_215),
.Y(n_295)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_241),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_240),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_239),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_234),
.Y(n_379)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_256),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B(n_253),
.Y(n_250)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_258),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_407),
.B(n_412),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_393),
.B(n_406),
.Y(n_259)
);

OAI21x1_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_356),
.B(n_392),
.Y(n_260)
);

AOI21x1_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_316),
.B(n_355),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_287),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_263),
.B(n_287),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_277),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_264),
.A2(n_277),
.B1(n_278),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_269),
.A3(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_271),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_308),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_288),
.B(n_309),
.C(n_315),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_301),
.Y(n_391)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_315),
.Y(n_308)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_317),
.A2(n_331),
.B(n_354),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_329),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_329),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_344),
.B(n_353),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_343),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_343),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_351),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_357),
.B(n_358),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_372),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_370),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_370),
.C(n_372),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_362),
.Y(n_403)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_390),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_390),
.Y(n_401)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_SL g406 ( 
.A(n_394),
.B(n_395),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_400),
.B2(n_405),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_401),
.C(n_402),
.Y(n_411)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_400),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_411),
.Y(n_412)
);


endmodule