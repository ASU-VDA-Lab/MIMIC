module real_jpeg_27431_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_0),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_0),
.A2(n_55),
.B1(n_57),
.B2(n_168),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_168),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_168),
.Y(n_306)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_3),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_55),
.B1(n_57),
.B2(n_132),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_132),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_132),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_5),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_5),
.A2(n_31),
.B1(n_55),
.B2(n_57),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_6),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_6),
.A2(n_35),
.B1(n_55),
.B2(n_57),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_8),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_55),
.B1(n_57),
.B2(n_84),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_84),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_84),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_57),
.Y(n_56)
);

A2O1A1O1Ixp25_ASAP7_75t_L g60 ( 
.A1(n_9),
.A2(n_56),
.B(n_57),
.C(n_61),
.D(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_9),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_9),
.A2(n_81),
.B(n_85),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_25),
.B(n_118),
.C(n_119),
.D(n_122),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_9),
.B(n_25),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_9),
.A2(n_23),
.B(n_24),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_102),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_10),
.A2(n_55),
.B1(n_57),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_77),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_77),
.Y(n_201)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_12),
.A2(n_55),
.B1(n_57),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_66),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_178)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_55),
.B1(n_57),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_15),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_15),
.A2(n_55),
.B1(n_57),
.B2(n_151),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_151),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_151),
.Y(n_296)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_16),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_30),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_21),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_21),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_21),
.A2(n_26),
.B1(n_201),
.B2(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_21),
.A2(n_26),
.B1(n_34),
.B2(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_22),
.A2(n_28),
.B(n_102),
.C(n_171),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_24),
.A2(n_57),
.A3(n_118),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_26),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_26),
.B(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_26),
.Y(n_241)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_33),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_33),
.B(n_333),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_332),
.B(n_334),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_320),
.B(n_331),
.Y(n_39)
);

OAI321xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_284),
.A3(n_313),
.B1(n_318),
.B2(n_319),
.C(n_336),
.Y(n_40)
);

AOI321xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_234),
.A3(n_273),
.B1(n_278),
.B2(n_283),
.C(n_337),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_188),
.C(n_230),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_159),
.B(n_187),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_138),
.B(n_158),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_113),
.B(n_137),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_89),
.B(n_112),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_68),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_48),
.B(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_60),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_60),
.Y(n_98)
);

AOI32xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.A3(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_50),
.B(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_55),
.B(n_135),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_59),
.B(n_62),
.C(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_61),
.A2(n_63),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_61),
.A2(n_63),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_61),
.A2(n_63),
.B1(n_250),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_67),
.A2(n_78),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_67),
.A2(n_155),
.B1(n_186),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_67),
.A2(n_155),
.B1(n_209),
.B2(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_67),
.A2(n_155),
.B(n_259),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_80),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_75),
.C(n_80),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_72),
.A2(n_119),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_72),
.A2(n_119),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_72),
.A2(n_119),
.B1(n_262),
.B2(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_72),
.A2(n_119),
.B(n_325),
.Y(n_324)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B(n_85),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_87),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_81),
.A2(n_97),
.B1(n_131),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_81),
.A2(n_97),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_81),
.A2(n_97),
.B1(n_207),
.B2(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_81),
.A2(n_97),
.B(n_224),
.Y(n_252)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_102),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_88),
.A2(n_94),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_111),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_98),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_97),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_105),
.B(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_106),
.B(n_110),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_101),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_128),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_125),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_125),
.C(n_128),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_124),
.A2(n_144),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_124),
.A2(n_196),
.B1(n_221),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_124),
.A2(n_196),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_139),
.B(n_140),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_152),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_153),
.C(n_154),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_147),
.C(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_148),
.A2(n_200),
.B(n_202),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_148),
.A2(n_202),
.B(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_148),
.A2(n_241),
.B1(n_269),
.B2(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_148),
.A2(n_241),
.B1(n_296),
.B2(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_173),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_163),
.B(n_164),
.C(n_173),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_172),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_181),
.C(n_184),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_177),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_183),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_189),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_211),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_190),
.B(n_211),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_204),
.C(n_210),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_194),
.C(n_203),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_203),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_199),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_210),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_208),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_211)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_222),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_213),
.B(n_222),
.C(n_229),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_217),
.C(n_219),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_218),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_227),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_232),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_254),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_254),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_246),
.C(n_253),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_246),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_245),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_243),
.C(n_245),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_252),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_252),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_267),
.B(n_270),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_272),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_264),
.B1(n_265),
.B2(n_271),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_260),
.B(n_263),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_260),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_263),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_263),
.A2(n_286),
.B1(n_287),
.B2(n_298),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_271),
.C(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_270),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_274),
.A2(n_279),
.B(n_282),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_301),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_301),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_298),
.C(n_299),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_295),
.B2(n_297),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_290),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_294),
.C(n_295),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_291),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_292),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_294),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_305),
.C(n_309),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_295),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_297),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_304),
.C(n_312),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_299),
.A2(n_300),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_312),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_306),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_311),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_322),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_330),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_326),
.B1(n_328),
.B2(n_329),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_324),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_326),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_329),
.C(n_330),
.Y(n_333)
);


endmodule