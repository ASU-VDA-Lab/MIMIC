module fake_jpeg_8182_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_SL g23 ( 
.A(n_18),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_12),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_1),
.C(n_3),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_11),
.B(n_18),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_28),
.A2(n_30),
.B(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_35),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_SL g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_41),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_18),
.B(n_19),
.C(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_19),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_20),
.B1(n_17),
.B2(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_38),
.B1(n_47),
.B2(n_40),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_20),
.B1(n_32),
.B2(n_34),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_33),
.B1(n_37),
.B2(n_25),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_60),
.Y(n_66)
);

OAI322xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_54),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_8),
.C2(n_9),
.Y(n_65)
);

NOR2x1p5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_55),
.C(n_51),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_15),
.B(n_13),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_55),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_14),
.C(n_59),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_59),
.B1(n_60),
.B2(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_8),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_15),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_71),
.B(n_69),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_72),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_70),
.A3(n_9),
.B1(n_6),
.B2(n_4),
.C(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_6),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_75),
.Y(n_79)
);


endmodule