module fake_jpeg_1194_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NAND2x1_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_60),
.Y(n_63)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_42),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_51),
.B1(n_49),
.B2(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_55),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_82),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_70),
.A2(n_59),
.B1(n_51),
.B2(n_41),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_47),
.B1(n_45),
.B2(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_22),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_44),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_84),
.B(n_82),
.Y(n_104)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_87),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_91),
.B1(n_17),
.B2(n_18),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_27),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_5),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_101),
.B1(n_81),
.B2(n_10),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_108),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_110),
.Y(n_126)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_26),
.Y(n_112)
);

OAI321xp33_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_117),
.A3(n_108),
.B1(n_102),
.B2(n_38),
.C(n_37),
.Y(n_125)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_118),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_96),
.B(n_10),
.Y(n_115)
);

XNOR2x1_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_117),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_14),
.C(n_15),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_36),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_16),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_101),
.B(n_24),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_124),
.C(n_129),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_21),
.B(n_28),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_32),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_128),
.B(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

AOI221xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_127),
.B1(n_119),
.B2(n_120),
.C(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_140),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_137),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_141),
.B(n_134),
.CI(n_131),
.CON(n_143),
.SN(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_131),
.C(n_138),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_142),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_142),
.B(n_143),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_148),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_132),
.Y(n_150)
);


endmodule