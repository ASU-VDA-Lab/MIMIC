module fake_ariane_675_n_1679 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1679);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1679;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_89),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_25),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_24),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_83),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_42),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_103),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_20),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_70),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_51),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_0),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_17),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_10),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_51),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_30),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_9),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_48),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_87),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_7),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_44),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_39),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_134),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_132),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_40),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_6),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_33),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_142),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_66),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_21),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_28),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_41),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_58),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_104),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_31),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_49),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_80),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_39),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_47),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_82),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_67),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_22),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_21),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_85),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_147),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_78),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_36),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_35),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_13),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_10),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_92),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_49),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_41),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_2),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_56),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_28),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_18),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_128),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_56),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_9),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_109),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_43),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_117),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_58),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_118),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_71),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_138),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_68),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_16),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_55),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_46),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_79),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_47),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_55),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_14),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_12),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_27),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_24),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_11),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_52),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_40),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_44),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_29),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_111),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_1),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_23),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_20),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_84),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_112),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_29),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_37),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_19),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_110),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_43),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_62),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_26),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_101),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_12),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_94),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_42),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_17),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_130),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_76),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_2),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_135),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_143),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_97),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_119),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_81),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_144),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_120),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_1),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_15),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_5),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_152),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_60),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_33),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_116),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_121),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_61),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_139),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_149),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_4),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_15),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_90),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_50),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_22),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_46),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_140),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_158),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_153),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_153),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_3),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_191),
.B(n_3),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_167),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_165),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_197),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_236),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_227),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_227),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_166),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_199),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_R g320 ( 
.A(n_288),
.B(n_303),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_200),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_166),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_169),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_169),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_171),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_172),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_171),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_160),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_174),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_164),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_207),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_174),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_191),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_179),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_168),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_179),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_170),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_186),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_261),
.B(n_4),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_186),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_187),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_173),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_172),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_192),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_221),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_172),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_175),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_225),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_194),
.B(n_5),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_176),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_194),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_195),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_180),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_195),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_209),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_294),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_294),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_202),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_181),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_183),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_209),
.B(n_6),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_184),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_210),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_190),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_193),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_204),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_204),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_294),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_201),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_205),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_211),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_216),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_204),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_210),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_294),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_217),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_223),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_305),
.B(n_177),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_306),
.B(n_223),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_306),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_318),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_319),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_312),
.B(n_223),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_312),
.B(n_234),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_326),
.B(n_234),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_322),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_323),
.B(n_238),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_315),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_324),
.B(n_325),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_325),
.B(n_238),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_358),
.B(n_225),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_350),
.A2(n_202),
.B1(n_301),
.B2(n_300),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_358),
.B(n_359),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_321),
.A2(n_302),
.B1(n_196),
.B2(n_208),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_329),
.B(n_239),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_344),
.B(n_375),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_344),
.B(n_263),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_330),
.B(n_239),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_329),
.Y(n_419)
);

BUFx8_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_332),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_371),
.B(n_256),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_334),
.Y(n_425)
);

BUFx8_ASAP7_75t_L g426 ( 
.A(n_379),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_336),
.B(n_263),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_336),
.B(n_155),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_359),
.B(n_256),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_341),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_341),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_342),
.B(n_260),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_345),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_379),
.B(n_346),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_316),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_328),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_350),
.A2(n_219),
.B1(n_298),
.B2(n_297),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_354),
.B(n_155),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_354),
.B(n_263),
.Y(n_448)
);

CKINVDCx6p67_ASAP7_75t_R g449 ( 
.A(n_386),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_404),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

BUFx4f_ASAP7_75t_L g453 ( 
.A(n_392),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_432),
.B(n_377),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_SL g456 ( 
.A(n_445),
.B(n_307),
.Y(n_456)
);

OAI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_381),
.A2(n_307),
.B(n_304),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_392),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_392),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_416),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_433),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

NAND3xp33_ASAP7_75t_L g468 ( 
.A(n_397),
.B(n_363),
.C(n_351),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_433),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_404),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_443),
.Y(n_473)
);

INVxp67_ASAP7_75t_R g474 ( 
.A(n_445),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_377),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_443),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_443),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_389),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_418),
.B(n_335),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_443),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_393),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_423),
.B(n_337),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_412),
.A2(n_339),
.B1(n_308),
.B2(n_304),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_446),
.B(n_343),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_393),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_446),
.B(n_349),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_393),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_393),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_414),
.B(n_308),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_410),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_409),
.B(n_352),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_401),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_L g498 ( 
.A(n_401),
.B(n_252),
.C(n_156),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_416),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_387),
.Y(n_500)
);

AND3x2_ASAP7_75t_L g501 ( 
.A(n_389),
.B(n_360),
.C(n_333),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_419),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_410),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_429),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_419),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_419),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_441),
.B(n_348),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_416),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_420),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_429),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_434),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_434),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_396),
.B(n_320),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_405),
.B(n_355),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_405),
.B(n_361),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_396),
.B(n_368),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_441),
.B(n_369),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_413),
.B(n_364),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_384),
.B(n_356),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_412),
.B(n_373),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_429),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_417),
.B(n_367),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_381),
.B(n_372),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_421),
.B(n_374),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_421),
.B(n_356),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_SL g531 ( 
.A(n_407),
.B(n_378),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_397),
.A2(n_376),
.B1(n_365),
.B2(n_357),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_387),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_387),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_421),
.B(n_370),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_395),
.A2(n_333),
.B1(n_360),
.B2(n_262),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_439),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_414),
.B(n_309),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_387),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_442),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_383),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_380),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_437),
.B(n_357),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_391),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_391),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_437),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_384),
.B(n_365),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_383),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_437),
.B(n_376),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_385),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_428),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_385),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_417),
.Y(n_560)
);

AND3x1_ASAP7_75t_L g561 ( 
.A(n_417),
.B(n_185),
.C(n_158),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_398),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_398),
.B(n_311),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_407),
.A2(n_250),
.B1(n_244),
.B2(n_241),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_399),
.B(n_313),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_399),
.B(n_260),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_384),
.B(n_225),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_428),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_420),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_384),
.B(n_225),
.Y(n_570)
);

BUFx4f_ASAP7_75t_L g571 ( 
.A(n_428),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_400),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_400),
.B(n_267),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_382),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_382),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_402),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_402),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_382),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_388),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_406),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_388),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_406),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_384),
.B(n_247),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_388),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_428),
.Y(n_585)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_394),
.Y(n_586)
);

INVxp67_ASAP7_75t_SL g587 ( 
.A(n_420),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_380),
.Y(n_588)
);

AO22x2_ASAP7_75t_L g589 ( 
.A1(n_420),
.A2(n_185),
.B1(n_196),
.B2(n_302),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_411),
.B(n_267),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_390),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_411),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_422),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_394),
.B(n_247),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_422),
.B(n_272),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_424),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_390),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_497),
.B(n_424),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_480),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_577),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_492),
.B(n_425),
.Y(n_601)
);

NAND2x1_ASAP7_75t_L g602 ( 
.A(n_558),
.B(n_425),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_503),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_497),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_450),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_480),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_483),
.B(n_430),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_492),
.B(n_430),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_507),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_528),
.B(n_420),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_577),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_577),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_524),
.B(n_431),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_524),
.B(n_431),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_524),
.B(n_435),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_468),
.A2(n_586),
.B1(n_488),
.B2(n_554),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_454),
.B(n_457),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_524),
.B(n_435),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_520),
.B(n_440),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_507),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_508),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_554),
.B(n_394),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_560),
.B(n_440),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_560),
.B(n_394),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_494),
.A2(n_426),
.B1(n_394),
.B2(n_427),
.Y(n_625)
);

OAI221xp5_ASAP7_75t_L g626 ( 
.A1(n_488),
.A2(n_257),
.B1(n_259),
.B2(n_246),
.C(n_255),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_547),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_509),
.B(n_522),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_508),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_492),
.B(n_426),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_513),
.Y(n_631)
);

BUFx8_ASAP7_75t_L g632 ( 
.A(n_450),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_492),
.B(n_426),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_555),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_481),
.B(n_331),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_513),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_557),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_494),
.A2(n_436),
.B1(n_415),
.B2(n_408),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_506),
.B(n_426),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_514),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_514),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_506),
.B(n_426),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_476),
.B(n_517),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_466),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_509),
.B(n_427),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_509),
.B(n_427),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_506),
.B(n_395),
.Y(n_647)
);

A2O1A1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_457),
.A2(n_436),
.B(n_415),
.C(n_408),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_L g649 ( 
.A(n_466),
.B(n_428),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_516),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_516),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_494),
.A2(n_448),
.B1(n_427),
.B2(n_428),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_509),
.B(n_522),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_588),
.A2(n_403),
.B(n_390),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_557),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_559),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_489),
.B(n_491),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_559),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_468),
.A2(n_403),
.B1(n_224),
.B2(n_291),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_487),
.B(n_427),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_586),
.B(n_448),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_522),
.B(n_448),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_522),
.B(n_448),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_506),
.B(n_448),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_586),
.A2(n_232),
.B1(n_230),
.B2(n_226),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_494),
.A2(n_447),
.B1(n_428),
.B2(n_247),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_490),
.B(n_428),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_490),
.B(n_428),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_518),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_482),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_476),
.A2(n_447),
.B1(n_272),
.B2(n_296),
.Y(n_671)
);

AND2x2_ASAP7_75t_SL g672 ( 
.A(n_569),
.B(n_561),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_490),
.B(n_502),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_562),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_502),
.B(n_447),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_466),
.Y(n_676)
);

OAI221xp5_ASAP7_75t_L g677 ( 
.A1(n_494),
.A2(n_208),
.B1(n_229),
.B2(n_222),
.C(n_218),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_482),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_519),
.A2(n_456),
.B1(n_554),
.B2(n_586),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_569),
.B(n_235),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_527),
.B(n_248),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_471),
.B(n_229),
.C(n_222),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_502),
.B(n_533),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_554),
.A2(n_447),
.B1(n_296),
.B2(n_293),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_518),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_558),
.B(n_281),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_532),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_532),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_563),
.Y(n_689)
);

BUFx6f_ASAP7_75t_SL g690 ( 
.A(n_461),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_562),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_572),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_572),
.B(n_576),
.Y(n_693)
);

AO22x1_ASAP7_75t_L g694 ( 
.A1(n_587),
.A2(n_273),
.B1(n_254),
.B2(n_258),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_449),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_474),
.B(n_347),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_545),
.Y(n_697)
);

INVxp67_ASAP7_75t_SL g698 ( 
.A(n_480),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_449),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_474),
.B(n_247),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_576),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_558),
.B(n_281),
.Y(n_702)
);

OAI221xp5_ASAP7_75t_L g703 ( 
.A1(n_561),
.A2(n_255),
.B1(n_212),
.B2(n_266),
.C(n_218),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_554),
.A2(n_268),
.B1(n_249),
.B2(n_271),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_580),
.B(n_447),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_565),
.B(n_286),
.C(n_285),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_L g708 ( 
.A1(n_525),
.A2(n_235),
.B1(n_240),
.B2(n_212),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_484),
.B(n_233),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_496),
.A2(n_531),
.B1(n_499),
.B2(n_510),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_558),
.B(n_282),
.Y(n_711)
);

BUFx5_ASAP7_75t_L g712 ( 
.A(n_486),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_527),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_589),
.A2(n_447),
.B1(n_277),
.B2(n_240),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_501),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_466),
.B(n_447),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_461),
.B(n_233),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_466),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_582),
.B(n_447),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_545),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_582),
.B(n_447),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_592),
.B(n_282),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_499),
.B(n_274),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_546),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_592),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_593),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_546),
.Y(n_727)
);

OAI21xp33_ASAP7_75t_L g728 ( 
.A1(n_510),
.A2(n_287),
.B(n_242),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_541),
.Y(n_729)
);

NOR2x1p5_ASAP7_75t_L g730 ( 
.A(n_525),
.B(n_242),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_523),
.B(n_290),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_500),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_593),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_596),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_568),
.B(n_290),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_536),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_596),
.A2(n_246),
.B1(n_245),
.B2(n_253),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_568),
.B(n_293),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_530),
.B(n_245),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_556),
.B(n_253),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_568),
.B(n_161),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_515),
.B(n_257),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_511),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_536),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_538),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_589),
.A2(n_277),
.B1(n_266),
.B2(n_259),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_529),
.B(n_567),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_486),
.B(n_154),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_493),
.B(n_157),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_537),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_SL g751 ( 
.A(n_553),
.B(n_277),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_493),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_568),
.B(n_161),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_538),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_540),
.Y(n_755)
);

BUFx8_ASAP7_75t_L g756 ( 
.A(n_495),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_504),
.B(n_505),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_539),
.A2(n_277),
.B1(n_228),
.B2(n_251),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_504),
.B(n_159),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_541),
.B(n_498),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_585),
.B(n_220),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_585),
.B(n_220),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_512),
.B(n_162),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_512),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_478),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_638),
.B(n_478),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_607),
.B(n_550),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_643),
.B(n_553),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_689),
.B(n_570),
.Y(n_769)
);

BUFx4f_ASAP7_75t_L g770 ( 
.A(n_604),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_616),
.A2(n_553),
.B1(n_521),
.B2(n_526),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_622),
.B(n_583),
.Y(n_772)
);

OAI21xp33_ASAP7_75t_L g773 ( 
.A1(n_681),
.A2(n_564),
.B(n_526),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_628),
.B(n_553),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_679),
.B(n_478),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_635),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_647),
.A2(n_534),
.B(n_500),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_617),
.A2(n_521),
.B(n_544),
.C(n_542),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_599),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_647),
.A2(n_534),
.B(n_500),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_617),
.A2(n_610),
.B1(n_672),
.B2(n_657),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_648),
.A2(n_455),
.B(n_452),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_713),
.B(n_594),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_693),
.A2(n_534),
.B(n_500),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_SL g785 ( 
.A(n_695),
.B(n_585),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_627),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_601),
.A2(n_534),
.B(n_453),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_601),
.A2(n_453),
.B(n_535),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_608),
.A2(n_453),
.B(n_535),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_653),
.B(n_540),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_712),
.B(n_478),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_SL g792 ( 
.A(n_699),
.B(n_585),
.Y(n_792)
);

OAI21xp33_ASAP7_75t_L g793 ( 
.A1(n_681),
.A2(n_595),
.B(n_590),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_673),
.A2(n_543),
.B(n_455),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_757),
.A2(n_543),
.B(n_458),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_610),
.A2(n_589),
.B1(n_544),
.B2(n_542),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_732),
.A2(n_458),
.B(n_473),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_672),
.A2(n_589),
.B1(n_462),
.B2(n_463),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_664),
.A2(n_452),
.B(n_467),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_743),
.B(n_571),
.Y(n_800)
);

OAI21xp33_ASAP7_75t_SL g801 ( 
.A1(n_664),
.A2(n_566),
.B(n_573),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_660),
.A2(n_462),
.B(n_571),
.C(n_463),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_657),
.A2(n_462),
.B1(n_463),
.B2(n_467),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_712),
.B(n_478),
.Y(n_804)
);

AOI21x1_ASAP7_75t_L g805 ( 
.A1(n_741),
.A2(n_477),
.B(n_475),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_632),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_731),
.B(n_462),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_619),
.A2(n_477),
.B(n_475),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_634),
.Y(n_809)
);

AOI21x1_ASAP7_75t_L g810 ( 
.A1(n_741),
.A2(n_469),
.B(n_473),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_645),
.B(n_548),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_606),
.A2(n_469),
.B(n_459),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_698),
.A2(n_451),
.B(n_459),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_603),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_644),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_646),
.B(n_548),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_678),
.B(n_451),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_609),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_667),
.A2(n_460),
.B(n_465),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_696),
.B(n_571),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_712),
.B(n_460),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_750),
.B(n_548),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_609),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_662),
.B(n_551),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_660),
.B(n_747),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_712),
.B(n_465),
.Y(n_826)
);

NOR2x2_ASAP7_75t_L g827 ( 
.A(n_680),
.B(n_470),
.Y(n_827)
);

NOR2x1_ASAP7_75t_L g828 ( 
.A(n_680),
.B(n_551),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_747),
.B(n_551),
.Y(n_829)
);

INVx11_ASAP7_75t_L g830 ( 
.A(n_632),
.Y(n_830)
);

BUFx8_ASAP7_75t_L g831 ( 
.A(n_690),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_663),
.B(n_470),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_661),
.B(n_472),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_668),
.A2(n_472),
.B(n_479),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_605),
.B(n_552),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_661),
.B(n_479),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_659),
.A2(n_703),
.B(n_648),
.C(n_624),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_706),
.A2(n_485),
.B(n_588),
.Y(n_838)
);

AND2x6_ASAP7_75t_L g839 ( 
.A(n_622),
.B(n_485),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_637),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_670),
.B(n_552),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_746),
.A2(n_277),
.B1(n_597),
.B2(n_578),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_742),
.B(n_574),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_675),
.A2(n_588),
.B(n_591),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_SL g845 ( 
.A(n_632),
.B(n_163),
.Y(n_845)
);

OAI21xp33_ASAP7_75t_L g846 ( 
.A1(n_723),
.A2(n_588),
.B(n_251),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_730),
.B(n_700),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_613),
.B(n_574),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_655),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_614),
.B(n_575),
.Y(n_850)
);

AO21x1_ASAP7_75t_L g851 ( 
.A1(n_630),
.A2(n_228),
.B(n_289),
.Y(n_851)
);

NOR2x1_ASAP7_75t_L g852 ( 
.A(n_680),
.B(n_575),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_620),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_602),
.A2(n_597),
.B(n_591),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_615),
.B(n_578),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_644),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_618),
.A2(n_581),
.B(n_579),
.C(n_584),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_752),
.A2(n_584),
.B(n_581),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_599),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_622),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_644),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_710),
.B(n_579),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_623),
.B(n_464),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_756),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_712),
.B(n_464),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_683),
.A2(n_289),
.B(n_8),
.C(n_11),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_723),
.B(n_464),
.Y(n_867)
);

O2A1O1Ixp5_ASAP7_75t_L g868 ( 
.A1(n_722),
.A2(n_549),
.B(n_464),
.C(n_380),
.Y(n_868)
);

O2A1O1Ixp5_ASAP7_75t_L g869 ( 
.A1(n_656),
.A2(n_549),
.B(n_464),
.C(n_380),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_598),
.A2(n_269),
.B1(n_182),
.B2(n_299),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_719),
.A2(n_549),
.B(n_265),
.Y(n_871)
);

BUFx2_ASAP7_75t_SL g872 ( 
.A(n_690),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_764),
.A2(n_744),
.B(n_736),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_620),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_626),
.A2(n_243),
.B1(n_295),
.B2(n_292),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_658),
.A2(n_726),
.B(n_725),
.C(n_733),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_712),
.B(n_380),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_744),
.A2(n_231),
.B(n_284),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_644),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_712),
.B(n_380),
.Y(n_880)
);

AO21x1_ASAP7_75t_L g881 ( 
.A1(n_630),
.A2(n_95),
.B(n_146),
.Y(n_881)
);

AO21x1_ASAP7_75t_L g882 ( 
.A1(n_633),
.A2(n_93),
.B(n_145),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_676),
.B(n_283),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_721),
.A2(n_654),
.B(n_745),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_677),
.A2(n_7),
.B(n_8),
.C(n_13),
.Y(n_885)
);

O2A1O1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_674),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_886)
);

BUFx4f_ASAP7_75t_L g887 ( 
.A(n_715),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_745),
.A2(n_280),
.B(n_279),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_691),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_754),
.A2(n_278),
.B(n_276),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_625),
.B(n_206),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_692),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_701),
.B(n_275),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_754),
.A2(n_270),
.B(n_237),
.Y(n_894)
);

AOI21xp33_ASAP7_75t_L g895 ( 
.A1(n_708),
.A2(n_215),
.B(n_214),
.Y(n_895)
);

BUFx12f_ASAP7_75t_L g896 ( 
.A(n_756),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_705),
.A2(n_213),
.B1(n_203),
.B2(n_198),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_734),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_717),
.B(n_652),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_694),
.B(n_189),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_682),
.A2(n_23),
.B(n_25),
.C(n_26),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_707),
.B(n_188),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_755),
.A2(n_178),
.B(n_65),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_709),
.B(n_27),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_714),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_755),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_906)
);

NOR2xp67_ASAP7_75t_L g907 ( 
.A(n_760),
.B(n_86),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_748),
.A2(n_73),
.B(n_133),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_739),
.B(n_740),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_621),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_600),
.B(n_34),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_749),
.A2(n_91),
.B(n_129),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_676),
.B(n_37),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_729),
.B(n_704),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_611),
.A2(n_72),
.B(n_127),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_612),
.A2(n_63),
.B(n_126),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_633),
.B(n_38),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_671),
.B(n_38),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_676),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_676),
.B(n_45),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_759),
.A2(n_96),
.B(n_123),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_665),
.A2(n_45),
.B(n_48),
.C(n_50),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_763),
.A2(n_105),
.B(n_122),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_753),
.A2(n_59),
.B(n_115),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_728),
.B(n_52),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_737),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_629),
.B(n_53),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_629),
.B(n_53),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_686),
.B(n_54),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_666),
.B(n_54),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_753),
.A2(n_761),
.B(n_762),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_765),
.A2(n_57),
.B1(n_108),
.B2(n_114),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_631),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_761),
.A2(n_136),
.B(n_57),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_684),
.B(n_631),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_636),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_762),
.A2(n_738),
.B(n_735),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_686),
.B(n_702),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_718),
.B(n_765),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_L g940 ( 
.A(n_702),
.B(n_711),
.C(n_738),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_758),
.A2(n_639),
.B(n_642),
.C(n_735),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_640),
.B(n_697),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_640),
.A2(n_688),
.B(n_641),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_641),
.A2(n_697),
.B(n_727),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_825),
.A2(n_639),
.B1(n_642),
.B2(n_765),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_786),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_825),
.A2(n_711),
.B(n_649),
.C(n_716),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_905),
.A2(n_650),
.B1(n_651),
.B2(n_669),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_817),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_781),
.A2(n_718),
.B1(n_765),
.B2(n_669),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_831),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_769),
.A2(n_650),
.B(n_651),
.C(n_685),
.Y(n_952)
);

CKINVDCx8_ASAP7_75t_R g953 ( 
.A(n_872),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_SL g954 ( 
.A1(n_926),
.A2(n_718),
.B1(n_687),
.B2(n_688),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_877),
.A2(n_880),
.B(n_804),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_SL g956 ( 
.A1(n_905),
.A2(n_718),
.B1(n_687),
.B2(n_685),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_860),
.B(n_720),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_909),
.B(n_720),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_769),
.B(n_724),
.Y(n_959)
);

CKINVDCx16_ASAP7_75t_R g960 ( 
.A(n_845),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_809),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_837),
.A2(n_724),
.B(n_727),
.C(n_751),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_831),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_776),
.B(n_847),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_SL g965 ( 
.A1(n_783),
.A2(n_806),
.B1(n_864),
.B2(n_906),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_835),
.B(n_783),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_830),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_829),
.B(n_917),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_814),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_770),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_818),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_SL g972 ( 
.A1(n_791),
.A2(n_804),
.B(n_865),
.C(n_880),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_929),
.Y(n_973)
);

CKINVDCx10_ASAP7_75t_R g974 ( 
.A(n_896),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_860),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_835),
.B(n_841),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_823),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_877),
.A2(n_791),
.B(n_867),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_853),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_772),
.B(n_828),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_766),
.A2(n_784),
.B(n_829),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_815),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_766),
.A2(n_826),
.B(n_821),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_874),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_827),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_930),
.A2(n_929),
.B1(n_899),
.B2(n_914),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_770),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_821),
.A2(n_826),
.B(n_793),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_900),
.B(n_822),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_772),
.A2(n_800),
.B1(n_875),
.B2(n_820),
.Y(n_990)
);

AND2x6_ASAP7_75t_L g991 ( 
.A(n_917),
.B(n_798),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_840),
.B(n_849),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_822),
.B(n_768),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_910),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_887),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_889),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_839),
.Y(n_997)
);

AO21x1_ASAP7_75t_L g998 ( 
.A1(n_775),
.A2(n_941),
.B(n_916),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_938),
.B(n_801),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_767),
.B(n_773),
.Y(n_1000)
);

OAI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_904),
.A2(n_906),
.B(n_918),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_892),
.B(n_790),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_938),
.B(n_774),
.Y(n_1003)
);

INVx6_ASAP7_75t_L g1004 ( 
.A(n_898),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_876),
.B(n_935),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_785),
.B(n_887),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_839),
.B(n_792),
.Y(n_1007)
);

NAND2x1_ASAP7_75t_L g1008 ( 
.A(n_861),
.B(n_919),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_873),
.A2(n_777),
.B(n_780),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_839),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_815),
.B(n_856),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_SL g1012 ( 
.A(n_901),
.B(n_886),
.C(n_902),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_L g1013 ( 
.A(n_922),
.B(n_885),
.C(n_866),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_839),
.Y(n_1014)
);

OA21x2_ASAP7_75t_L g1015 ( 
.A1(n_884),
.A2(n_782),
.B(n_778),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_913),
.A2(n_920),
.B(n_893),
.C(n_925),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_844),
.A2(n_865),
.B(n_794),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_796),
.B(n_940),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_862),
.B(n_833),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_862),
.B(n_907),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_863),
.A2(n_795),
.B(n_787),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_836),
.B(n_811),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_815),
.Y(n_1023)
);

O2A1O1Ixp5_ASAP7_75t_L g1024 ( 
.A1(n_913),
.A2(n_920),
.B(n_868),
.C(n_934),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_928),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_779),
.B(n_859),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_779),
.B(n_859),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_815),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_937),
.A2(n_846),
.B(n_915),
.C(n_931),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_775),
.A2(n_911),
.B(n_803),
.C(n_927),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_816),
.B(n_824),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_933),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_856),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_856),
.B(n_879),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_857),
.A2(n_802),
.B(n_799),
.C(n_869),
.Y(n_1035)
);

OR2x6_ASAP7_75t_L g1036 ( 
.A(n_852),
.B(n_891),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_936),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_771),
.A2(n_897),
.B(n_895),
.C(n_883),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_843),
.B(n_832),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_883),
.A2(n_807),
.B(n_890),
.C(n_888),
.Y(n_1040)
);

OAI22x1_ASAP7_75t_L g1041 ( 
.A1(n_870),
.A2(n_939),
.B1(n_861),
.B2(n_919),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_942),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_788),
.A2(n_789),
.B(n_819),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_856),
.B(n_879),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_848),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_834),
.A2(n_808),
.B(n_812),
.Y(n_1046)
);

BUFx8_ASAP7_75t_SL g1047 ( 
.A(n_879),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_850),
.B(n_855),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_879),
.B(n_939),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_943),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_881),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_878),
.A2(n_894),
.B(n_932),
.C(n_838),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_944),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_858),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_805),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_871),
.B(n_842),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_842),
.B(n_797),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_L g1058 ( 
.A(n_908),
.B(n_912),
.C(n_923),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_810),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_813),
.B(n_854),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_851),
.B(n_903),
.Y(n_1061)
);

INVx8_ASAP7_75t_L g1062 ( 
.A(n_882),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_869),
.A2(n_868),
.B(n_921),
.C(n_924),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_SL g1064 ( 
.A1(n_845),
.A2(n_414),
.B1(n_589),
.B2(n_511),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_825),
.B(n_643),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_825),
.A2(n_689),
.B1(n_483),
.B2(n_481),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_860),
.Y(n_1067)
);

NOR2xp67_ASAP7_75t_SL g1068 ( 
.A(n_872),
.B(n_450),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_825),
.A2(n_483),
.B(n_689),
.C(n_487),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_825),
.B(n_643),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_896),
.B(n_386),
.Y(n_1071)
);

NAND3xp33_ASAP7_75t_SL g1072 ( 
.A(n_781),
.B(n_483),
.C(n_689),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_831),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_825),
.B(n_689),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_825),
.B(n_781),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_825),
.A2(n_689),
.B1(n_483),
.B2(n_481),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_770),
.B(n_604),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_825),
.B(n_643),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_776),
.B(n_476),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_825),
.B(n_781),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_946),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1082)
);

INVxp67_ASAP7_75t_SL g1083 ( 
.A(n_1019),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_1069),
.A2(n_973),
.B(n_1018),
.C(n_1019),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_998),
.A2(n_1055),
.A3(n_1029),
.B(n_1061),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_L g1086 ( 
.A(n_1072),
.B(n_1074),
.C(n_973),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1018),
.A2(n_1001),
.B(n_1038),
.C(n_1080),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1066),
.A2(n_1076),
.B1(n_1074),
.B2(n_1072),
.Y(n_1088)
);

AOI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1017),
.A2(n_1043),
.B(n_1020),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_999),
.A2(n_1080),
.B(n_1075),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1021),
.A2(n_1046),
.B(n_1009),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1065),
.B(n_1070),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_1030),
.A2(n_1041),
.A3(n_1035),
.B(n_983),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1003),
.B(n_1075),
.Y(n_1094)
);

AO31x2_ASAP7_75t_L g1095 ( 
.A1(n_978),
.A2(n_1050),
.A3(n_1053),
.B(n_988),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_1024),
.A2(n_1060),
.B(n_955),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1003),
.B(n_1078),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_SL g1098 ( 
.A(n_960),
.B(n_991),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1048),
.B(n_1045),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1014),
.B(n_995),
.Y(n_1100)
);

CKINVDCx8_ASAP7_75t_R g1101 ( 
.A(n_974),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1079),
.B(n_964),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1048),
.B(n_966),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_L g1104 ( 
.A(n_1000),
.B(n_1013),
.C(n_1012),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_SL g1105 ( 
.A1(n_1016),
.A2(n_1005),
.B(n_959),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_961),
.Y(n_1106)
);

AOI221x1_ASAP7_75t_L g1107 ( 
.A1(n_1000),
.A2(n_956),
.B1(n_954),
.B2(n_945),
.C(n_965),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1054),
.A2(n_1024),
.B(n_1052),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_993),
.B(n_1022),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1058),
.A2(n_1049),
.B(n_1040),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1022),
.A2(n_993),
.B(n_972),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_987),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_997),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1002),
.B(n_986),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_986),
.B(n_1039),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_L g1116 ( 
.A(n_1012),
.B(n_968),
.C(n_947),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_967),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_SL g1118 ( 
.A1(n_968),
.A2(n_1008),
.B(n_1011),
.C(n_1034),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_1049),
.A2(n_1011),
.B(n_1034),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_962),
.A2(n_1031),
.A3(n_1057),
.B(n_1042),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1031),
.A2(n_1056),
.B(n_958),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_1044),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_952),
.A2(n_950),
.B(n_1015),
.Y(n_1123)
);

OA21x2_ASAP7_75t_L g1124 ( 
.A1(n_948),
.A2(n_1037),
.B(n_989),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1015),
.A2(n_1062),
.B(n_992),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1062),
.A2(n_1026),
.B(n_1027),
.Y(n_1126)
);

OAI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1071),
.A2(n_976),
.B1(n_990),
.B2(n_1025),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1007),
.A2(n_997),
.B(n_948),
.Y(n_1128)
);

AO32x2_ASAP7_75t_L g1129 ( 
.A1(n_1064),
.A2(n_991),
.A3(n_949),
.B1(n_1062),
.B2(n_1059),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1064),
.A2(n_991),
.B1(n_980),
.B2(n_1068),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_996),
.A2(n_957),
.B(n_1010),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_980),
.B(n_967),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_957),
.A2(n_1051),
.B(n_1044),
.Y(n_1133)
);

AOI221xp5_ASAP7_75t_L g1134 ( 
.A1(n_1077),
.A2(n_970),
.B1(n_949),
.B2(n_963),
.C(n_951),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_975),
.A2(n_1067),
.B1(n_1023),
.B2(n_1028),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1006),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_969),
.A2(n_971),
.B(n_994),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_975),
.B(n_1067),
.Y(n_1138)
);

BUFx4_ASAP7_75t_SL g1139 ( 
.A(n_1073),
.Y(n_1139)
);

AOI221x1_ASAP7_75t_L g1140 ( 
.A1(n_1059),
.A2(n_977),
.B1(n_979),
.B2(n_984),
.C(n_982),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1036),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1059),
.A2(n_991),
.A3(n_1036),
.B(n_1044),
.Y(n_1142)
);

AOI221xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1059),
.A2(n_982),
.B1(n_1033),
.B2(n_985),
.C(n_991),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_982),
.A2(n_1033),
.B(n_1036),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_982),
.A2(n_1033),
.B(n_1004),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1006),
.A2(n_689),
.B1(n_1074),
.B2(n_483),
.C(n_1072),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1004),
.A2(n_689),
.B(n_483),
.C(n_1072),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_953),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_SL g1149 ( 
.A1(n_1075),
.A2(n_1080),
.B(n_1072),
.C(n_1065),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_966),
.B(n_825),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1074),
.B(n_1066),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_946),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_998),
.A2(n_1055),
.A3(n_851),
.B(n_1029),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1017),
.A2(n_1043),
.B(n_1021),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_1075),
.A2(n_1080),
.B(n_1072),
.C(n_1065),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1069),
.A2(n_825),
.B(n_973),
.C(n_1018),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1160)
);

BUFx8_ASAP7_75t_L g1161 ( 
.A(n_970),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_L g1162 ( 
.A(n_1072),
.B(n_483),
.C(n_689),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1079),
.B(n_678),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_964),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_987),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1019),
.B(n_825),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1074),
.B(n_1066),
.Y(n_1168)
);

CKINVDCx11_ASAP7_75t_R g1169 ( 
.A(n_953),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1019),
.B(n_825),
.Y(n_1170)
);

AO32x2_ASAP7_75t_L g1171 ( 
.A1(n_954),
.A2(n_956),
.A3(n_965),
.B1(n_945),
.B2(n_414),
.Y(n_1171)
);

BUFx24_ASAP7_75t_L g1172 ( 
.A(n_974),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1069),
.A2(n_825),
.B(n_973),
.C(n_1018),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_960),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_998),
.A2(n_1055),
.A3(n_851),
.B(n_1029),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_SL g1177 ( 
.A(n_1044),
.B(n_1075),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1075),
.A2(n_825),
.B(n_1080),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1017),
.A2(n_1043),
.B(n_1021),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_998),
.A2(n_1055),
.A3(n_851),
.B(n_1029),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1069),
.A2(n_825),
.B(n_973),
.C(n_1018),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1183)
);

NAND3x1_ASAP7_75t_L g1184 ( 
.A(n_1066),
.B(n_1076),
.C(n_1074),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1017),
.A2(n_1043),
.B(n_1021),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1017),
.A2(n_1043),
.B(n_1021),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1072),
.A2(n_689),
.B(n_483),
.C(n_1069),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_946),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_SL g1190 ( 
.A(n_1066),
.B(n_1076),
.C(n_483),
.Y(n_1190)
);

AOI221x1_ASAP7_75t_L g1191 ( 
.A1(n_1001),
.A2(n_1072),
.B1(n_1013),
.B2(n_589),
.C(n_1041),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1079),
.B(n_678),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1064),
.A2(n_541),
.B1(n_991),
.B2(n_494),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1079),
.B(n_678),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1014),
.B(n_860),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1019),
.B(n_825),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1069),
.A2(n_825),
.B(n_973),
.C(n_1018),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_946),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1079),
.B(n_678),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1075),
.A2(n_1080),
.B(n_1072),
.C(n_1065),
.Y(n_1202)
);

AOI21x1_ASAP7_75t_L g1203 ( 
.A1(n_981),
.A2(n_1017),
.B(n_1061),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1019),
.B(n_825),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1021),
.A2(n_1043),
.B(n_981),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1064),
.A2(n_541),
.B1(n_991),
.B2(n_494),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_981),
.A2(n_999),
.B(n_1046),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1017),
.A2(n_1043),
.B(n_1021),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1047),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1075),
.A2(n_825),
.B(n_1080),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_999),
.A2(n_981),
.B(n_1063),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1032),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1081),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1152),
.A2(n_1168),
.B1(n_1088),
.B2(n_1184),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1167),
.A2(n_1204),
.B1(n_1170),
.B2(n_1198),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1194),
.A2(n_1206),
.B1(n_1190),
.B2(n_1204),
.Y(n_1216)
);

INVx6_ASAP7_75t_L g1217 ( 
.A(n_1161),
.Y(n_1217)
);

INVx6_ASAP7_75t_L g1218 ( 
.A(n_1161),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1167),
.A2(n_1170),
.B1(n_1198),
.B2(n_1104),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1106),
.Y(n_1220)
);

INVx4_ASAP7_75t_L g1221 ( 
.A(n_1169),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1101),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1083),
.B(n_1109),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_SL g1224 ( 
.A1(n_1104),
.A2(n_1146),
.B(n_1187),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1114),
.A2(n_1115),
.B1(n_1098),
.B2(n_1109),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_1098),
.A2(n_1114),
.B1(n_1115),
.B2(n_1116),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1172),
.Y(n_1227)
);

CKINVDCx11_ASAP7_75t_R g1228 ( 
.A(n_1209),
.Y(n_1228)
);

INVx8_ASAP7_75t_L g1229 ( 
.A(n_1209),
.Y(n_1229)
);

BUFx12f_ASAP7_75t_L g1230 ( 
.A(n_1209),
.Y(n_1230)
);

INVxp67_ASAP7_75t_L g1231 ( 
.A(n_1116),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1084),
.A2(n_1146),
.B1(n_1159),
.B2(n_1174),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1139),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1182),
.A2(n_1199),
.B1(n_1094),
.B2(n_1097),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1127),
.A2(n_1130),
.B1(n_1086),
.B2(n_1210),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1197),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_1112),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1197),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1092),
.B(n_1103),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1163),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1132),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1175),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1094),
.A2(n_1097),
.B1(n_1087),
.B2(n_1162),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1148),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1178),
.A2(n_1210),
.B1(n_1151),
.B2(n_1103),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1178),
.A2(n_1111),
.B1(n_1147),
.B2(n_1090),
.Y(n_1246)
);

NAND2x1p5_ASAP7_75t_L g1247 ( 
.A(n_1122),
.B(n_1136),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1153),
.A2(n_1156),
.B1(n_1173),
.B2(n_1099),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1099),
.A2(n_1102),
.B1(n_1165),
.B2(n_1192),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_1117),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1117),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1166),
.Y(n_1252)
);

BUFx4_ASAP7_75t_SL g1253 ( 
.A(n_1195),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1165),
.A2(n_1201),
.B1(n_1105),
.B2(n_1212),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1107),
.A2(n_1191),
.B1(n_1200),
.B2(n_1189),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1154),
.B(n_1149),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1100),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1124),
.A2(n_1121),
.B1(n_1141),
.B2(n_1171),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1124),
.A2(n_1171),
.B1(n_1129),
.B2(n_1134),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1171),
.A2(n_1129),
.B1(n_1134),
.B2(n_1131),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1137),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1129),
.A2(n_1135),
.B1(n_1122),
.B2(n_1131),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1135),
.A2(n_1138),
.B1(n_1211),
.B2(n_1181),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1100),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1145),
.Y(n_1265)
);

CKINVDCx11_ASAP7_75t_R g1266 ( 
.A(n_1158),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1138),
.A2(n_1202),
.B1(n_1133),
.B2(n_1113),
.Y(n_1267)
);

BUFx12f_ASAP7_75t_L g1268 ( 
.A(n_1144),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1143),
.A2(n_1133),
.B1(n_1113),
.B2(n_1125),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1123),
.A2(n_1128),
.B1(n_1150),
.B2(n_1164),
.Y(n_1270)
);

BUFx2_ASAP7_75t_SL g1271 ( 
.A(n_1126),
.Y(n_1271)
);

INVxp67_ASAP7_75t_SL g1272 ( 
.A(n_1096),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1142),
.B(n_1120),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1082),
.A2(n_1188),
.B1(n_1193),
.B2(n_1196),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1177),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1118),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1119),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1096),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1123),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1143),
.B(n_1120),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1160),
.A2(n_1183),
.B1(n_1207),
.B2(n_1108),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1207),
.A2(n_1110),
.B(n_1089),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1205),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1095),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1140),
.Y(n_1285)
);

BUFx8_ASAP7_75t_L g1286 ( 
.A(n_1093),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1093),
.Y(n_1287)
);

INVx6_ASAP7_75t_L g1288 ( 
.A(n_1093),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_1205),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1203),
.A2(n_1085),
.B1(n_1176),
.B2(n_1155),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1085),
.B(n_1180),
.Y(n_1291)
);

CKINVDCx11_ASAP7_75t_R g1292 ( 
.A(n_1176),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1091),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1157),
.A2(n_1179),
.B1(n_1185),
.B2(n_1186),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1208),
.Y(n_1295)
);

INVx6_ASAP7_75t_L g1296 ( 
.A(n_1161),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1161),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1169),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1081),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1152),
.A2(n_1168),
.B1(n_1088),
.B2(n_1066),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_1163),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1101),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1161),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1098),
.A2(n_991),
.B1(n_589),
.B2(n_414),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1152),
.A2(n_1168),
.B1(n_1088),
.B2(n_1066),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1081),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1083),
.B(n_1109),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1083),
.B(n_1109),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1209),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1167),
.A2(n_1198),
.B1(n_1170),
.B2(n_1204),
.Y(n_1310)
);

BUFx8_ASAP7_75t_SL g1311 ( 
.A(n_1209),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1167),
.A2(n_1198),
.B1(n_1170),
.B2(n_1204),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1081),
.Y(n_1313)
);

INVx4_ASAP7_75t_L g1314 ( 
.A(n_1169),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1161),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1280),
.B(n_1213),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1261),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1291),
.B(n_1287),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1284),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_L g1320 ( 
.A(n_1300),
.B(n_1305),
.C(n_1224),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1284),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1291),
.B(n_1287),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1273),
.B(n_1288),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1220),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1283),
.B(n_1272),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1269),
.B(n_1265),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1278),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1223),
.B(n_1307),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1299),
.Y(n_1329)
);

AOI21xp33_ASAP7_75t_L g1330 ( 
.A1(n_1214),
.A2(n_1232),
.B(n_1304),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1306),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1215),
.B(n_1310),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1313),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1308),
.B(n_1249),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1295),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1290),
.A2(n_1282),
.B(n_1272),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1277),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1236),
.B(n_1238),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1248),
.B(n_1231),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_SL g1340 ( 
.A(n_1231),
.B(n_1262),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1274),
.A2(n_1270),
.B(n_1293),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1290),
.A2(n_1255),
.B(n_1262),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1248),
.B(n_1225),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1286),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1270),
.A2(n_1258),
.B(n_1259),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1246),
.A2(n_1263),
.B(n_1258),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1259),
.A2(n_1256),
.B(n_1225),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1289),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1271),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1285),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1285),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1285),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1304),
.A2(n_1260),
.B1(n_1279),
.B2(n_1226),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1281),
.B(n_1260),
.Y(n_1354)
);

CKINVDCx6p67_ASAP7_75t_R g1355 ( 
.A(n_1266),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1234),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1292),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1292),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1226),
.A2(n_1216),
.B1(n_1235),
.B2(n_1266),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1268),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1243),
.A2(n_1235),
.B(n_1216),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1310),
.B(n_1312),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1222),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1217),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1312),
.B(n_1219),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1254),
.A2(n_1245),
.B(n_1247),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1239),
.B(n_1242),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1222),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1267),
.Y(n_1369)
);

AO21x2_ASAP7_75t_L g1370 ( 
.A1(n_1255),
.A2(n_1294),
.B(n_1281),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1254),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1294),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1249),
.B(n_1301),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1245),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1240),
.A2(n_1227),
.B1(n_1218),
.B2(n_1296),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1238),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1276),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1250),
.A2(n_1251),
.B(n_1257),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1275),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1275),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1264),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1217),
.A2(n_1218),
.B1(n_1296),
.B2(n_1241),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1217),
.A2(n_1218),
.B1(n_1296),
.B2(n_1252),
.Y(n_1383)
);

AOI221x1_ASAP7_75t_SL g1384 ( 
.A1(n_1320),
.A2(n_1228),
.B1(n_1253),
.B2(n_1311),
.C(n_1229),
.Y(n_1384)
);

NAND4xp25_ASAP7_75t_L g1385 ( 
.A(n_1320),
.B(n_1250),
.C(n_1251),
.D(n_1221),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1357),
.B(n_1315),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1328),
.B(n_1303),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1361),
.A2(n_1297),
.B(n_1244),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_SL g1389 ( 
.A1(n_1361),
.A2(n_1221),
.B(n_1314),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1353),
.A2(n_1330),
.B1(n_1354),
.B2(n_1359),
.Y(n_1390)
);

AND2x2_ASAP7_75t_SL g1391 ( 
.A(n_1340),
.B(n_1314),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_SL g1392 ( 
.A1(n_1378),
.A2(n_1309),
.B(n_1237),
.C(n_1229),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1325),
.B(n_1237),
.Y(n_1393)
);

O2A1O1Ixp5_ASAP7_75t_L g1394 ( 
.A1(n_1330),
.A2(n_1311),
.B(n_1302),
.C(n_1230),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1332),
.B(n_1302),
.C(n_1233),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1340),
.A2(n_1298),
.B1(n_1369),
.B2(n_1365),
.Y(n_1396)
);

AO32x2_ASAP7_75t_L g1397 ( 
.A1(n_1364),
.A2(n_1328),
.A3(n_1316),
.B1(n_1334),
.B2(n_1371),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1332),
.A2(n_1362),
.B(n_1365),
.C(n_1369),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1357),
.B(n_1358),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1362),
.A2(n_1354),
.B1(n_1356),
.B2(n_1374),
.C(n_1343),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1376),
.B(n_1339),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1334),
.B(n_1324),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1377),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1356),
.A2(n_1346),
.B(n_1354),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1376),
.Y(n_1405)
);

AOI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1374),
.A2(n_1343),
.B1(n_1339),
.B2(n_1372),
.C(n_1342),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1346),
.A2(n_1366),
.B(n_1341),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1342),
.A2(n_1367),
.B1(n_1347),
.B2(n_1355),
.Y(n_1408)
);

AO32x2_ASAP7_75t_L g1409 ( 
.A1(n_1364),
.A2(n_1371),
.A3(n_1373),
.B1(n_1347),
.B2(n_1342),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1346),
.A2(n_1366),
.B(n_1377),
.C(n_1326),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1366),
.A2(n_1341),
.B(n_1347),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1318),
.B(n_1322),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1355),
.A2(n_1382),
.B1(n_1375),
.B2(n_1364),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1342),
.A2(n_1347),
.B1(n_1355),
.B2(n_1326),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1349),
.B(n_1347),
.C(n_1337),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1368),
.B(n_1363),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1370),
.A2(n_1349),
.B(n_1381),
.C(n_1379),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1338),
.B(n_1380),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1329),
.B(n_1331),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1370),
.A2(n_1381),
.B(n_1319),
.C(n_1336),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1382),
.A2(n_1375),
.B1(n_1383),
.B2(n_1373),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1363),
.Y(n_1422)
);

AO32x2_ASAP7_75t_L g1423 ( 
.A1(n_1345),
.A2(n_1319),
.A3(n_1333),
.B1(n_1331),
.B2(n_1329),
.Y(n_1423)
);

OR2x6_ASAP7_75t_L g1424 ( 
.A(n_1323),
.B(n_1326),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1370),
.A2(n_1333),
.B1(n_1317),
.B2(n_1321),
.C(n_1336),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1352),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1412),
.B(n_1322),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1423),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1412),
.B(n_1352),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1408),
.A2(n_1363),
.B(n_1344),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1401),
.B(n_1336),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1404),
.B(n_1336),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1404),
.B(n_1341),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1423),
.Y(n_1434)
);

NOR2xp67_ASAP7_75t_L g1435 ( 
.A(n_1415),
.B(n_1348),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1390),
.A2(n_1345),
.B1(n_1370),
.B2(n_1360),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1423),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1403),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1419),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1419),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1398),
.A2(n_1345),
.B1(n_1360),
.B2(n_1351),
.C(n_1350),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1397),
.B(n_1335),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1402),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1397),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1407),
.B(n_1345),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1405),
.B(n_1327),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1425),
.B(n_1417),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1406),
.B(n_1317),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1407),
.B(n_1345),
.Y(n_1449)
);

INVxp67_ASAP7_75t_SL g1450 ( 
.A(n_1415),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1442),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1446),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1446),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1431),
.B(n_1410),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1446),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1431),
.B(n_1414),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1431),
.B(n_1411),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1433),
.B(n_1411),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1436),
.A2(n_1406),
.B1(n_1400),
.B2(n_1391),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1442),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1450),
.B(n_1387),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1428),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1436),
.A2(n_1400),
.B1(n_1396),
.B2(n_1421),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1444),
.B(n_1387),
.Y(n_1464)
);

NOR3xp33_ASAP7_75t_L g1465 ( 
.A(n_1450),
.B(n_1388),
.C(n_1420),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1442),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1433),
.B(n_1418),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1428),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1433),
.B(n_1409),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1432),
.B(n_1409),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1434),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1432),
.B(n_1409),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1434),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1438),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1434),
.B(n_1399),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1434),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1432),
.B(n_1426),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1427),
.B(n_1424),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1427),
.B(n_1393),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1437),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1437),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1461),
.B(n_1452),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1471),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1461),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1477),
.B(n_1427),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1478),
.B(n_1435),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1451),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1477),
.B(n_1435),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1451),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1452),
.B(n_1439),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1463),
.A2(n_1421),
.B1(n_1447),
.B2(n_1413),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1453),
.B(n_1439),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1474),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1471),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1460),
.B(n_1437),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1453),
.B(n_1440),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1464),
.B(n_1440),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1455),
.B(n_1465),
.Y(n_1498)
);

AND2x4_ASAP7_75t_SL g1499 ( 
.A(n_1478),
.B(n_1429),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1474),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1476),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1455),
.B(n_1465),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1464),
.B(n_1443),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1476),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1464),
.B(n_1443),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1462),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1498),
.A2(n_1481),
.B(n_1480),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1501),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1503),
.B(n_1475),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1501),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1491),
.B(n_1458),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1503),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1503),
.B(n_1475),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1491),
.A2(n_1463),
.B1(n_1447),
.B2(n_1441),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1505),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1505),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1499),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1484),
.B(n_1458),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1505),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1484),
.B(n_1458),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1500),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1499),
.B(n_1467),
.Y(n_1522)
);

NOR2xp67_ASAP7_75t_SL g1523 ( 
.A(n_1500),
.B(n_1395),
.Y(n_1523)
);

AOI211xp5_ASAP7_75t_L g1524 ( 
.A1(n_1498),
.A2(n_1430),
.B(n_1413),
.C(n_1441),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1502),
.B(n_1458),
.Y(n_1525)
);

NAND2x1_ASAP7_75t_L g1526 ( 
.A(n_1488),
.B(n_1474),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1502),
.A2(n_1463),
.B(n_1454),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1499),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1482),
.B(n_1457),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1482),
.B(n_1457),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1506),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1499),
.B(n_1467),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1485),
.B(n_1488),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1497),
.B(n_1475),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1487),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1506),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1490),
.B(n_1457),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1490),
.B(n_1457),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1483),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1485),
.B(n_1467),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1492),
.B(n_1454),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1497),
.B(n_1466),
.Y(n_1542)
);

AOI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1486),
.A2(n_1459),
.B1(n_1469),
.B2(n_1445),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1486),
.A2(n_1459),
.B1(n_1469),
.B2(n_1445),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1485),
.B(n_1479),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1486),
.A2(n_1469),
.B1(n_1445),
.B2(n_1449),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1504),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1422),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1539),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1539),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1507),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1522),
.B(n_1532),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1508),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1507),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1510),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1522),
.B(n_1488),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1532),
.B(n_1500),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1540),
.B(n_1500),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1540),
.B(n_1546),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1523),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1512),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1546),
.B(n_1500),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1515),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1525),
.B(n_1492),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1527),
.B(n_1504),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1507),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1516),
.B(n_1496),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1519),
.B(n_1496),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1526),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1517),
.B(n_1493),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1535),
.A2(n_1494),
.B(n_1483),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1541),
.B(n_1497),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1518),
.B(n_1462),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1531),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1520),
.B(n_1509),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1521),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1536),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1545),
.B(n_1548),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1513),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1534),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1521),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1535),
.Y(n_1583)
);

NOR2xp67_ASAP7_75t_L g1584 ( 
.A(n_1570),
.B(n_1517),
.Y(n_1584)
);

AOI22x1_ASAP7_75t_SL g1585 ( 
.A1(n_1577),
.A2(n_1493),
.B1(n_1385),
.B2(n_1494),
.Y(n_1585)
);

NAND2xp33_ASAP7_75t_R g1586 ( 
.A(n_1582),
.B(n_1493),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1566),
.B(n_1543),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1550),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1567),
.A2(n_1472),
.B1(n_1470),
.B2(n_1388),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1550),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1582),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1566),
.A2(n_1514),
.B(n_1524),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1561),
.A2(n_1544),
.B1(n_1547),
.B2(n_1514),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1551),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1577),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1567),
.A2(n_1472),
.B1(n_1470),
.B2(n_1454),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1551),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1552),
.A2(n_1472),
.B1(n_1470),
.B2(n_1449),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1580),
.B(n_1529),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1560),
.B(n_1528),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1579),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1561),
.A2(n_1528),
.B1(n_1530),
.B2(n_1537),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_L g1603 ( 
.A(n_1552),
.B(n_1395),
.C(n_1394),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1571),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1580),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1552),
.A2(n_1538),
.B(n_1472),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1579),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1562),
.Y(n_1608)
);

O2A1O1Ixp33_ASAP7_75t_L g1609 ( 
.A1(n_1592),
.A2(n_1555),
.B(n_1556),
.C(n_1554),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1595),
.B(n_1549),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1605),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1586),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1608),
.Y(n_1613)
);

OAI32xp33_ASAP7_75t_L g1614 ( 
.A1(n_1587),
.A2(n_1555),
.A3(n_1565),
.B1(n_1581),
.B2(n_1573),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1588),
.Y(n_1615)
);

AOI21xp33_ASAP7_75t_L g1616 ( 
.A1(n_1593),
.A2(n_1555),
.B(n_1562),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1591),
.B(n_1581),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1589),
.A2(n_1583),
.B(n_1556),
.Y(n_1618)
);

OAI32xp33_ASAP7_75t_L g1619 ( 
.A1(n_1603),
.A2(n_1565),
.A3(n_1573),
.B1(n_1576),
.B2(n_1568),
.Y(n_1619)
);

NAND2xp33_ASAP7_75t_SL g1620 ( 
.A(n_1600),
.B(n_1558),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1601),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1591),
.B(n_1554),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1589),
.A2(n_1583),
.B(n_1572),
.Y(n_1623)
);

AOI222xp33_ASAP7_75t_L g1624 ( 
.A1(n_1607),
.A2(n_1564),
.B1(n_1456),
.B2(n_1575),
.C1(n_1578),
.C2(n_1448),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1596),
.A2(n_1456),
.B1(n_1449),
.B2(n_1572),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1590),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1604),
.B(n_1560),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1627),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1618),
.A2(n_1606),
.B1(n_1598),
.B2(n_1603),
.C(n_1602),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1618),
.A2(n_1584),
.B(n_1599),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1617),
.Y(n_1631)
);

XNOR2x2_ASAP7_75t_L g1632 ( 
.A(n_1623),
.B(n_1594),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1622),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1611),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1613),
.Y(n_1635)
);

AOI21xp33_ASAP7_75t_SL g1636 ( 
.A1(n_1609),
.A2(n_1597),
.B(n_1578),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1615),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1626),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1629),
.A2(n_1625),
.B1(n_1612),
.B2(n_1610),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1631),
.A2(n_1616),
.B1(n_1624),
.B2(n_1585),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1628),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1631),
.B(n_1576),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1633),
.B(n_1614),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1630),
.B(n_1621),
.Y(n_1644)
);

AND4x1_ASAP7_75t_L g1645 ( 
.A(n_1634),
.B(n_1416),
.C(n_1558),
.D(n_1553),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1636),
.B(n_1620),
.C(n_1575),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1632),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1642),
.Y(n_1648)
);

NOR4xp25_ASAP7_75t_L g1649 ( 
.A(n_1647),
.B(n_1644),
.C(n_1643),
.D(n_1639),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1641),
.B(n_1635),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1640),
.A2(n_1638),
.B1(n_1637),
.B2(n_1572),
.C(n_1564),
.Y(n_1651)
);

OAI211xp5_ASAP7_75t_L g1652 ( 
.A1(n_1646),
.A2(n_1619),
.B(n_1570),
.C(n_1572),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1649),
.B(n_1645),
.C(n_1571),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1648),
.Y(n_1654)
);

NAND4xp75_ASAP7_75t_L g1655 ( 
.A(n_1652),
.B(n_1572),
.C(n_1563),
.D(n_1553),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1650),
.Y(n_1656)
);

NOR2xp67_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_1570),
.Y(n_1657)
);

AO22x2_ASAP7_75t_L g1658 ( 
.A1(n_1652),
.A2(n_1570),
.B1(n_1559),
.B2(n_1563),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1654),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1656),
.B(n_1521),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1653),
.B(n_1559),
.Y(n_1661)
);

XNOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1655),
.B(n_1574),
.Y(n_1662)
);

NAND4xp75_ASAP7_75t_L g1663 ( 
.A(n_1657),
.B(n_1560),
.C(n_1557),
.D(n_1568),
.Y(n_1663)
);

OAI211xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1659),
.A2(n_1658),
.B(n_1569),
.C(n_1574),
.Y(n_1664)
);

INVxp33_ASAP7_75t_SL g1665 ( 
.A(n_1660),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1662),
.A2(n_1569),
.B1(n_1557),
.B2(n_1495),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1665),
.B(n_1661),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1667),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1668),
.B(n_1664),
.Y(n_1669)
);

OAI21xp33_ASAP7_75t_L g1670 ( 
.A1(n_1668),
.A2(n_1666),
.B(n_1663),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1669),
.A2(n_1468),
.B1(n_1473),
.B2(n_1481),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1670),
.B(n_1483),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1672),
.A2(n_1671),
.B(n_1533),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1672),
.A2(n_1542),
.B1(n_1494),
.B2(n_1533),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1542),
.B1(n_1487),
.B2(n_1489),
.Y(n_1675)
);

NOR2xp67_ASAP7_75t_L g1676 ( 
.A(n_1675),
.B(n_1673),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1473),
.B1(n_1468),
.B2(n_1480),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_R g1678 ( 
.A1(n_1677),
.A2(n_1493),
.B1(n_1384),
.B2(n_1392),
.C(n_1389),
.Y(n_1678)
);

AOI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1385),
.B(n_1386),
.C(n_1493),
.Y(n_1679)
);


endmodule