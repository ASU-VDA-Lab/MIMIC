module fake_netlist_6_4095_n_6 (n_1, n_0, n_2, n_6);

input n_1;
input n_0;
input n_2;

output n_6;

wire n_4;
wire n_3;
wire n_5;

INVx3_ASAP7_75t_L g3 ( 
.A(n_2),
.Y(n_3)
);

CKINVDCx6p67_ASAP7_75t_R g4 ( 
.A(n_1),
.Y(n_4)
);

AOI22xp5_ASAP7_75t_L g5 ( 
.A1(n_4),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);


endmodule