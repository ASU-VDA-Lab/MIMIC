module fake_jpeg_15815_n_357 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_357);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_357;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_2),
.B(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_0),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_53),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_36),
.B1(n_29),
.B2(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_24),
.B1(n_58),
.B2(n_51),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_64),
.B(n_66),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_36),
.B1(n_33),
.B2(n_23),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_58),
.B1(n_51),
.B2(n_36),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_43),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_91),
.Y(n_99)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_33),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_52),
.Y(n_109)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

OR2x4_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_26),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_92),
.A2(n_114),
.B1(n_67),
.B2(n_40),
.Y(n_143)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_100),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_50),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_57),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

CKINVDCx12_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_111),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_108),
.Y(n_132)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_115),
.Y(n_128)
);

CKINVDCx6p67_ASAP7_75t_R g110 ( 
.A(n_77),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_49),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_58),
.B1(n_24),
.B2(n_56),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_90),
.B1(n_70),
.B2(n_72),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_123),
.Y(n_130)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_78),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_80),
.B1(n_73),
.B2(n_81),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_68),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_145),
.C(n_56),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_81),
.B1(n_74),
.B2(n_86),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_141),
.B1(n_121),
.B2(n_122),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_136),
.A2(n_139),
.B1(n_142),
.B2(n_35),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_147),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_80),
.B1(n_65),
.B2(n_32),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_143),
.B1(n_148),
.B2(n_149),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_70),
.B1(n_67),
.B2(n_57),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_32),
.B1(n_41),
.B2(n_40),
.Y(n_142)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_102),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_85),
.C(n_53),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_88),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_28),
.B1(n_41),
.B2(n_25),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_157),
.B(n_178),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_164),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_147),
.C(n_140),
.Y(n_191)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_165),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_85),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_116),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_171),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_25),
.B(n_35),
.C(n_34),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_94),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_103),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_176),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_22),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_148),
.B1(n_145),
.B2(n_128),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_179),
.A2(n_199),
.B1(n_170),
.B2(n_124),
.Y(n_214)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_131),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_172),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_125),
.B(n_127),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_197),
.B(n_158),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_194),
.C(n_198),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_166),
.A2(n_126),
.B1(n_110),
.B2(n_127),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_167),
.B1(n_159),
.B2(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_137),
.C(n_151),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_126),
.C(n_137),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_129),
.C(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_177),
.A2(n_146),
.B1(n_124),
.B2(n_57),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_213),
.B1(n_56),
.B2(n_55),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_205),
.Y(n_227)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_207),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_179),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_210),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_214),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_165),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_180),
.B(n_164),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_189),
.A2(n_188),
.B(n_195),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_218),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_157),
.B1(n_175),
.B2(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_176),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_156),
.B(n_178),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_161),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_161),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_221),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_187),
.B(n_186),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_222),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_168),
.B1(n_34),
.B2(n_38),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_1),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_190),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_181),
.B1(n_191),
.B2(n_194),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_236),
.B1(n_200),
.B2(n_213),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_246),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_198),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_234),
.C(n_205),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_197),
.C(n_187),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_181),
.B1(n_197),
.B2(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_110),
.B(n_2),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_249),
.B(n_98),
.Y(n_271)
);

NOR4xp25_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_22),
.C(n_38),
.D(n_169),
.Y(n_239)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_239),
.A2(n_39),
.B(n_214),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_84),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_82),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_204),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_202),
.B(n_169),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_226),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_254),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_201),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_260),
.C(n_262),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_243),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_265),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_210),
.B1(n_216),
.B2(n_221),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_207),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_42),
.B1(n_2),
.B2(n_3),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_206),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_206),
.C(n_203),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_169),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_93),
.C(n_133),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_93),
.C(n_133),
.Y(n_269)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_39),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_246),
.B(n_241),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_271),
.A2(n_53),
.B(n_27),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_250),
.A2(n_233),
.B1(n_235),
.B2(n_237),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_272),
.A2(n_281),
.B1(n_282),
.B2(n_1),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_268),
.A2(n_229),
.B1(n_231),
.B2(n_242),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_245),
.B1(n_238),
.B2(n_246),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_260),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_253),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_278),
.B(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

XNOR2x2_ASAP7_75t_SL g297 ( 
.A(n_277),
.B(n_252),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g319 ( 
.A(n_297),
.B(n_283),
.Y(n_319)
);

AOI221xp5_ASAP7_75t_L g300 ( 
.A1(n_281),
.A2(n_254),
.B1(n_266),
.B2(n_262),
.C(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_278),
.B(n_1),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_303),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_282),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_152),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_27),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_306),
.C(n_279),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_98),
.C(n_82),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_297),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_276),
.B1(n_288),
.B2(n_284),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_308),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_284),
.C(n_287),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_318),
.C(n_306),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_285),
.B(n_273),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_311),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_294),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_283),
.B1(n_290),
.B2(n_272),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_286),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_293),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_321),
.A2(n_316),
.B(n_309),
.C(n_307),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_295),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_292),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_327),
.C(n_55),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_55),
.C(n_27),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_313),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_329),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_315),
.B(n_4),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_42),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_318),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_325),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_332),
.A2(n_324),
.B1(n_10),
.B2(n_11),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_333),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_42),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_327),
.A2(n_6),
.B(n_7),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_335),
.A2(n_9),
.B(n_11),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_339),
.C(n_340),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_7),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_330),
.A2(n_9),
.B(n_10),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_322),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_343),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_336),
.C(n_50),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_345),
.A2(n_9),
.B(n_12),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_346),
.A2(n_333),
.B(n_340),
.Y(n_348)
);

AO21x1_ASAP7_75t_L g351 ( 
.A1(n_348),
.A2(n_349),
.B(n_350),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_347),
.A2(n_342),
.B(n_341),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_12),
.C(n_13),
.Y(n_353)
);

AOI211xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_351),
.B(n_13),
.C(n_14),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_12),
.Y(n_355)
);

AOI321xp33_ASAP7_75t_L g356 ( 
.A1(n_355),
.A2(n_16),
.A3(n_17),
.B1(n_42),
.B2(n_50),
.C(n_345),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_16),
.B(n_17),
.Y(n_357)
);


endmodule