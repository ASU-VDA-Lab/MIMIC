module real_jpeg_908_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_202;
wire n_167;
wire n_128;
wire n_295;
wire n_179;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_44),
.B1(n_50),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_2),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_85),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_2),
.A2(n_29),
.B1(n_35),
.B2(n_85),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_29),
.B1(n_35),
.B2(n_73),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_44),
.B1(n_50),
.B2(n_73),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_4),
.A2(n_50),
.B(n_81),
.C(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_4),
.B(n_50),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_12),
.B(n_50),
.C(n_199),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_8),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_44),
.B1(n_50),
.B2(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_71),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_10),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_10),
.A2(n_44),
.B1(n_50),
.B2(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_149),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_149),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_11),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_44),
.B1(n_50),
.B2(n_104),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_104),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_11),
.A2(n_29),
.B1(n_35),
.B2(n_104),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_12),
.B(n_40),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_12),
.B(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_12),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_12),
.B(n_82),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_12),
.A2(n_44),
.B1(n_50),
.B2(n_200),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_12),
.B(n_29),
.C(n_66),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_200),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_12),
.B(n_32),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_12),
.B(n_98),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_42),
.B1(n_44),
.B2(n_50),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_14),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_14),
.A2(n_29),
.B1(n_35),
.B2(n_42),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_15),
.A2(n_44),
.B1(n_50),
.B2(n_54),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_15),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_15),
.A2(n_29),
.B1(n_35),
.B2(n_54),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_125),
.B1(n_297),
.B2(n_298),
.Y(n_18)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_19),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_108),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_21),
.B(n_108),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_89),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_22),
.A2(n_23),
.B1(n_75),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_74),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_57),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_26),
.A2(n_38),
.B(n_74),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_26),
.A2(n_57),
.B1(n_59),
.B2(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_27),
.A2(n_32),
.B1(n_94),
.B2(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_27),
.A2(n_200),
.B(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_28),
.A2(n_31),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_28),
.A2(n_31),
.B1(n_175),
.B2(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_28),
.B(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_28),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_28),
.A2(n_31),
.B1(n_231),
.B2(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_29),
.A2(n_35),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_29),
.B(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_31),
.A2(n_190),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_31),
.B(n_204),
.Y(n_233)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_32),
.A2(n_203),
.B(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_51),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_39),
.A2(n_43),
.B1(n_105),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI32xp33_ASAP7_75t_L g170 ( 
.A1(n_41),
.A2(n_47),
.A3(n_50),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_41),
.A2(n_105),
.B(n_200),
.C(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_43),
.B(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_43),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_43),
.A2(n_51),
.B(n_164),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_43)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_44),
.B(n_48),
.Y(n_172)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_55),
.A2(n_103),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_59),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_68),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_60),
.A2(n_68),
.B1(n_193),
.B2(n_227),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_60),
.A2(n_195),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_70),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_61),
.A2(n_98),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_97),
.B1(n_98),
.B2(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_61),
.A2(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_61),
.B(n_196),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_63),
.A2(n_83),
.B(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_64),
.B(n_245),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_68),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_68),
.A2(n_216),
.B(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B(n_88),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_78),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_84),
.B1(n_86),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_86),
.B1(n_87),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_79),
.A2(n_166),
.B(n_168),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_79),
.A2(n_168),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_80),
.A2(n_82),
.B1(n_167),
.B2(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_82),
.B(n_146),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_100),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_86),
.A2(n_145),
.B(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.C(n_101),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_91),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_161),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_92),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_98),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_101),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B(n_106),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_107),
.B(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_122),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_121),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_125),
.Y(n_298)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_151),
.B(n_296),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_127),
.B(n_130),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_136),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.C(n_147),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_138),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_139),
.B(n_141),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_140),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_177),
.B(n_295),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_153),
.B(n_155),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_162),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_156),
.B(n_160),
.Y(n_280)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_162),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_169),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_163),
.B(n_165),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_169),
.B(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI31xp33_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_277),
.A3(n_287),
.B(n_292),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_221),
.B(n_276),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_205),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_180),
.B(n_205),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.C(n_197),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_181),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_186),
.C(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_191),
.B(n_197),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_201),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_217),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_206),
.B(n_218),
.C(n_220),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_207),
.B(n_212),
.C(n_213),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_271),
.B(n_275),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_240),
.B(n_270),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_234),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_234),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_229),
.A2(n_230),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_252),
.B(n_269),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_263),
.B(n_268),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B(n_262),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_266),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_274),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_281),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_284),
.Y(n_290)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_291),
.Y(n_293)
);


endmodule