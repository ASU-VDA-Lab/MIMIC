module fake_ariane_1782_n_1930 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1930);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1930;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1803;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_925;
wire n_246;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_134),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_18),
.Y(n_159)
);

BUFx2_ASAP7_75t_SL g160 ( 
.A(n_58),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_97),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_69),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_59),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_21),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_56),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_51),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_5),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_39),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_76),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_75),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_11),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_39),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_8),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_73),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_21),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_49),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_44),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_42),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_137),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_7),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_52),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_85),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_91),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_96),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_41),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_81),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_124),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_88),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_62),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_140),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_144),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_0),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_93),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_22),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_60),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_54),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_24),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_50),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_13),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_22),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_150),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_105),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_28),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_80),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_13),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_26),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_1),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_64),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_104),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_157),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_127),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_38),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_28),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_47),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_98),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_31),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_37),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_128),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_70),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_31),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_156),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_10),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_10),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_130),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_101),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_8),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_121),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_87),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_15),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_1),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_78),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_131),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_114),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_4),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_95),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_138),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_18),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_120),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_79),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_107),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_61),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_154),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_27),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_35),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_16),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_7),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_117),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_143),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_48),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_46),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_84),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_103),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_112),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_71),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_26),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_11),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_67),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_92),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_40),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_68),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_44),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_153),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_30),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_6),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_135),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_41),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_99),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_77),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_14),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_111),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_37),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_115),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_3),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_109),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_24),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_20),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_30),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_34),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_65),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_20),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_106),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_53),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_33),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_25),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_55),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_12),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_90),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_133),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_19),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_2),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_212),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_206),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_180),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_250),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_162),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_162),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_163),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_163),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_167),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_169),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_171),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_179),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_172),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_179),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_172),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_170),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_173),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_201),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_186),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_179),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_180),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_173),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_239),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_178),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_220),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_178),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_270),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_293),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_185),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_159),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_219),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_185),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_187),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_187),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_228),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_195),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_250),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_212),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_257),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_195),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_175),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_196),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_181),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_196),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_188),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_239),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_192),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_197),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_197),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_250),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_215),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_199),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_215),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_264),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_179),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_179),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_224),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_224),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_226),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_226),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_207),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_235),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_230),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_210),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_230),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_264),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_213),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_236),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_217),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_236),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_377),
.A2(n_189),
.B(n_262),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_377),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_319),
.A2(n_299),
.B1(n_252),
.B2(n_244),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_326),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_314),
.B(n_166),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_320),
.B(n_166),
.Y(n_397)
);

AND2x6_ASAP7_75t_L g398 ( 
.A(n_316),
.B(n_189),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_314),
.B(n_319),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_381),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_328),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_316),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_316),
.B(n_237),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_355),
.B(n_237),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_335),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_355),
.B(n_240),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_355),
.B(n_240),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_345),
.A2(n_309),
.B1(n_312),
.B2(n_303),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_337),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_317),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_354),
.B(n_256),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_R g418 ( 
.A(n_359),
.B(n_158),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_317),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_317),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_329),
.B(n_262),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_354),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_331),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_342),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_344),
.Y(n_427)
);

CKINVDCx8_ASAP7_75t_R g428 ( 
.A(n_369),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_333),
.B(n_279),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_361),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_374),
.B(n_272),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_333),
.B(n_279),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_336),
.A2(n_225),
.B1(n_245),
.B2(n_249),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_363),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_321),
.A2(n_189),
.B(n_272),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_369),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_348),
.B(n_227),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_375),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_315),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_317),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_315),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_321),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_322),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_317),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_322),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_317),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_373),
.B(n_295),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_373),
.B(n_295),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_323),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_385),
.A2(n_356),
.B1(n_367),
.B2(n_338),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_323),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_365),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_324),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_385),
.B(n_304),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_324),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_325),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_380),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_325),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_405),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_410),
.B(n_304),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_391),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_429),
.B(n_327),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_418),
.B(n_383),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_392),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_410),
.B(n_305),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_415),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_399),
.B(n_447),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_419),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_425),
.B(n_327),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

INVxp33_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_425),
.B(n_330),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_438),
.B(n_405),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_422),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_422),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_401),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_446),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_406),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_432),
.A2(n_367),
.B1(n_340),
.B2(n_364),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_448),
.B(n_386),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_388),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_330),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_411),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_442),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_416),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_395),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_434),
.B(n_332),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_434),
.B(n_332),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_398),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_414),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_410),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_397),
.B(n_334),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_443),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_394),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_445),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_395),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_394),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_445),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_432),
.B(n_334),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_449),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_458),
.B(n_339),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_424),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_394),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_444),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_L g518 ( 
.A1(n_433),
.A2(n_245),
.B1(n_242),
.B2(n_253),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_444),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_404),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_437),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_453),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_444),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_457),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_409),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_458),
.B(n_339),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_457),
.Y(n_530)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_450),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_396),
.B(n_341),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_441),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_441),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_439),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_407),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_430),
.B(n_341),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_413),
.B(n_343),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_439),
.B(n_343),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_417),
.B(n_408),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_412),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_423),
.B(n_346),
.Y(n_543)
);

AND3x2_ASAP7_75t_L g544 ( 
.A(n_452),
.B(n_455),
.C(n_402),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_431),
.B(n_439),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_451),
.B(n_346),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_456),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_452),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_416),
.Y(n_550)
);

INVx8_ASAP7_75t_L g551 ( 
.A(n_398),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_398),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_416),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_398),
.A2(n_389),
.B1(n_387),
.B2(n_384),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_420),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_455),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_435),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_403),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_420),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_420),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_398),
.B(n_305),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_420),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_435),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_400),
.B(n_349),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_398),
.A2(n_289),
.B1(n_292),
.B2(n_294),
.Y(n_567)
);

AOI21x1_ASAP7_75t_L g568 ( 
.A1(n_420),
.A2(n_351),
.B(n_350),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_436),
.B(n_266),
.Y(n_569)
);

AO22x2_ASAP7_75t_L g570 ( 
.A1(n_393),
.A2(n_389),
.B1(n_387),
.B2(n_384),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_421),
.B(n_353),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_421),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_421),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_421),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_428),
.A2(n_267),
.B1(n_268),
.B2(n_278),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_421),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_440),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_428),
.B(n_353),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_440),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_440),
.B(n_358),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_440),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_404),
.B(n_358),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_440),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_426),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_426),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_427),
.B(n_360),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_427),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_392),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_392),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_391),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_392),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_425),
.B(n_360),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_392),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_392),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_392),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_399),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_405),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_390),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_392),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_405),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_418),
.B(n_362),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_409),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_405),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_392),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_392),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_398),
.B(n_362),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_392),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_437),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_500),
.B(n_366),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_525),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_500),
.B(n_366),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_548),
.B(n_379),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_494),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_560),
.B(n_368),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_525),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_492),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_492),
.B(n_379),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_484),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_541),
.B(n_282),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_597),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_477),
.B(n_164),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_503),
.Y(n_622)
);

AO22x2_ASAP7_75t_L g623 ( 
.A1(n_570),
.A2(n_378),
.B1(n_376),
.B2(n_372),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_503),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_504),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_471),
.B(n_286),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_548),
.B(n_378),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_504),
.B(n_368),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_505),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_505),
.B(n_376),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_507),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_526),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_602),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_507),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_597),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_510),
.B(n_370),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_560),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_551),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_477),
.B(n_370),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_510),
.B(n_372),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_494),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_170),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_486),
.B(n_298),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_512),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_512),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_513),
.B(n_204),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_484),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_558),
.B(n_582),
.Y(n_649)
);

CKINVDCx8_ASAP7_75t_R g650 ( 
.A(n_515),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_558),
.B(n_183),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_513),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_489),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_489),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_582),
.B(n_183),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_551),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_502),
.A2(n_190),
.B1(n_307),
.B2(n_306),
.Y(n_657)
);

OR2x2_ASAP7_75t_SL g658 ( 
.A(n_515),
.B(n_184),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_522),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_487),
.B(n_182),
.Y(n_660)
);

BUFx10_ASAP7_75t_L g661 ( 
.A(n_508),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_522),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_536),
.B(n_218),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_582),
.Y(n_664)
);

INVx3_ASAP7_75t_R g665 ( 
.A(n_521),
.Y(n_665)
);

BUFx4f_ASAP7_75t_L g666 ( 
.A(n_462),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_529),
.B(n_184),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_490),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_508),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_490),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_459),
.B(n_190),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_459),
.B(n_216),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_523),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_523),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_530),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_569),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_530),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_533),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_533),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_529),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_534),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_534),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_464),
.B(n_216),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_566),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_498),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_598),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_498),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_551),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_535),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_462),
.A2(n_221),
.B1(n_307),
.B2(n_306),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_462),
.A2(n_468),
.B1(n_538),
.B2(n_570),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_566),
.B(n_221),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_551),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_535),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_545),
.B(n_202),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_499),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_584),
.B(n_223),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_463),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_481),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_536),
.B(n_238),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_461),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_499),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_464),
.B(n_223),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

NAND3x1_ASAP7_75t_L g705 ( 
.A(n_584),
.B(n_269),
.C(n_231),
.Y(n_705)
);

OAI221xp5_ASAP7_75t_L g706 ( 
.A1(n_532),
.A2(n_231),
.B1(n_301),
.B2(n_300),
.C(n_296),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_461),
.Y(n_707)
);

INVx8_ASAP7_75t_L g708 ( 
.A(n_462),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_584),
.B(n_234),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_511),
.B(n_234),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_477),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_SL g712 ( 
.A(n_585),
.B(n_269),
.C(n_287),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_501),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_520),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_462),
.A2(n_283),
.B1(n_160),
.B2(n_308),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_542),
.B(n_202),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_462),
.A2(n_283),
.B1(n_160),
.B2(n_302),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_467),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_587),
.B(n_287),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_511),
.B(n_296),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_470),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_470),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_501),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_520),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_474),
.Y(n_725)
);

BUFx4f_ASAP7_75t_L g726 ( 
.A(n_462),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_578),
.B(n_300),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_506),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_474),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_542),
.B(n_251),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_506),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_477),
.B(n_251),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_468),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_544),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_497),
.B(n_255),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_495),
.B(n_301),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_596),
.B(n_260),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_496),
.B(n_241),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_509),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_587),
.B(n_264),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_589),
.Y(n_741)
);

CKINVDCx16_ASAP7_75t_R g742 ( 
.A(n_569),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_509),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_516),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_497),
.B(n_255),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_516),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_585),
.B(n_2),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_466),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_466),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_469),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_589),
.Y(n_751)
);

NAND2x1p5_ASAP7_75t_L g752 ( 
.A(n_497),
.B(n_241),
.Y(n_752)
);

AO22x2_ASAP7_75t_L g753 ( 
.A1(n_570),
.A2(n_265),
.B1(n_285),
.B2(n_274),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_593),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_596),
.B(n_5),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_539),
.B(n_265),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_469),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_468),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_593),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_467),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_598),
.Y(n_761)
);

NAND2x1p5_ASAP7_75t_L g762 ( 
.A(n_497),
.B(n_274),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_539),
.B(n_161),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_594),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_514),
.B(n_285),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_596),
.B(n_6),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_528),
.B(n_311),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_547),
.B(n_165),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_586),
.B(n_311),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_521),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_594),
.Y(n_771)
);

OR2x2_ASAP7_75t_SL g772 ( 
.A(n_531),
.B(n_206),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_601),
.B(n_12),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_595),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_595),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_538),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_570),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_596),
.Y(n_778)
);

AND2x6_ASAP7_75t_L g779 ( 
.A(n_567),
.B(n_206),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_537),
.B(n_17),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_472),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_538),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_649),
.B(n_460),
.Y(n_784)
);

AND2x2_ASAP7_75t_SL g785 ( 
.A(n_691),
.B(n_567),
.Y(n_785)
);

OAI21xp33_ASAP7_75t_L g786 ( 
.A1(n_619),
.A2(n_465),
.B(n_518),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_648),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_660),
.A2(n_468),
.B1(n_538),
.B2(n_460),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_619),
.B(n_468),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_666),
.B(n_598),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_699),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_666),
.B(n_726),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_660),
.B(n_468),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_653),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_644),
.A2(n_543),
.B(n_607),
.C(n_599),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_616),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_622),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_647),
.A2(n_604),
.B(n_599),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_624),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_625),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_614),
.B(n_608),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_630),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_708),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_632),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_SL g805 ( 
.A(n_644),
.B(n_475),
.C(n_608),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_726),
.B(n_598),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_654),
.Y(n_807)
);

AO21x2_ASAP7_75t_L g808 ( 
.A1(n_647),
.A2(n_607),
.B(n_604),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_663),
.B(n_468),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_663),
.B(n_473),
.Y(n_810)
);

AND3x1_ASAP7_75t_L g811 ( 
.A(n_780),
.B(n_485),
.C(n_546),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_708),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_668),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_737),
.B(n_538),
.C(n_575),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_777),
.A2(n_547),
.B1(n_549),
.B2(n_527),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_708),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_609),
.B(n_476),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_711),
.B(n_598),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_664),
.B(n_478),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_670),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_711),
.A2(n_559),
.B(n_565),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_635),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_686),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_686),
.A2(n_559),
.B(n_565),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_633),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_609),
.B(n_488),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_685),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_611),
.B(n_737),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_613),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_611),
.B(n_592),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_645),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_634),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_649),
.B(n_603),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_740),
.B(n_697),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_642),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_638),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_638),
.B(n_603),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_687),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_646),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_777),
.A2(n_549),
.B1(n_527),
.B2(n_472),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_709),
.B(n_600),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_652),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_669),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_696),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_684),
.B(n_479),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_777),
.A2(n_480),
.B1(n_605),
.B2(n_591),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_691),
.A2(n_623),
.B1(n_753),
.B2(n_779),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_640),
.B(n_467),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_718),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_698),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_700),
.B(n_479),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_770),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_700),
.B(n_480),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_732),
.A2(n_491),
.B(n_482),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_702),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_706),
.A2(n_684),
.B1(n_712),
.B2(n_664),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_SL g857 ( 
.A(n_778),
.B(n_482),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_612),
.B(n_588),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_623),
.A2(n_605),
.B1(n_591),
.B2(n_588),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_612),
.B(n_483),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_713),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_627),
.B(n_553),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_718),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_627),
.B(n_555),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_633),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_640),
.B(n_483),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_723),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_680),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_659),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_643),
.B(n_563),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_662),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_673),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_716),
.B(n_563),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_680),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_674),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_716),
.B(n_563),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_623),
.A2(n_563),
.B1(n_606),
.B2(n_580),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_675),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_667),
.B(n_571),
.Y(n_879)
);

BUFx4f_ASAP7_75t_L g880 ( 
.A(n_724),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_730),
.B(n_563),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_753),
.A2(n_563),
.B1(n_540),
.B2(n_483),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_SL g883 ( 
.A1(n_706),
.A2(n_776),
.B1(n_782),
.B2(n_773),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_677),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_730),
.B(n_563),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_610),
.B(n_540),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_650),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_615),
.B(n_540),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_661),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_763),
.B(n_517),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_763),
.B(n_517),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_620),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_620),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_753),
.A2(n_519),
.B1(n_524),
.B2(n_491),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_SL g895 ( 
.A1(n_676),
.A2(n_211),
.B1(n_203),
.B2(n_200),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_678),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_661),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_719),
.B(n_519),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_773),
.A2(n_214),
.B1(n_205),
.B2(n_198),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_692),
.B(n_524),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_626),
.B(n_552),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_671),
.B(n_552),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_714),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_626),
.B(n_552),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_772),
.B(n_554),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_679),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_655),
.B(n_755),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_681),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_682),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_655),
.B(n_554),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_733),
.B(n_554),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_701),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_755),
.B(n_562),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_779),
.A2(n_583),
.B1(n_581),
.B2(n_550),
.Y(n_914)
);

AND2x6_ASAP7_75t_SL g915 ( 
.A(n_651),
.B(n_574),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_714),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_671),
.B(n_562),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_707),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_721),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_620),
.Y(n_920)
);

BUFx4f_ASAP7_75t_L g921 ( 
.A(n_636),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_779),
.A2(n_583),
.B1(n_581),
.B2(n_550),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_704),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_748),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_672),
.B(n_579),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_733),
.B(n_562),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_766),
.A2(n_574),
.B1(n_579),
.B2(n_557),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_704),
.B(n_579),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_722),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_749),
.Y(n_930)
);

OAI22x1_ASAP7_75t_R g931 ( 
.A1(n_676),
.A2(n_194),
.B1(n_310),
.B2(n_297),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_758),
.B(n_568),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_766),
.B(n_557),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_725),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_672),
.B(n_568),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_729),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_741),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_686),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_SL g939 ( 
.A(n_747),
.B(n_493),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_636),
.B(n_561),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_SL g941 ( 
.A1(n_742),
.A2(n_177),
.B1(n_291),
.B2(n_290),
.Y(n_941)
);

CKINVDCx8_ASAP7_75t_R g942 ( 
.A(n_651),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_760),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_751),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_636),
.B(n_561),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_760),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_734),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_734),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_683),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_688),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_629),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_683),
.B(n_564),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_779),
.A2(n_577),
.B1(n_573),
.B2(n_572),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_703),
.B(n_564),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_703),
.B(n_572),
.Y(n_955)
);

AND2x6_ASAP7_75t_SL g956 ( 
.A(n_780),
.B(n_17),
.Y(n_956)
);

BUFx6f_ASAP7_75t_SL g957 ( 
.A(n_710),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_689),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_768),
.B(n_573),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_761),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_754),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_710),
.B(n_577),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_750),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_657),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_779),
.A2(n_254),
.B1(n_176),
.B2(n_191),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_657),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_720),
.B(n_576),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_720),
.B(n_576),
.Y(n_968)
);

BUFx4f_ASAP7_75t_L g969 ( 
.A(n_736),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_690),
.A2(n_758),
.B1(n_712),
.B2(n_736),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_SL g971 ( 
.A1(n_617),
.A2(n_19),
.B(n_23),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_690),
.A2(n_206),
.B1(n_168),
.B2(n_248),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_694),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_761),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_688),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_964),
.B(n_665),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_783),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_832),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_786),
.A2(n_617),
.B(n_641),
.C(n_637),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_783),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_832),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_791),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_812),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_829),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_787),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_789),
.B(n_761),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_810),
.B(n_727),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_787),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_794),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_966),
.B(n_658),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_828),
.B(n_727),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_834),
.B(n_628),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_791),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_801),
.B(n_969),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_796),
.Y(n_995)
);

AOI221xp5_ASAP7_75t_L g996 ( 
.A1(n_856),
.A2(n_738),
.B1(n_765),
.B2(n_767),
.C(n_769),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_845),
.B(n_628),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_817),
.B(n_631),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_812),
.Y(n_999)
);

O2A1O1Ixp5_ASAP7_75t_L g1000 ( 
.A1(n_795),
.A2(n_621),
.B(n_768),
.C(n_637),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_826),
.B(n_631),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_830),
.B(n_879),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_812),
.B(n_629),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_856),
.B(n_641),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_887),
.Y(n_1005)
);

AND3x1_ASAP7_75t_SL g1006 ( 
.A(n_956),
.B(n_759),
.C(n_764),
.Y(n_1006)
);

OA22x2_ASAP7_75t_L g1007 ( 
.A1(n_949),
.A2(n_767),
.B1(n_765),
.B2(n_738),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_860),
.B(n_756),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_812),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_836),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_797),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_794),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_948),
.B(n_629),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_860),
.B(n_756),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_807),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_835),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_807),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_821),
.A2(n_693),
.B(n_656),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_907),
.B(n_771),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_813),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_819),
.B(n_774),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_813),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_836),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_819),
.B(n_775),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_950),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_951),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_825),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_820),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_837),
.B(n_769),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_799),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_865),
.Y(n_1031)
);

NAND2x1_ASAP7_75t_L g1032 ( 
.A(n_951),
.B(n_757),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_784),
.B(n_695),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_903),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_800),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_824),
.A2(n_639),
.B(n_693),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_820),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_843),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_784),
.B(n_695),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_923),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_827),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_833),
.B(n_705),
.Y(n_1042)
);

NOR2x1p5_ASAP7_75t_L g1043 ( 
.A(n_887),
.B(n_781),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_923),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_827),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_803),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_809),
.B(n_621),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_844),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_948),
.B(n_629),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_844),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_814),
.B(n_728),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_889),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_855),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_880),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_802),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_855),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_793),
.B(n_715),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_788),
.B(n_717),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_833),
.B(n_731),
.Y(n_1059)
);

CKINVDCx16_ASAP7_75t_R g1060 ( 
.A(n_931),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_804),
.Y(n_1061)
);

OR2x6_ASAP7_75t_L g1062 ( 
.A(n_852),
.B(n_752),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_822),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_831),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_938),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_938),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_L g1067 ( 
.A(n_795),
.B(n_745),
.C(n_732),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_880),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_839),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_842),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_869),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_969),
.B(n_739),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_921),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_921),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_941),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_924),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_803),
.B(n_639),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_816),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_SL g1079 ( 
.A1(n_785),
.A2(n_762),
.B1(n_752),
.B2(n_639),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_816),
.B(n_639),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_924),
.Y(n_1081)
);

BUFx8_ASAP7_75t_L g1082 ( 
.A(n_957),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_SL g1083 ( 
.A1(n_895),
.A2(n_762),
.B1(n_261),
.B2(n_259),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_871),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_872),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_868),
.B(n_746),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_875),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_878),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_884),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_902),
.B(n_693),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_805),
.A2(n_745),
.B1(n_735),
.B2(n_743),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_930),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_902),
.B(n_693),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_896),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_957),
.A2(n_735),
.B1(n_744),
.B2(n_656),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_906),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_917),
.B(n_656),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_970),
.B(n_576),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_792),
.B(n_656),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_970),
.B(n_576),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_SL g1101 ( 
.A1(n_899),
.A2(n_277),
.B1(n_193),
.B2(n_209),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_874),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_858),
.B(n_917),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_942),
.B(n_883),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_950),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_925),
.Y(n_1106)
);

BUFx2_ASAP7_75t_SL g1107 ( 
.A(n_916),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_930),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_963),
.Y(n_1109)
);

NAND2xp33_ASAP7_75t_L g1110 ( 
.A(n_938),
.B(n_576),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_925),
.B(n_556),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_908),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_909),
.B(n_556),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_892),
.B(n_556),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_950),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_950),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_938),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_933),
.B(n_556),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_912),
.Y(n_1119)
);

AND3x1_ASAP7_75t_L g1120 ( 
.A(n_897),
.B(n_23),
.C(n_25),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_892),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_932),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_963),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_838),
.Y(n_1124)
);

NOR2x1_ASAP7_75t_L g1125 ( 
.A(n_893),
.B(n_556),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_918),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_850),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_928),
.B(n_493),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_919),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_1004),
.B(n_811),
.C(n_971),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_995),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_978),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1021),
.B(n_785),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1011),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_984),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1082),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1030),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1035),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_998),
.B(n_851),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1055),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1001),
.B(n_853),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_990),
.A2(n_905),
.B1(n_935),
.B2(n_864),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1024),
.B(n_847),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_979),
.A2(n_818),
.B(n_848),
.C(n_866),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_979),
.A2(n_933),
.B(n_905),
.C(n_959),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_1082),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1061),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1110),
.A2(n_986),
.B(n_818),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1082),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_984),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1063),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1074),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_997),
.B(n_847),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1074),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_992),
.B(n_929),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1124),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1019),
.A2(n_815),
.B1(n_840),
.B2(n_846),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1090),
.Y(n_1158)
);

AO22x2_ASAP7_75t_L g1159 ( 
.A1(n_1058),
.A2(n_815),
.B1(n_840),
.B2(n_846),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_978),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1002),
.B(n_934),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1090),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1010),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_994),
.B(n_990),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_982),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1064),
.Y(n_1166)
);

INVx8_ASAP7_75t_L g1167 ( 
.A(n_1013),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_981),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_SL g1169 ( 
.A(n_981),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_1060),
.A2(n_882),
.B1(n_862),
.B2(n_937),
.Y(n_1170)
);

BUFx8_ASAP7_75t_SL g1171 ( 
.A(n_1031),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1023),
.B(n_947),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_SL g1173 ( 
.A1(n_1075),
.A2(n_882),
.B1(n_961),
.B2(n_936),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_996),
.A2(n_972),
.B1(n_894),
.B2(n_859),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1069),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1090),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1016),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1040),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1093),
.B(n_893),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1070),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_977),
.Y(n_1181)
);

OAI22x1_ASAP7_75t_L g1182 ( 
.A1(n_1104),
.A2(n_944),
.B1(n_965),
.B2(n_935),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1093),
.B(n_920),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1093),
.B(n_920),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_982),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1027),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_987),
.A2(n_972),
.B1(n_894),
.B2(n_859),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_1025),
.Y(n_1188)
);

AND3x1_ASAP7_75t_SL g1189 ( 
.A(n_1006),
.B(n_27),
.C(n_29),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1005),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1031),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1005),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1054),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1033),
.B(n_958),
.Y(n_1194)
);

CKINVDCx11_ASAP7_75t_R g1195 ( 
.A(n_1075),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1097),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_977),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1008),
.A2(n_973),
.B1(n_958),
.B2(n_900),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_976),
.A2(n_973),
.B1(n_870),
.B2(n_939),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1016),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_980),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1039),
.B(n_798),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1014),
.A2(n_841),
.B1(n_877),
.B2(n_914),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1038),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1043),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_993),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_980),
.Y(n_1207)
);

AOI221x1_ASAP7_75t_L g1208 ( 
.A1(n_1051),
.A2(n_913),
.B1(n_901),
.B2(n_904),
.C(n_959),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_991),
.B(n_798),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1071),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1120),
.B(n_968),
.C(n_967),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_985),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1000),
.A2(n_888),
.B(n_886),
.C(n_885),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_985),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_976),
.A2(n_910),
.B1(n_952),
.B2(n_962),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1084),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1068),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1085),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1013),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1087),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1088),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1083),
.A2(n_955),
.B1(n_954),
.B2(n_792),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1106),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1089),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1007),
.A2(n_898),
.B1(n_808),
.B2(n_867),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1097),
.B(n_849),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1094),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_1038),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1121),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1102),
.A2(n_866),
.B1(n_848),
.B2(n_863),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1007),
.A2(n_808),
.B1(n_861),
.B2(n_891),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1107),
.B(n_1097),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1044),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1110),
.A2(n_790),
.B(n_806),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1052),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1051),
.B(n_890),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_SL g1237 ( 
.A1(n_1046),
.A2(n_857),
.B(n_888),
.C(n_886),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1025),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1096),
.B(n_849),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1025),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_988),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1121),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1052),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1103),
.B(n_863),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1065),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1112),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1101),
.A2(n_943),
.B1(n_946),
.B2(n_945),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1098),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1104),
.A2(n_877),
.B1(n_873),
.B2(n_876),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1065),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1100),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_988),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1013),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_989),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_989),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1034),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_986),
.A2(n_790),
.B(n_806),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_1118),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1003),
.A2(n_881),
.B(n_823),
.Y(n_1259)
);

AOI33xp33_ASAP7_75t_L g1260 ( 
.A1(n_1119),
.A2(n_29),
.A3(n_32),
.B1(n_33),
.B2(n_34),
.B3(n_35),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1012),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1127),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1122),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1012),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1126),
.B(n_943),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1058),
.A2(n_922),
.B1(n_914),
.B2(n_953),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1029),
.A2(n_922),
.B1(n_953),
.B2(n_926),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1122),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1015),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1015),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1065),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1129),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1065),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1086),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1049),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1072),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1017),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1017),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1018),
.A2(n_974),
.B(n_960),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1020),
.B(n_946),
.Y(n_1280)
);

INVx4_ASAP7_75t_L g1281 ( 
.A(n_1049),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1020),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1042),
.B(n_945),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1172),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1145),
.A2(n_1057),
.B(n_1118),
.C(n_1047),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1234),
.A2(n_1036),
.B(n_854),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1130),
.A2(n_1067),
.B1(n_1091),
.B2(n_1079),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1213),
.A2(n_1057),
.B(n_1047),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1173),
.A2(n_1059),
.B1(n_1123),
.B2(n_1081),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1163),
.B(n_1022),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1164),
.B(n_1073),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1173),
.A2(n_1053),
.B1(n_1123),
.B2(n_1048),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1208),
.A2(n_927),
.B(n_1113),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1131),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1248),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1234),
.A2(n_1099),
.B(n_1125),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1133),
.B(n_1281),
.Y(n_1297)
);

AOI221xp5_ASAP7_75t_L g1298 ( 
.A1(n_1157),
.A2(n_1006),
.B1(n_940),
.B2(n_911),
.C(n_926),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1174),
.A2(n_1062),
.B1(n_1095),
.B2(n_1078),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1148),
.A2(n_1099),
.B(n_1032),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1148),
.A2(n_1009),
.B(n_983),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1156),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1262),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1181),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1134),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1144),
.A2(n_960),
.B(n_974),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1190),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_SL g1308 ( 
.A1(n_1237),
.A2(n_911),
.B(n_1026),
.C(n_1046),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1135),
.Y(n_1309)
);

AO21x2_ASAP7_75t_L g1310 ( 
.A1(n_1209),
.A2(n_1202),
.B(n_1257),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1161),
.B(n_915),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1279),
.A2(n_1009),
.B(n_983),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1137),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1161),
.B(n_1049),
.Y(n_1314)
);

NOR2x1_ASAP7_75t_SL g1315 ( 
.A(n_1232),
.B(n_1122),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1281),
.B(n_1122),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1167),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1197),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1283),
.B(n_1142),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1139),
.A2(n_1111),
.B(n_1128),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1174),
.A2(n_1170),
.B1(n_1211),
.B2(n_1199),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1248),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1201),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1138),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1132),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1259),
.B(n_1062),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1279),
.A2(n_1009),
.B(n_983),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1140),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1139),
.A2(n_940),
.B(n_1114),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1260),
.A2(n_1266),
.B(n_1141),
.C(n_1143),
.Y(n_1330)
);

NOR2x1_ASAP7_75t_SL g1331 ( 
.A(n_1232),
.B(n_1062),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1171),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1143),
.A2(n_932),
.B1(n_1116),
.B2(n_1115),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1167),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1147),
.Y(n_1335)
);

NOR4xp25_ASAP7_75t_L g1336 ( 
.A(n_1274),
.B(n_1078),
.C(n_1022),
.D(n_1028),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1257),
.A2(n_999),
.B(n_1026),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1233),
.B(n_32),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1266),
.A2(n_1003),
.B(n_975),
.C(n_1115),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1191),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1280),
.A2(n_999),
.B(n_1026),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1253),
.B(n_1066),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1280),
.A2(n_1105),
.B(n_1116),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1253),
.B(n_1066),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1141),
.A2(n_1157),
.B(n_1170),
.C(n_1236),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1236),
.A2(n_1114),
.B(n_1105),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1187),
.A2(n_1003),
.B(n_975),
.C(n_1077),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1151),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1159),
.A2(n_1053),
.B1(n_1028),
.B2(n_1109),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1166),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1159),
.A2(n_1056),
.B1(n_1050),
.B2(n_1109),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1198),
.A2(n_1037),
.B(n_1076),
.Y(n_1352)
);

AO32x2_ASAP7_75t_L g1353 ( 
.A1(n_1198),
.A2(n_1056),
.A3(n_1037),
.B1(n_1108),
.B2(n_1092),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1163),
.B(n_36),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1175),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1209),
.A2(n_1050),
.B(n_1076),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1202),
.A2(n_1081),
.B(n_1048),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1238),
.A2(n_1045),
.B(n_1108),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1238),
.A2(n_1045),
.B(n_1041),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1192),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1240),
.A2(n_1041),
.B(n_1092),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_SL g1362 ( 
.A1(n_1239),
.A2(n_1117),
.B(n_1066),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1165),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1240),
.A2(n_960),
.B(n_974),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1155),
.A2(n_1114),
.B(n_932),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1180),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1258),
.A2(n_974),
.B(n_960),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1159),
.A2(n_1117),
.B1(n_1066),
.B2(n_1077),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1258),
.A2(n_1080),
.B(n_1077),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1192),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1182),
.A2(n_1268),
.B(n_1263),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1210),
.Y(n_1372)
);

AO31x2_ASAP7_75t_L g1373 ( 
.A1(n_1203),
.A2(n_1117),
.A3(n_1080),
.B(n_493),
.Y(n_1373)
);

INVx8_ASAP7_75t_L g1374 ( 
.A(n_1167),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1231),
.A2(n_1117),
.B(n_1080),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1231),
.A2(n_493),
.B(n_146),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1155),
.A2(n_493),
.B(n_206),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1251),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_L g1379 ( 
.A(n_1168),
.B(n_1185),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_SL g1380 ( 
.A1(n_1237),
.A2(n_36),
.B(n_38),
.C(n_40),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1263),
.A2(n_288),
.B(n_281),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1219),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1247),
.A2(n_280),
.B1(n_276),
.B2(n_275),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1244),
.A2(n_273),
.B(n_271),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_SL g1385 ( 
.A(n_1146),
.B(n_1204),
.Y(n_1385)
);

BUFx12f_ASAP7_75t_L g1386 ( 
.A(n_1150),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1192),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1177),
.Y(n_1388)
);

INVx4_ASAP7_75t_L g1389 ( 
.A(n_1200),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1189),
.A2(n_263),
.B1(n_258),
.B2(n_247),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1216),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1225),
.A2(n_119),
.B(n_151),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1225),
.A2(n_113),
.B(n_149),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1249),
.A2(n_100),
.B(n_145),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1203),
.A2(n_94),
.A3(n_141),
.B(n_129),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1249),
.A2(n_89),
.B(n_123),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1187),
.A2(n_1244),
.B(n_1222),
.C(n_1153),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1207),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1218),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1212),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1153),
.A2(n_246),
.B1(n_243),
.B2(n_233),
.Y(n_1401)
);

OAI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1194),
.A2(n_232),
.B1(n_229),
.B2(n_222),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1239),
.A2(n_72),
.B(n_86),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1230),
.A2(n_208),
.B(n_43),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1229),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1265),
.A2(n_57),
.B(n_66),
.Y(n_1406)
);

AOI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1268),
.A2(n_1194),
.B(n_1265),
.Y(n_1407)
);

OAI211xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1178),
.A2(n_1215),
.B(n_1189),
.C(n_1220),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1282),
.A2(n_74),
.B(n_83),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1214),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1221),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1278),
.A2(n_42),
.B(n_43),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1219),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1275),
.B(n_45),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_SL g1415 ( 
.A1(n_1136),
.A2(n_45),
.B(n_1149),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1178),
.A2(n_1186),
.B(n_1224),
.C(n_1227),
.Y(n_1416)
);

AOI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1246),
.A2(n_1272),
.B1(n_1223),
.B2(n_1205),
.C(n_1251),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1267),
.A2(n_1277),
.B(n_1270),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_SL g1419 ( 
.A1(n_1267),
.A2(n_1261),
.B(n_1241),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1252),
.A2(n_1254),
.B(n_1255),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1188),
.A2(n_1217),
.B(n_1193),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1169),
.A2(n_1232),
.B1(n_1219),
.B2(n_1158),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1264),
.A2(n_1269),
.B(n_1226),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1275),
.A2(n_1176),
.B(n_1158),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1162),
.A2(n_1196),
.B(n_1176),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1179),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1226),
.A2(n_1276),
.B(n_1184),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1245),
.Y(n_1428)
);

BUFx2_ASAP7_75t_SL g1429 ( 
.A(n_1169),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1229),
.Y(n_1430)
);

NAND2xp33_ASAP7_75t_R g1431 ( 
.A(n_1427),
.B(n_1183),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1360),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1345),
.A2(n_1162),
.B1(n_1196),
.B2(n_1206),
.Y(n_1433)
);

BUFx8_ASAP7_75t_SL g1434 ( 
.A(n_1332),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1321),
.A2(n_1256),
.B1(n_1195),
.B2(n_1160),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1408),
.A2(n_1160),
.B1(n_1152),
.B2(n_1154),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1290),
.B(n_1160),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1363),
.B(n_1229),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1408),
.A2(n_1152),
.B1(n_1154),
.B2(n_1242),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1345),
.A2(n_1188),
.B1(n_1243),
.B2(n_1235),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1302),
.Y(n_1441)
);

AOI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1377),
.A2(n_1184),
.B(n_1179),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1388),
.Y(n_1443)
);

NAND2x1p5_ASAP7_75t_L g1444 ( 
.A(n_1316),
.B(n_1188),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1291),
.B(n_1242),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1295),
.B(n_1242),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1289),
.A2(n_1152),
.B1(n_1154),
.B2(n_1183),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1317),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1325),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1295),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1377),
.A2(n_1245),
.B(n_1250),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1294),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1386),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1325),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1332),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1305),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1378),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1289),
.A2(n_1228),
.B1(n_1245),
.B2(n_1250),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1313),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1288),
.A2(n_1188),
.B(n_1250),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1309),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1324),
.Y(n_1462)
);

AOI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1330),
.A2(n_1397),
.B1(n_1404),
.B2(n_1287),
.C(n_1319),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1326),
.B(n_1427),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1340),
.B(n_1228),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1319),
.A2(n_1271),
.B1(n_1273),
.B2(n_1299),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1378),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1292),
.A2(n_1271),
.B1(n_1273),
.B2(n_1427),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1316),
.B(n_1271),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1360),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1322),
.B(n_1273),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1284),
.B(n_1354),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1292),
.A2(n_1311),
.B1(n_1368),
.B2(n_1383),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1373),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1328),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1340),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1368),
.A2(n_1349),
.B1(n_1298),
.B2(n_1401),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1349),
.A2(n_1401),
.B1(n_1351),
.B2(n_1417),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1335),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1421),
.B(n_1370),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1374),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_SL g1482 ( 
.A(n_1390),
.B(n_1416),
.C(n_1384),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1416),
.B(n_1397),
.C(n_1330),
.Y(n_1483)
);

AO31x2_ASAP7_75t_L g1484 ( 
.A1(n_1339),
.A2(n_1347),
.A3(n_1288),
.B(n_1400),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1348),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1350),
.Y(n_1486)
);

AOI221xp5_ASAP7_75t_L g1487 ( 
.A1(n_1380),
.A2(n_1285),
.B1(n_1402),
.B2(n_1347),
.C(n_1338),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1286),
.A2(n_1341),
.B(n_1343),
.Y(n_1488)
);

BUFx8_ASAP7_75t_L g1489 ( 
.A(n_1317),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1307),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1370),
.B(n_1387),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1309),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1355),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1366),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1376),
.A2(n_1306),
.B(n_1312),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1389),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1387),
.B(n_1405),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1405),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1314),
.B(n_1372),
.Y(n_1499)
);

AOI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1380),
.A2(n_1285),
.B1(n_1402),
.B2(n_1339),
.C(n_1333),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1391),
.B(n_1399),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1394),
.A2(n_1396),
.B(n_1306),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1411),
.B(n_1322),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1304),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1310),
.B(n_1336),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1326),
.B(n_1375),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1310),
.B(n_1333),
.Y(n_1507)
);

NAND2x1p5_ASAP7_75t_L g1508 ( 
.A(n_1422),
.B(n_1379),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1365),
.B(n_1430),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1326),
.B(n_1426),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1351),
.A2(n_1418),
.B1(n_1419),
.B2(n_1423),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1369),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1297),
.B(n_1426),
.Y(n_1513)
);

AND2x4_ASAP7_75t_SL g1514 ( 
.A(n_1389),
.B(n_1334),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1304),
.Y(n_1515)
);

BUFx5_ASAP7_75t_L g1516 ( 
.A(n_1342),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1317),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1369),
.Y(n_1518)
);

AND4x1_ASAP7_75t_L g1519 ( 
.A(n_1385),
.B(n_1414),
.C(n_1297),
.D(n_1346),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1423),
.A2(n_1329),
.B1(n_1318),
.B2(n_1410),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1318),
.Y(n_1521)
);

INVx4_ASAP7_75t_SL g1522 ( 
.A(n_1373),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_SL g1523 ( 
.A(n_1429),
.B(n_1374),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1407),
.B(n_1373),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1373),
.B(n_1426),
.Y(n_1525)
);

CKINVDCx11_ASAP7_75t_R g1526 ( 
.A(n_1303),
.Y(n_1526)
);

BUFx4f_ASAP7_75t_L g1527 ( 
.A(n_1317),
.Y(n_1527)
);

AOI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1293),
.A2(n_1392),
.B(n_1393),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1413),
.B(n_1382),
.Y(n_1529)
);

AO31x2_ASAP7_75t_L g1530 ( 
.A1(n_1323),
.A2(n_1398),
.A3(n_1400),
.B(n_1410),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1323),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1374),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1334),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1420),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1426),
.Y(n_1535)
);

AOI211xp5_ASAP7_75t_L g1536 ( 
.A1(n_1414),
.A2(n_1320),
.B(n_1308),
.C(n_1412),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1357),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1423),
.B(n_1293),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1420),
.A2(n_1293),
.B1(n_1382),
.B2(n_1356),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1352),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1382),
.A2(n_1415),
.B1(n_1413),
.B2(n_1344),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1331),
.B(n_1315),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1428),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1371),
.B(n_1361),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1428),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1342),
.B(n_1344),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1382),
.A2(n_1334),
.B1(n_1362),
.B2(n_1359),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1367),
.Y(n_1548)
);

AOI221x1_ASAP7_75t_SL g1549 ( 
.A1(n_1395),
.A2(n_1308),
.B1(n_1381),
.B2(n_1353),
.C(n_1403),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1353),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1463),
.A2(n_1483),
.B1(n_1482),
.B2(n_1433),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1490),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1463),
.A2(n_1334),
.B1(n_1395),
.B2(n_1424),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1472),
.B(n_1425),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1434),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1440),
.A2(n_1395),
.B1(n_1409),
.B2(n_1406),
.Y(n_1556)
);

CKINVDCx16_ASAP7_75t_R g1557 ( 
.A(n_1453),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1530),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1440),
.A2(n_1395),
.B(n_1353),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1454),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1445),
.B(n_1364),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1457),
.Y(n_1562)
);

NAND2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1481),
.B(n_1337),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1457),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1482),
.A2(n_1358),
.B1(n_1296),
.B2(n_1301),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1452),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1513),
.B(n_1327),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1456),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1470),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1443),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1501),
.B(n_1353),
.Y(n_1571)
);

AOI21xp33_ASAP7_75t_L g1572 ( 
.A1(n_1433),
.A2(n_1300),
.B(n_1505),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1487),
.A2(n_1500),
.B(n_1435),
.C(n_1536),
.Y(n_1573)
);

NAND2xp33_ASAP7_75t_R g1574 ( 
.A(n_1464),
.B(n_1506),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1476),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1448),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1491),
.Y(n_1577)
);

NOR3xp33_ASAP7_75t_SL g1578 ( 
.A(n_1455),
.B(n_1492),
.C(n_1496),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1477),
.A2(n_1478),
.B1(n_1487),
.B2(n_1466),
.Y(n_1579)
);

CKINVDCx16_ASAP7_75t_R g1580 ( 
.A(n_1461),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1499),
.B(n_1438),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1459),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_R g1583 ( 
.A(n_1523),
.B(n_1489),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1467),
.B(n_1450),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1480),
.B(n_1467),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1462),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1450),
.B(n_1446),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1480),
.B(n_1525),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_R g1589 ( 
.A(n_1523),
.B(n_1489),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1530),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1531),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_R g1592 ( 
.A(n_1464),
.B(n_1506),
.Y(n_1592)
);

OR2x6_ASAP7_75t_L g1593 ( 
.A(n_1464),
.B(n_1506),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1500),
.A2(n_1473),
.B1(n_1466),
.B2(n_1436),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1485),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1495),
.A2(n_1502),
.B(n_1442),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1503),
.B(n_1486),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1505),
.A2(n_1507),
.B(n_1524),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1519),
.B(n_1460),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_R g1600 ( 
.A(n_1526),
.B(n_1432),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_SL g1601 ( 
.A1(n_1465),
.A2(n_1471),
.B(n_1446),
.C(n_1460),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1438),
.B(n_1497),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1546),
.B(n_1432),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1508),
.B(n_1542),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1475),
.B(n_1479),
.Y(n_1605)
);

NOR2x1p5_ASAP7_75t_L g1606 ( 
.A(n_1481),
.B(n_1532),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1449),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1449),
.Y(n_1608)
);

NOR3xp33_ASAP7_75t_SL g1609 ( 
.A(n_1529),
.B(n_1502),
.C(n_1471),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1493),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1504),
.Y(n_1611)
);

NOR3xp33_ASAP7_75t_SL g1612 ( 
.A(n_1528),
.B(n_1507),
.C(n_1514),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1494),
.B(n_1437),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1498),
.B(n_1545),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1498),
.B(n_1516),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1535),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1515),
.Y(n_1617)
);

CKINVDCx16_ASAP7_75t_R g1618 ( 
.A(n_1431),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1521),
.Y(n_1619)
);

XOR2xp5_ASAP7_75t_L g1620 ( 
.A(n_1508),
.B(n_1509),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1543),
.Y(n_1621)
);

AO31x2_ASAP7_75t_L g1622 ( 
.A1(n_1524),
.A2(n_1534),
.A3(n_1538),
.B(n_1550),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1441),
.Y(n_1623)
);

AND2x4_ASAP7_75t_SL g1624 ( 
.A(n_1542),
.B(n_1510),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1593),
.B(n_1522),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1622),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1571),
.B(n_1522),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1622),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1622),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1558),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1567),
.B(n_1522),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1558),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1598),
.B(n_1474),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1598),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1622),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_1474),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1609),
.B(n_1488),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1562),
.B(n_1518),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1564),
.B(n_1518),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1566),
.Y(n_1640)
);

A2O1A1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1573),
.A2(n_1559),
.B(n_1551),
.C(n_1579),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1584),
.B(n_1538),
.Y(n_1642)
);

NAND3xp33_ASAP7_75t_L g1643 ( 
.A(n_1551),
.B(n_1439),
.C(n_1528),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1609),
.B(n_1549),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1568),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1554),
.B(n_1582),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1586),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1590),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1610),
.B(n_1488),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1590),
.Y(n_1650)
);

INVxp67_ASAP7_75t_R g1651 ( 
.A(n_1596),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1587),
.B(n_1549),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1569),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1617),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1585),
.B(n_1484),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1605),
.B(n_1484),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1597),
.B(n_1537),
.Y(n_1658)
);

BUFx3_ASAP7_75t_L g1659 ( 
.A(n_1604),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1611),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1611),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1619),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1603),
.B(n_1548),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1581),
.B(n_1484),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1593),
.B(n_1540),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1604),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1591),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1601),
.B(n_1512),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1577),
.B(n_1512),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1612),
.B(n_1561),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1612),
.B(n_1451),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_SL g1672 ( 
.A1(n_1641),
.A2(n_1599),
.B(n_1604),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1644),
.B(n_1600),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1653),
.B(n_1569),
.Y(n_1674)
);

OAI221xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1641),
.A2(n_1579),
.B1(n_1556),
.B2(n_1458),
.C(n_1541),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1670),
.B(n_1654),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1644),
.B(n_1599),
.C(n_1594),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1643),
.A2(n_1560),
.B1(n_1552),
.B2(n_1618),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1670),
.B(n_1602),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1653),
.B(n_1553),
.C(n_1572),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1643),
.A2(n_1607),
.B1(n_1620),
.B2(n_1615),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1670),
.B(n_1600),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1659),
.B(n_1624),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1642),
.B(n_1601),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1634),
.A2(n_1613),
.B1(n_1595),
.B2(n_1623),
.C(n_1565),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1654),
.B(n_1580),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1642),
.B(n_1614),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1654),
.B(n_1621),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1657),
.B(n_1608),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1654),
.B(n_1588),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1637),
.A2(n_1565),
.B1(n_1447),
.B2(n_1593),
.C(n_1511),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_SL g1692 ( 
.A1(n_1637),
.A2(n_1624),
.B(n_1589),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1634),
.B(n_1578),
.C(n_1616),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1657),
.B(n_1588),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1637),
.A2(n_1583),
.B1(n_1589),
.B2(n_1510),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1664),
.B(n_1583),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1668),
.A2(n_1563),
.B(n_1527),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1646),
.B(n_1576),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1671),
.A2(n_1576),
.B(n_1557),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1627),
.A2(n_1468),
.B1(n_1544),
.B2(n_1520),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1663),
.B(n_1578),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1633),
.B(n_1543),
.C(n_1547),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1668),
.A2(n_1539),
.B1(n_1592),
.B2(n_1574),
.C(n_1544),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1663),
.B(n_1576),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1646),
.B(n_1576),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1663),
.B(n_1516),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1646),
.B(n_1516),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1652),
.B(n_1664),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1638),
.B(n_1516),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1652),
.B(n_1664),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1652),
.B(n_1516),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_L g1712 ( 
.A(n_1649),
.B(n_1532),
.C(n_1533),
.D(n_1575),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1659),
.B(n_1555),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1659),
.B(n_1570),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1638),
.B(n_1516),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1708),
.B(n_1649),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1684),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1708),
.B(n_1649),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1687),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1689),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1680),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1710),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1710),
.B(n_1651),
.Y(n_1723)
);

NOR2x1_ASAP7_75t_SL g1724 ( 
.A(n_1682),
.B(n_1666),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1676),
.B(n_1651),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1676),
.B(n_1651),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1679),
.B(n_1671),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1679),
.B(n_1671),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1680),
.B(n_1658),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1709),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1715),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1706),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1701),
.B(n_1633),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1701),
.B(n_1633),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1674),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1706),
.B(n_1636),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1688),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1677),
.B(n_1675),
.C(n_1678),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1677),
.B(n_1645),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1704),
.B(n_1636),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1702),
.B(n_1658),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1702),
.B(n_1658),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1673),
.B(n_1640),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1688),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1704),
.B(n_1636),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1690),
.B(n_1711),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1694),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1690),
.B(n_1627),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1707),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1685),
.B(n_1645),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1711),
.B(n_1627),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1698),
.B(n_1647),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1705),
.B(n_1647),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1739),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1717),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1739),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1729),
.B(n_1639),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1724),
.B(n_1686),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1681),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1729),
.B(n_1719),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1721),
.B(n_1693),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1724),
.B(n_1699),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1719),
.B(n_1735),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1750),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1750),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1720),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1746),
.B(n_1713),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1720),
.B(n_1639),
.Y(n_1768)
);

BUFx2_ASAP7_75t_SL g1769 ( 
.A(n_1725),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1746),
.B(n_1693),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1735),
.B(n_1747),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1741),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1752),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1747),
.B(n_1645),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1722),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1743),
.B(n_1647),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1722),
.B(n_1696),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1752),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1752),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1722),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1753),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1741),
.B(n_1640),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1753),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1746),
.B(n_1714),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1753),
.Y(n_1785)
);

OAI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1738),
.A2(n_1672),
.B(n_1712),
.C(n_1692),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1742),
.B(n_1640),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1737),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1737),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1740),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1742),
.B(n_1655),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1744),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1730),
.B(n_1662),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1730),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1738),
.B(n_1712),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1755),
.B(n_1733),
.Y(n_1796)
);

NOR2xp67_ASAP7_75t_L g1797 ( 
.A(n_1786),
.B(n_1728),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1754),
.B(n_1733),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1762),
.B(n_1727),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1756),
.B(n_1733),
.Y(n_1800)
);

NOR2x1_ASAP7_75t_L g1801 ( 
.A(n_1761),
.B(n_1672),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1790),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1762),
.B(n_1727),
.Y(n_1803)
);

OAI32xp33_ASAP7_75t_L g1804 ( 
.A1(n_1795),
.A2(n_1734),
.A3(n_1726),
.B1(n_1725),
.B2(n_1727),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1764),
.A2(n_1703),
.B1(n_1723),
.B2(n_1725),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1761),
.A2(n_1691),
.B(n_1734),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1795),
.B(n_1734),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_SL g1808 ( 
.A(n_1758),
.B(n_1666),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1765),
.B(n_1716),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1772),
.B(n_1749),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1760),
.B(n_1771),
.Y(n_1811)
);

OAI31xp33_ASAP7_75t_L g1812 ( 
.A1(n_1759),
.A2(n_1728),
.A3(n_1726),
.B(n_1723),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1766),
.Y(n_1813)
);

AOI221xp5_ASAP7_75t_L g1814 ( 
.A1(n_1770),
.A2(n_1728),
.B1(n_1731),
.B2(n_1749),
.C(n_1723),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1769),
.B(n_1770),
.Y(n_1815)
);

AO221x1_ASAP7_75t_L g1816 ( 
.A1(n_1775),
.A2(n_1732),
.B1(n_1731),
.B2(n_1726),
.C(n_1629),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1777),
.A2(n_1695),
.B1(n_1732),
.B2(n_1683),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1763),
.B(n_1716),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1790),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1792),
.B(n_1716),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1788),
.B(n_1718),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1789),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1782),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1767),
.A2(n_1751),
.B1(n_1748),
.B2(n_1732),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1776),
.B(n_1718),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1767),
.B(n_1794),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1782),
.Y(n_1827)
);

NAND2x1p5_ASAP7_75t_L g1828 ( 
.A(n_1758),
.B(n_1683),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1787),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1777),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1830),
.B(n_1779),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1830),
.B(n_1784),
.Y(n_1832)
);

OAI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1806),
.A2(n_1757),
.B1(n_1787),
.B2(n_1791),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1815),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1807),
.B(n_1773),
.Y(n_1835)
);

NAND2x1_ASAP7_75t_L g1836 ( 
.A(n_1816),
.B(n_1777),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1815),
.B(n_1784),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1799),
.B(n_1778),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1813),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1828),
.B(n_1781),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1801),
.A2(n_1791),
.B(n_1780),
.Y(n_1841)
);

OAI332xp33_ASAP7_75t_L g1842 ( 
.A1(n_1817),
.A2(n_1785),
.A3(n_1783),
.B1(n_1768),
.B2(n_1780),
.B3(n_1774),
.C1(n_1793),
.C2(n_1635),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1806),
.A2(n_1797),
.B1(n_1805),
.B2(n_1808),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1822),
.Y(n_1844)
);

AOI222xp33_ASAP7_75t_L g1845 ( 
.A1(n_1814),
.A2(n_1626),
.B1(n_1628),
.B2(n_1629),
.C1(n_1635),
.C2(n_1775),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1823),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1799),
.B(n_1775),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1826),
.B(n_1768),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1803),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1827),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1803),
.B(n_1718),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1829),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1811),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1828),
.B(n_1748),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1796),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1849),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1849),
.Y(n_1857)
);

OAI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1843),
.A2(n_1812),
.B1(n_1810),
.B2(n_1809),
.C(n_1798),
.Y(n_1858)
);

O2A1O1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1833),
.A2(n_1804),
.B(n_1824),
.C(n_1800),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1834),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1837),
.B(n_1818),
.Y(n_1861)
);

OAI322xp33_ASAP7_75t_L g1862 ( 
.A1(n_1833),
.A2(n_1819),
.A3(n_1802),
.B1(n_1821),
.B2(n_1820),
.C1(n_1825),
.C2(n_1697),
.Y(n_1862)
);

OAI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1836),
.A2(n_1819),
.B1(n_1802),
.B2(n_1656),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1834),
.A2(n_1700),
.B1(n_1635),
.B2(n_1629),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1832),
.Y(n_1865)
);

OAI321xp33_ASAP7_75t_L g1866 ( 
.A1(n_1841),
.A2(n_1656),
.A3(n_1628),
.B1(n_1626),
.B2(n_1736),
.C(n_1740),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1844),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1832),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1832),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1839),
.Y(n_1870)
);

OAI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1845),
.A2(n_1628),
.B1(n_1626),
.B2(n_1736),
.C(n_1740),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1837),
.B(n_1745),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_SL g1873 ( 
.A(n_1853),
.B(n_1683),
.Y(n_1873)
);

AO22x1_ASAP7_75t_L g1874 ( 
.A1(n_1847),
.A2(n_1748),
.B1(n_1745),
.B2(n_1751),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1868),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1868),
.Y(n_1876)
);

OAI211xp5_ASAP7_75t_L g1877 ( 
.A1(n_1859),
.A2(n_1855),
.B(n_1854),
.C(n_1831),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1868),
.Y(n_1878)
);

INVxp67_ASAP7_75t_SL g1879 ( 
.A(n_1860),
.Y(n_1879)
);

AOI322xp5_ASAP7_75t_L g1880 ( 
.A1(n_1863),
.A2(n_1842),
.A3(n_1848),
.B1(n_1854),
.B2(n_1850),
.C1(n_1852),
.C2(n_1846),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1869),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1869),
.Y(n_1882)
);

OAI21xp5_ASAP7_75t_SL g1883 ( 
.A1(n_1863),
.A2(n_1840),
.B(n_1847),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1861),
.B(n_1838),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1865),
.B(n_1838),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1862),
.A2(n_1858),
.B(n_1867),
.C(n_1870),
.Y(n_1886)
);

AOI222xp33_ASAP7_75t_L g1887 ( 
.A1(n_1877),
.A2(n_1866),
.B1(n_1871),
.B2(n_1864),
.C1(n_1857),
.C2(n_1856),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1886),
.A2(n_1873),
.B(n_1874),
.Y(n_1888)
);

AOI221xp5_ASAP7_75t_L g1889 ( 
.A1(n_1883),
.A2(n_1881),
.B1(n_1880),
.B2(n_1882),
.C(n_1885),
.Y(n_1889)
);

OAI222xp33_ASAP7_75t_L g1890 ( 
.A1(n_1881),
.A2(n_1864),
.B1(n_1872),
.B2(n_1835),
.C1(n_1847),
.C2(n_1851),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1884),
.A2(n_1872),
.B1(n_1851),
.B2(n_1736),
.Y(n_1891)
);

NOR2x1_ASAP7_75t_L g1892 ( 
.A(n_1876),
.B(n_1745),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1885),
.Y(n_1893)
);

OAI21xp33_ASAP7_75t_L g1894 ( 
.A1(n_1884),
.A2(n_1751),
.B(n_1662),
.Y(n_1894)
);

NAND3xp33_ASAP7_75t_L g1895 ( 
.A(n_1875),
.B(n_1655),
.C(n_1662),
.Y(n_1895)
);

OAI211xp5_ASAP7_75t_L g1896 ( 
.A1(n_1879),
.A2(n_1533),
.B(n_1666),
.C(n_1659),
.Y(n_1896)
);

AOI22x1_ASAP7_75t_SL g1897 ( 
.A1(n_1893),
.A2(n_1876),
.B1(n_1878),
.B2(n_1889),
.Y(n_1897)
);

AOI211x1_ASAP7_75t_L g1898 ( 
.A1(n_1890),
.A2(n_1878),
.B(n_1655),
.C(n_1669),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1887),
.A2(n_1631),
.B1(n_1669),
.B2(n_1666),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1888),
.A2(n_1527),
.B(n_1448),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1892),
.B(n_1606),
.Y(n_1901)
);

OAI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1898),
.A2(n_1900),
.B(n_1899),
.C(n_1897),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1901),
.Y(n_1903)
);

O2A1O1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1897),
.A2(n_1896),
.B(n_1891),
.C(n_1894),
.Y(n_1904)
);

NOR4xp25_ASAP7_75t_L g1905 ( 
.A(n_1897),
.B(n_1895),
.C(n_1669),
.D(n_1661),
.Y(n_1905)
);

NOR4xp25_ASAP7_75t_L g1906 ( 
.A(n_1897),
.B(n_1660),
.C(n_1661),
.D(n_1631),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1900),
.B(n_1631),
.C(n_1661),
.Y(n_1907)
);

NAND4xp75_ASAP7_75t_L g1908 ( 
.A(n_1903),
.B(n_1451),
.C(n_1660),
.D(n_1661),
.Y(n_1908)
);

NOR3xp33_ASAP7_75t_L g1909 ( 
.A(n_1902),
.B(n_1660),
.C(n_1625),
.Y(n_1909)
);

NAND4xp75_ASAP7_75t_L g1910 ( 
.A(n_1906),
.B(n_1660),
.C(n_1632),
.D(n_1648),
.Y(n_1910)
);

NOR2x1_ASAP7_75t_L g1911 ( 
.A(n_1904),
.B(n_1905),
.Y(n_1911)
);

NOR3xp33_ASAP7_75t_L g1912 ( 
.A(n_1907),
.B(n_1625),
.C(n_1667),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1911),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1909),
.B(n_1448),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1910),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1913),
.A2(n_1912),
.B1(n_1908),
.B2(n_1517),
.Y(n_1916)
);

AOI221x1_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1915),
.B1(n_1914),
.B2(n_1517),
.C(n_1630),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1917),
.A2(n_1914),
.B1(n_1517),
.B2(n_1667),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1917),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1919),
.B(n_1667),
.Y(n_1920)
);

NOR3xp33_ASAP7_75t_SL g1921 ( 
.A(n_1918),
.B(n_1592),
.C(n_1574),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1920),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1921),
.A2(n_1667),
.B1(n_1625),
.B2(n_1630),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1922),
.A2(n_1625),
.B(n_1650),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1924),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1925),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1926),
.A2(n_1923),
.B1(n_1625),
.B2(n_1665),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1927),
.A2(n_1625),
.B1(n_1650),
.B2(n_1648),
.Y(n_1928)
);

AOI22xp33_ASAP7_75t_SL g1929 ( 
.A1(n_1928),
.A2(n_1444),
.B1(n_1469),
.B2(n_1665),
.Y(n_1929)
);

AOI211xp5_ASAP7_75t_L g1930 ( 
.A1(n_1929),
.A2(n_1665),
.B(n_1630),
.C(n_1632),
.Y(n_1930)
);


endmodule