module fake_jpeg_13779_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_1),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_47),
.B1(n_36),
.B2(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_67),
.B1(n_20),
.B2(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_42),
.CON(n_62),
.SN(n_62)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_56),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_18),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_74),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_62),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_61),
.C(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_71),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_41),
.C(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_2),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_3),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_6),
.B(n_7),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_6),
.B1(n_10),
.B2(n_13),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_4),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_24),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_87),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_94)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_87),
.B1(n_85),
.B2(n_26),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_101),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_82),
.B(n_84),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_92),
.C(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_104),
.C(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_100),
.B(n_97),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_107),
.B1(n_103),
.B2(n_102),
.Y(n_108)
);

AOI31xp67_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_96),
.A3(n_23),
.B(n_28),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_17),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_29),
.A3(n_30),
.B1(n_31),
.B2(n_32),
.C1(n_33),
.C2(n_35),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);


endmodule