module fake_jpeg_32172_n_527 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_527);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_60),
.Y(n_114)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_57),
.Y(n_164)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_59),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_0),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_66),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_17),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_70),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_31),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_2),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_74),
.B(n_76),
.Y(n_130)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_85),
.Y(n_140)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_18),
.B(n_2),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_18),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_101),
.B(n_20),
.Y(n_158)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_43),
.B1(n_47),
.B2(n_50),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_107),
.A2(n_131),
.B1(n_157),
.B2(n_57),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_58),
.A2(n_43),
.B1(n_29),
.B2(n_45),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_110),
.A2(n_25),
.B(n_21),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_37),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_85),
.B1(n_74),
.B2(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_47),
.B1(n_50),
.B2(n_45),
.Y(n_131)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_66),
.B(n_35),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_76),
.B(n_35),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_155),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_53),
.B(n_20),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_55),
.A2(n_47),
.B1(n_29),
.B2(n_26),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_37),
.Y(n_189)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_112),
.B(n_38),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_167),
.B(n_176),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_174),
.Y(n_220)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_126),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

INVx4_ASAP7_75t_SL g257 ( 
.A(n_173),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_140),
.C(n_130),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_177),
.A2(n_40),
.B1(n_42),
.B2(n_151),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_114),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_189),
.Y(n_222)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_138),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_181),
.B(n_182),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_119),
.A2(n_21),
.B(n_25),
.C(n_26),
.Y(n_182)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

NAND2x1p5_ASAP7_75t_L g188 ( 
.A(n_119),
.B(n_120),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_199),
.Y(n_243)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_191),
.Y(n_249)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_121),
.Y(n_193)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_120),
.B(n_39),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_218),
.Y(n_223)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_154),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_203),
.Y(n_227)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_108),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_130),
.B(n_68),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_206),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_155),
.B(n_28),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_202),
.A2(n_210),
.B(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_207),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_109),
.B1(n_118),
.B2(n_137),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_80),
.C(n_100),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_212),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_98),
.B1(n_163),
.B2(n_135),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_209),
.A2(n_211),
.B1(n_217),
.B2(n_144),
.Y(n_228)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_110),
.A2(n_23),
.B(n_28),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_139),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_214),
.Y(n_248)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_149),
.B(n_40),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_216),
.Y(n_247)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_118),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_123),
.B(n_39),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_229),
.B(n_236),
.Y(n_291)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_131),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_231),
.A2(n_182),
.B(n_206),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_173),
.A2(n_145),
.B1(n_160),
.B2(n_153),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_238),
.B1(n_243),
.B2(n_260),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_205),
.A2(n_217),
.B1(n_204),
.B2(n_199),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_234),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_175),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_242),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_177),
.A2(n_132),
.B1(n_128),
.B2(n_127),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_184),
.A2(n_116),
.B1(n_105),
.B2(n_115),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_239),
.B(n_142),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_134),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_201),
.A2(n_84),
.B1(n_72),
.B2(n_95),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_190),
.B1(n_170),
.B2(n_186),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_188),
.B(n_94),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_180),
.Y(n_281)
);

AO22x2_ASAP7_75t_L g258 ( 
.A1(n_209),
.A2(n_77),
.B1(n_78),
.B2(n_88),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_185),
.B1(n_169),
.B2(n_198),
.Y(n_296)
);

CKINVDCx9p33_ASAP7_75t_R g260 ( 
.A(n_187),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_260),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_261),
.Y(n_323)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_268),
.A2(n_293),
.B1(n_251),
.B2(n_245),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_223),
.B(n_222),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_272),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_270),
.A2(n_229),
.B(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_223),
.B(n_178),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_225),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_273),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_172),
.C(n_183),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_242),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_157),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_278),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g304 ( 
.A1(n_277),
.A2(n_285),
.B1(n_296),
.B2(n_239),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_230),
.B(n_166),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_227),
.B(n_200),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_280),
.B(n_286),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_287),
.Y(n_303)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_282),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_220),
.B(n_42),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_283),
.B(n_288),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_195),
.C(n_196),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_281),
.C(n_292),
.Y(n_313)
);

NAND2x1_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_214),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_237),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_221),
.B(n_192),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_187),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_208),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_243),
.B(n_255),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_329),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_275),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_231),
.B(n_236),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_306),
.A2(n_308),
.B(n_296),
.Y(n_352)
);

OAI32xp33_ASAP7_75t_L g307 ( 
.A1(n_274),
.A2(n_250),
.A3(n_254),
.B1(n_229),
.B2(n_258),
.Y(n_307)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_307),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_257),
.B(n_229),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_322),
.B(n_291),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_273),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_312),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_285),
.Y(n_332)
);

OAI22x1_ASAP7_75t_SL g315 ( 
.A1(n_291),
.A2(n_258),
.B1(n_257),
.B2(n_219),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_315),
.A2(n_316),
.B1(n_321),
.B2(n_328),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_276),
.A2(n_258),
.B1(n_219),
.B2(n_247),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_258),
.B1(n_219),
.B2(n_171),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_251),
.B(n_247),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_266),
.A2(n_290),
.B1(n_271),
.B2(n_286),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_326),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_265),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_274),
.A2(n_246),
.B1(n_253),
.B2(n_233),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_259),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_332),
.B(n_343),
.C(n_348),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_333),
.A2(n_345),
.B(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_337),
.B(n_352),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_283),
.Y(n_339)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_320),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_342),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_279),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_313),
.B(n_285),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_266),
.B(n_293),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_321),
.A2(n_293),
.B1(n_296),
.B2(n_268),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_347),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_277),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_320),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_349),
.Y(n_381)
);

OAI22x1_ASAP7_75t_SL g350 ( 
.A1(n_315),
.A2(n_296),
.B1(n_261),
.B2(n_253),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_353),
.B1(n_324),
.B2(n_322),
.Y(n_364)
);

OAI32xp33_ASAP7_75t_L g351 ( 
.A1(n_310),
.A2(n_315),
.A3(n_303),
.B1(n_318),
.B2(n_304),
.Y(n_351)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_316),
.A2(n_263),
.B1(n_264),
.B2(n_294),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_355),
.B(n_360),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_287),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_356),
.B(n_362),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_306),
.A2(n_261),
.B1(n_246),
.B2(n_245),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_357),
.A2(n_361),
.B1(n_323),
.B2(n_244),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_299),
.B(n_282),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_358),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_330),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_359),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_310),
.B(n_330),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_326),
.A2(n_225),
.B1(n_241),
.B2(n_244),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_267),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_364),
.A2(n_367),
.B1(n_377),
.B2(n_395),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_334),
.A2(n_303),
.B1(n_307),
.B2(n_311),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_344),
.A2(n_304),
.B1(n_319),
.B2(n_328),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_386),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_319),
.C(n_304),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_378),
.C(n_370),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_344),
.A2(n_298),
.B1(n_304),
.B2(n_309),
.Y(n_376)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_334),
.A2(n_298),
.B1(n_309),
.B2(n_300),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_300),
.C(n_312),
.Y(n_378)
);

AOI22x1_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_325),
.B1(n_317),
.B2(n_297),
.Y(n_384)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_384),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_325),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_335),
.B(n_317),
.Y(n_388)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_388),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_331),
.A2(n_323),
.B1(n_297),
.B2(n_241),
.Y(n_390)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_391),
.A2(n_347),
.B1(n_354),
.B2(n_355),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_346),
.B(n_262),
.Y(n_392)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_392),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_333),
.A2(n_211),
.B(n_32),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_393),
.B(n_340),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_3),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_336),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_331),
.A2(n_47),
.B1(n_32),
.B2(n_5),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_363),
.Y(n_396)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_396),
.Y(n_425)
);

AOI221xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_351),
.B1(n_366),
.B2(n_385),
.C(n_367),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_417),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_401),
.Y(n_428)
);

A2O1A1O1Ixp25_ASAP7_75t_L g401 ( 
.A1(n_366),
.A2(n_363),
.B(n_352),
.C(n_348),
.D(n_337),
.Y(n_401)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_383),
.A2(n_340),
.B1(n_357),
.B2(n_361),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_405),
.A2(n_391),
.B1(n_384),
.B2(n_369),
.Y(n_433)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_406),
.A2(n_393),
.B(n_373),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_362),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_409),
.B(n_410),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_380),
.B(n_356),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_353),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_411),
.B(n_365),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_412),
.A2(n_383),
.B1(n_395),
.B2(n_379),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_371),
.B(n_3),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_420),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_47),
.C(n_19),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_419),
.C(n_368),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_19),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_3),
.Y(n_418)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_418),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_365),
.B(n_19),
.C(n_4),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_372),
.B(n_3),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_421),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_392),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_422),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_4),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_394),
.Y(n_426)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_407),
.A2(n_384),
.B1(n_374),
.B2(n_386),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_437),
.Y(n_452)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_430),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_407),
.A2(n_382),
.B1(n_388),
.B2(n_387),
.Y(n_435)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_402),
.A2(n_386),
.B1(n_368),
.B2(n_382),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_446),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_412),
.A2(n_403),
.B1(n_413),
.B2(n_414),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_443),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_386),
.Y(n_441)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_441),
.Y(n_456)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_414),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_434),
.B(n_399),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_447),
.B(n_444),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_411),
.C(n_417),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_454),
.C(n_458),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_400),
.C(n_416),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_400),
.B(n_403),
.C(n_413),
.Y(n_457)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_398),
.C(n_413),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_398),
.C(n_405),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_465),
.C(n_430),
.Y(n_480)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_419),
.C(n_401),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_SL g467 ( 
.A(n_461),
.B(n_438),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_467),
.A2(n_451),
.B1(n_456),
.B2(n_427),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_425),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_472),
.Y(n_484)
);

FAx1_ASAP7_75t_SL g469 ( 
.A(n_454),
.B(n_440),
.CI(n_429),
.CON(n_469),
.SN(n_469)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_459),
.B(n_437),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_471),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_439),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_448),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_476),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_431),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_478),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_452),
.B(n_426),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_465),
.A2(n_443),
.B(n_442),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_477),
.A2(n_457),
.B(n_462),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_424),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_480),
.B(n_481),
.Y(n_485)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_464),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_427),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_455),
.C(n_450),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_483),
.B(n_487),
.Y(n_501)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_486),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_480),
.A2(n_455),
.B(n_463),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_490),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_473),
.A2(n_450),
.B1(n_463),
.B2(n_456),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_489),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_445),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_471),
.A2(n_459),
.B(n_6),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_491),
.A2(n_484),
.B(n_493),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_4),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_6),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_478),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_9),
.Y(n_506)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_498),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g499 ( 
.A(n_494),
.B(n_475),
.C(n_470),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_486),
.B(n_491),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_466),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_502),
.B(n_503),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_466),
.C(n_19),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_508),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_492),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_505),
.B(n_506),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_501),
.A2(n_485),
.B(n_497),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_511),
.A2(n_498),
.B(n_496),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_507),
.B(n_488),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_10),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_514),
.A2(n_500),
.B(n_499),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_516),
.Y(n_521)
);

AOI21xp33_ASAP7_75t_L g520 ( 
.A1(n_517),
.A2(n_518),
.B(n_519),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_510),
.A2(n_10),
.B(n_13),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_521),
.B(n_515),
.C(n_509),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_520),
.B(n_513),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_14),
.C(n_15),
.Y(n_524)
);

MAJx2_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_14),
.C(n_15),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_525),
.B(n_15),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_16),
.B(n_19),
.Y(n_527)
);


endmodule