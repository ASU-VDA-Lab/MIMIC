module fake_jpeg_29453_n_44 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_44);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_3),
.B1(n_5),
.B2(n_22),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_28),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_23),
.B1(n_35),
.B2(n_15),
.Y(n_41)
);

A2O1A1O1Ixp25_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_15),
.B(n_29),
.C(n_13),
.D(n_28),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_36),
.B(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.C(n_16),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_13),
.C(n_23),
.Y(n_44)
);


endmodule