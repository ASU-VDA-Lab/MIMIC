module fake_netlist_6_2380_n_1414 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_340, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1414);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1414;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1309;
wire n_1123;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_474;
wire n_1207;
wire n_1368;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1362;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g342 ( 
.A(n_28),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_254),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_51),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_135),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_108),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_217),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_49),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_52),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_27),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_172),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_327),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_109),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_95),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_18),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_72),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_330),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_154),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_120),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_67),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_232),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_128),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_335),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_273),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_306),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_224),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_191),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_153),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_9),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_99),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_183),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_17),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_200),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_11),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_41),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_144),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_313),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_9),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_325),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_309),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_105),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_298),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_15),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_287),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_28),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_43),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_220),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_80),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_6),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_12),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_16),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_115),
.Y(n_394)
);

BUFx10_ASAP7_75t_L g395 ( 
.A(n_107),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_20),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_307),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_6),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_241),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_138),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_188),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_219),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_274),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_234),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_34),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_73),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_302),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_315),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_85),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_0),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_291),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_271),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_110),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_211),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_129),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_238),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_213),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_146),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_123),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_151),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_53),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_323),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_55),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_26),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_156),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_164),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_68),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_303),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_324),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_155),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_103),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_339),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_82),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_29),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_190),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_244),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_331),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_35),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_215),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_161),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_338),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_296),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_39),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_280),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_253),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_264),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_314),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_310),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_236),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_24),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_35),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_30),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_160),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_83),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_255),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_93),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_5),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_305),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_60),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_133),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_50),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_148),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_165),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_12),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_185),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_276),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_312),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_221),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_205),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_13),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_30),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_304),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_64),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_84),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_311),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_289),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_136),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_184),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_114),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_260),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_119),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_61),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_157),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_270),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_89),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_125),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_252),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_229),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_38),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_262),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_333),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_139),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_266),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_301),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_269),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_17),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_23),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_158),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_34),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_130),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_209),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_26),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_113),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_228),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_237),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_91),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_181),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_300),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_169),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_75),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_235),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_170),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_201),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_197),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_24),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_149),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_222),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_32),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_46),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_23),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_308),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_78),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_134),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_230),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_207),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_116),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_147),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_286),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_212),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_39),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_46),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_299),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_444),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_405),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_376),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_345),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_343),
.B(n_0),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_347),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_376),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_349),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_531),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_519),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_453),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_531),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_351),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_405),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_R g548 ( 
.A(n_348),
.B(n_1),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_374),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_377),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_405),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_405),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_342),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_356),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_371),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_353),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_380),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_385),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_387),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_391),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_388),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_354),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_357),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_392),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_393),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_358),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_398),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_359),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_361),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_362),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_410),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_396),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_343),
.B(n_1),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_364),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_367),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_368),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_426),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_451),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_425),
.Y(n_579)
);

NOR2xp67_ASAP7_75t_L g580 ( 
.A(n_520),
.B(n_2),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_465),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_484),
.B(n_2),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_435),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_370),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_373),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_498),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_426),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_452),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_439),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_344),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_346),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_350),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_352),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_488),
.B(n_3),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_369),
.B(n_401),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_355),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_378),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_360),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_363),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_412),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_458),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_379),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_407),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_407),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_382),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_365),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_383),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_471),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_372),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_490),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_500),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_375),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_386),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_389),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_390),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_468),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_L g619 ( 
.A(n_462),
.B(n_3),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_397),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_394),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_399),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_503),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_403),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_406),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_414),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_516),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_415),
.Y(n_628)
);

INVxp33_ASAP7_75t_SL g629 ( 
.A(n_521),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_417),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_418),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_366),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_400),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_402),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_420),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_546),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_535),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_547),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_535),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_546),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_551),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_552),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_551),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_590),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_557),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_534),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_559),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_557),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_564),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_610),
.B(n_623),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_564),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_592),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_577),
.B(n_432),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_593),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_594),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_595),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_597),
.B(n_441),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_573),
.B(n_508),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_598),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_600),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_601),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_608),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_611),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_537),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_614),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_578),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_615),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_577),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_550),
.Y(n_670)
);

OA21x2_ASAP7_75t_L g671 ( 
.A1(n_617),
.A2(n_462),
.B(n_429),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_620),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_596),
.B(n_413),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_577),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_624),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_553),
.Y(n_676)
);

AND2x2_ASAP7_75t_SL g677 ( 
.A(n_538),
.B(n_413),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_626),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_628),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_560),
.B(n_395),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_630),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_631),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_635),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_554),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_555),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_565),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_603),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_558),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_567),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_571),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_605),
.B(n_424),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_R g692 ( 
.A(n_549),
.B(n_532),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_579),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_581),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_582),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_584),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_588),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_536),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_540),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_589),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_542),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_545),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_583),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_625),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_634),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_539),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_561),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_602),
.A2(n_384),
.B1(n_436),
.B2(n_381),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_541),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_556),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_606),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_619),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_591),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_580),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_612),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_613),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_576),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_618),
.B(n_413),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_549),
.Y(n_719)
);

AND2x6_ASAP7_75t_L g720 ( 
.A(n_658),
.B(n_413),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_704),
.B(n_445),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_706),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_698),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_644),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_703),
.B(n_562),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_703),
.B(n_563),
.Y(n_726)
);

AND2x6_ASAP7_75t_L g727 ( 
.A(n_658),
.B(n_475),
.Y(n_727)
);

CKINVDCx8_ASAP7_75t_R g728 ( 
.A(n_706),
.Y(n_728)
);

AND2x6_ASAP7_75t_L g729 ( 
.A(n_653),
.B(n_475),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_703),
.B(n_566),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_638),
.Y(n_731)
);

NAND2x1p5_ASAP7_75t_L g732 ( 
.A(n_706),
.B(n_475),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_648),
.Y(n_733)
);

INVx5_ASAP7_75t_L g734 ( 
.A(n_718),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_677),
.A2(n_692),
.B1(n_650),
.B2(n_686),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_648),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_677),
.B(n_568),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_644),
.B(n_569),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_704),
.B(n_570),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_669),
.B(n_674),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_669),
.B(n_574),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_713),
.B(n_544),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_669),
.B(n_575),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_684),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_703),
.B(n_586),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_706),
.B(n_587),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_719),
.B(n_599),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_648),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_648),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_647),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_685),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_651),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_669),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_674),
.B(n_657),
.Y(n_754)
);

INVx4_ASAP7_75t_SL g755 ( 
.A(n_718),
.Y(n_755)
);

INVx4_ASAP7_75t_SL g756 ( 
.A(n_718),
.Y(n_756)
);

OR2x2_ASAP7_75t_SL g757 ( 
.A(n_647),
.B(n_632),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_651),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_711),
.B(n_482),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_705),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_651),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_651),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_674),
.B(n_604),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_711),
.B(n_483),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_680),
.B(n_607),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_693),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_646),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_705),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_694),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_692),
.A2(n_629),
.B1(n_616),
.B2(n_621),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_701),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_700),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_674),
.B(n_609),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_695),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_717),
.B(n_622),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_653),
.B(n_504),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_696),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_646),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_713),
.B(n_633),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_700),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_641),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_701),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_650),
.B(n_629),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_657),
.B(n_404),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_691),
.A2(n_511),
.B1(n_525),
.B2(n_475),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_691),
.A2(n_525),
.B1(n_526),
.B2(n_511),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_697),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_665),
.B(n_550),
.Y(n_788)
);

NAND2x1p5_ASAP7_75t_L g789 ( 
.A(n_709),
.B(n_511),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_642),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_718),
.B(n_673),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_718),
.B(n_408),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_652),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_665),
.B(n_572),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_673),
.B(n_700),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_700),
.B(n_643),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_687),
.B(n_428),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_709),
.B(n_511),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_654),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_641),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_710),
.B(n_548),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_686),
.B(n_572),
.Y(n_802)
);

NAND2x1p5_ASAP7_75t_L g803 ( 
.A(n_710),
.B(n_525),
.Y(n_803)
);

INVx5_ASAP7_75t_L g804 ( 
.A(n_701),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_641),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_655),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_641),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_687),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_656),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_754),
.B(n_716),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_731),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_731),
.Y(n_812)
);

NAND2x1p5_ASAP7_75t_L g813 ( 
.A(n_722),
.B(n_690),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_737),
.A2(n_715),
.B1(n_708),
.B2(n_473),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_790),
.Y(n_815)
);

AO22x2_ASAP7_75t_L g816 ( 
.A1(n_724),
.A2(n_543),
.B1(n_534),
.B2(n_707),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_790),
.Y(n_817)
);

CKINVDCx14_ASAP7_75t_R g818 ( 
.A(n_788),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_722),
.B(n_690),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_753),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_760),
.B(n_699),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_739),
.B(n_671),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_738),
.B(n_712),
.Y(n_823)
);

AO22x2_ASAP7_75t_L g824 ( 
.A1(n_797),
.A2(n_714),
.B1(n_431),
.B2(n_443),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_768),
.B(n_702),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_744),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_728),
.Y(n_827)
);

AO22x2_ASAP7_75t_L g828 ( 
.A1(n_783),
.A2(n_437),
.B1(n_455),
.B2(n_449),
.Y(n_828)
);

AO22x2_ASAP7_75t_L g829 ( 
.A1(n_776),
.A2(n_543),
.B1(n_456),
.B2(n_485),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_767),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_753),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_735),
.A2(n_627),
.B1(n_585),
.B2(n_659),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_802),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_751),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_766),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_808),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_769),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_753),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_778),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_774),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_777),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_808),
.B(n_636),
.Y(n_842)
);

AO22x2_ASAP7_75t_L g843 ( 
.A1(n_776),
.A2(n_476),
.B1(n_489),
.B2(n_486),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_787),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_793),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_742),
.B(n_640),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_799),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_750),
.B(n_670),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_806),
.Y(n_849)
);

NAND2x1p5_ASAP7_75t_L g850 ( 
.A(n_734),
.B(n_660),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_809),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_772),
.Y(n_852)
);

BUFx8_ASAP7_75t_L g853 ( 
.A(n_779),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_723),
.Y(n_854)
);

AO22x2_ASAP7_75t_L g855 ( 
.A1(n_759),
.A2(n_764),
.B1(n_801),
.B2(n_721),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_796),
.Y(n_856)
);

BUFx8_ASAP7_75t_L g857 ( 
.A(n_765),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_721),
.A2(n_501),
.B1(n_515),
.B2(n_427),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_759),
.B(n_661),
.Y(n_859)
);

OAI221xp5_ASAP7_75t_L g860 ( 
.A1(n_784),
.A2(n_786),
.B1(n_785),
.B2(n_666),
.C(n_668),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_775),
.A2(n_627),
.B1(n_585),
.B2(n_662),
.Y(n_861)
);

AO22x2_ASAP7_75t_L g862 ( 
.A1(n_764),
.A2(n_492),
.B1(n_493),
.B2(n_491),
.Y(n_862)
);

AO21x1_ASAP7_75t_L g863 ( 
.A1(n_791),
.A2(n_505),
.B(n_502),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_740),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_794),
.Y(n_865)
);

CKINVDCx16_ASAP7_75t_R g866 ( 
.A(n_770),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_734),
.B(n_664),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_747),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_805),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_795),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_748),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_734),
.B(n_548),
.Y(n_872)
);

AO22x2_ASAP7_75t_L g873 ( 
.A1(n_725),
.A2(n_507),
.B1(n_514),
.B2(n_506),
.Y(n_873)
);

AO22x2_ASAP7_75t_L g874 ( 
.A1(n_726),
.A2(n_522),
.B1(n_523),
.B2(n_518),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_746),
.B(n_672),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_730),
.Y(n_876)
);

AO22x2_ASAP7_75t_L g877 ( 
.A1(n_745),
.A2(n_527),
.B1(n_529),
.B2(n_524),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_749),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_741),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_743),
.A2(n_678),
.B1(n_679),
.B2(n_675),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_763),
.B(n_681),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_773),
.B(n_682),
.Y(n_882)
);

AO22x2_ASAP7_75t_L g883 ( 
.A1(n_757),
.A2(n_533),
.B1(n_7),
.B2(n_4),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_752),
.Y(n_884)
);

AO22x2_ASAP7_75t_L g885 ( 
.A1(n_755),
.A2(n_683),
.B1(n_7),
.B2(n_4),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_758),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_792),
.B(n_701),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_729),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_761),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_805),
.Y(n_890)
);

AO22x2_ASAP7_75t_L g891 ( 
.A1(n_755),
.A2(n_10),
.B1(n_5),
.B2(n_8),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_781),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_800),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_771),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_789),
.B(n_676),
.Y(n_895)
);

AO22x2_ASAP7_75t_L g896 ( 
.A1(n_756),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_896)
);

OAI22xp33_ASAP7_75t_L g897 ( 
.A1(n_803),
.A2(n_689),
.B1(n_688),
.B2(n_667),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_780),
.B(n_649),
.Y(n_898)
);

BUFx8_ASAP7_75t_L g899 ( 
.A(n_729),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_732),
.A2(n_416),
.B1(n_419),
.B2(n_411),
.Y(n_900)
);

OAI221xp5_ASAP7_75t_L g901 ( 
.A1(n_782),
.A2(n_645),
.B1(n_663),
.B2(n_649),
.C(n_671),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_733),
.Y(n_902)
);

AO22x2_ASAP7_75t_L g903 ( 
.A1(n_756),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_903)
);

NAND2xp33_ASAP7_75t_SL g904 ( 
.A(n_827),
.B(n_421),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_821),
.B(n_825),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_868),
.B(n_780),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_881),
.B(n_805),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_876),
.B(n_807),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_879),
.B(n_807),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_865),
.B(n_807),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_882),
.B(n_804),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_823),
.B(n_663),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_SL g913 ( 
.A(n_814),
.B(n_422),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_SL g914 ( 
.A(n_810),
.B(n_423),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_870),
.B(n_720),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_856),
.B(n_720),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_833),
.B(n_804),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_861),
.B(n_804),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_836),
.B(n_729),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_859),
.B(n_736),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_818),
.B(n_395),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_811),
.B(n_762),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_812),
.B(n_430),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_815),
.B(n_433),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_817),
.B(n_434),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_832),
.B(n_438),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_840),
.B(n_440),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_864),
.B(n_720),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_864),
.B(n_727),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_826),
.B(n_727),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_834),
.B(n_727),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_SL g932 ( 
.A(n_888),
.B(n_442),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_844),
.B(n_798),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_835),
.B(n_446),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_837),
.B(n_841),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_845),
.B(n_447),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_855),
.B(n_409),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_847),
.B(n_448),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_849),
.B(n_798),
.Y(n_939)
);

NAND2xp33_ASAP7_75t_SL g940 ( 
.A(n_872),
.B(n_450),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_851),
.B(n_798),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_854),
.B(n_454),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_822),
.B(n_457),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_852),
.B(n_459),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_880),
.B(n_460),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_887),
.B(n_461),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_873),
.B(n_463),
.Y(n_947)
);

AND2x2_ASAP7_75t_SL g948 ( 
.A(n_866),
.B(n_525),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_846),
.B(n_875),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_873),
.B(n_464),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_848),
.B(n_466),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_813),
.B(n_467),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_874),
.B(n_469),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_830),
.B(n_470),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_819),
.B(n_474),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_894),
.B(n_637),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_895),
.B(n_897),
.Y(n_957)
);

NAND2xp33_ASAP7_75t_SL g958 ( 
.A(n_839),
.B(n_858),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_874),
.B(n_477),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_902),
.B(n_478),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_853),
.B(n_479),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_899),
.B(n_820),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_877),
.B(n_480),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_831),
.B(n_838),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_869),
.B(n_481),
.Y(n_965)
);

NAND2xp33_ASAP7_75t_SL g966 ( 
.A(n_890),
.B(n_487),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_SL g967 ( 
.A(n_900),
.B(n_494),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_857),
.B(n_495),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_863),
.B(n_496),
.Y(n_969)
);

NAND2xp33_ASAP7_75t_SL g970 ( 
.A(n_871),
.B(n_499),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_878),
.B(n_509),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_SL g972 ( 
.A(n_884),
.B(n_510),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_886),
.B(n_512),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_889),
.B(n_513),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_892),
.B(n_517),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_913),
.A2(n_860),
.B(n_893),
.C(n_901),
.Y(n_976)
);

OA21x2_ASAP7_75t_L g977 ( 
.A1(n_943),
.A2(n_639),
.B(n_637),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_905),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_912),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_935),
.B(n_828),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_915),
.A2(n_898),
.B(n_867),
.Y(n_981)
);

OA21x2_ASAP7_75t_L g982 ( 
.A1(n_969),
.A2(n_639),
.B(n_530),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_905),
.B(n_842),
.Y(n_983)
);

AO21x2_ASAP7_75t_L g984 ( 
.A1(n_957),
.A2(n_877),
.B(n_828),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_SL g985 ( 
.A(n_948),
.B(n_842),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_916),
.A2(n_862),
.B(n_528),
.C(n_526),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_958),
.A2(n_862),
.B(n_528),
.C(n_526),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_911),
.A2(n_843),
.B(n_885),
.Y(n_988)
);

CKINVDCx8_ASAP7_75t_R g989 ( 
.A(n_956),
.Y(n_989)
);

AO32x2_ASAP7_75t_L g990 ( 
.A1(n_948),
.A2(n_824),
.A3(n_885),
.B1(n_891),
.B2(n_896),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_946),
.B(n_824),
.Y(n_991)
);

BUFx2_ASAP7_75t_R g992 ( 
.A(n_962),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_928),
.A2(n_850),
.B(n_891),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_929),
.A2(n_896),
.B(n_528),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_930),
.A2(n_903),
.B(n_883),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_964),
.A2(n_48),
.B(n_47),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_921),
.B(n_829),
.Y(n_997)
);

OA21x2_ASAP7_75t_L g998 ( 
.A1(n_931),
.A2(n_528),
.B(n_526),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_956),
.Y(n_999)
);

NAND2x1p5_ASAP7_75t_L g1000 ( 
.A(n_907),
.B(n_816),
.Y(n_1000)
);

O2A1O1Ixp5_ASAP7_75t_SL g1001 ( 
.A1(n_918),
.A2(n_409),
.B(n_16),
.C(n_18),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_920),
.B(n_54),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_906),
.B(n_14),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_922),
.A2(n_57),
.B(n_56),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_939),
.A2(n_59),
.B(n_58),
.Y(n_1005)
);

BUFx10_ASAP7_75t_L g1006 ( 
.A(n_933),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_952),
.A2(n_63),
.B(n_62),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_909),
.A2(n_66),
.B(n_65),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_941),
.A2(n_70),
.B(n_69),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_919),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_955),
.A2(n_74),
.B(n_71),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_908),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_965),
.A2(n_77),
.B(n_76),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_947),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_1014)
);

OA21x2_ASAP7_75t_L g1015 ( 
.A1(n_950),
.A2(n_81),
.B(n_79),
.Y(n_1015)
);

NAND3xp33_ASAP7_75t_L g1016 ( 
.A(n_926),
.B(n_19),
.C(n_21),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_944),
.A2(n_87),
.B(n_86),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_949),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_910),
.A2(n_90),
.B(n_88),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_970),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_933),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_953),
.A2(n_22),
.B(n_25),
.C(n_27),
.Y(n_1022)
);

AO31x2_ASAP7_75t_L g1023 ( 
.A1(n_959),
.A2(n_22),
.A3(n_25),
.B(n_29),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_960),
.A2(n_94),
.B(n_92),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_951),
.B(n_31),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_971),
.A2(n_97),
.B(n_96),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_975),
.A2(n_100),
.B(n_98),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_973),
.Y(n_1028)
);

O2A1O1Ixp5_ASAP7_75t_L g1029 ( 
.A1(n_923),
.A2(n_216),
.B(n_340),
.C(n_337),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_974),
.A2(n_102),
.B(n_101),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_917),
.A2(n_925),
.B(n_924),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_927),
.A2(n_106),
.B(n_104),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_934),
.A2(n_938),
.B(n_936),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_937),
.B(n_942),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_963),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_985),
.B(n_904),
.Y(n_1036)
);

OAI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_979),
.A2(n_968),
.B1(n_961),
.B2(n_945),
.Y(n_1037)
);

INVx5_ASAP7_75t_L g1038 ( 
.A(n_1006),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_979),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_996),
.A2(n_966),
.B(n_972),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_976),
.A2(n_914),
.B(n_967),
.Y(n_1041)
);

NAND2x1p5_ASAP7_75t_L g1042 ( 
.A(n_1018),
.B(n_932),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_1004),
.A2(n_940),
.B(n_954),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1012),
.Y(n_1044)
);

AO21x2_ASAP7_75t_L g1045 ( 
.A1(n_986),
.A2(n_987),
.B(n_1005),
.Y(n_1045)
);

AOI21xp33_ASAP7_75t_SL g1046 ( 
.A1(n_1000),
.A2(n_31),
.B(n_32),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_991),
.B(n_33),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1034),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_SL g1049 ( 
.A1(n_981),
.A2(n_225),
.B(n_336),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_1028),
.B(n_341),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_983),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1021),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1016),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1021),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1035),
.B(n_40),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_989),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_1006),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_980),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_984),
.A2(n_1025),
.B1(n_1034),
.B2(n_994),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1010),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_999),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1003),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1008),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_1009),
.A2(n_226),
.B(n_332),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_1019),
.A2(n_223),
.B(n_329),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_1013),
.A2(n_218),
.B(n_322),
.Y(n_1066)
);

OA21x2_ASAP7_75t_L g1067 ( 
.A1(n_1031),
.A2(n_214),
.B(n_321),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_978),
.B(n_334),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1002),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_983),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_984),
.B(n_1028),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_978),
.Y(n_1072)
);

OAI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_995),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_1032),
.A2(n_227),
.B(n_319),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1002),
.Y(n_1075)
);

AO21x1_ASAP7_75t_L g1076 ( 
.A1(n_993),
.A2(n_42),
.B(n_43),
.Y(n_1076)
);

INVx6_ASAP7_75t_L g1077 ( 
.A(n_978),
.Y(n_1077)
);

INVx4_ASAP7_75t_SL g1078 ( 
.A(n_1023),
.Y(n_1078)
);

BUFx12f_ASAP7_75t_L g1079 ( 
.A(n_1020),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1022),
.A2(n_44),
.B1(n_45),
.B2(n_111),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_997),
.B(n_112),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1026),
.A2(n_233),
.B(n_318),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1033),
.B(n_44),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1027),
.A2(n_1030),
.B(n_1024),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_990),
.B(n_45),
.Y(n_1085)
);

BUFx2_ASAP7_75t_SL g1086 ( 
.A(n_982),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_977),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_977),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_988),
.B(n_117),
.Y(n_1089)
);

AOI21x1_ASAP7_75t_L g1090 ( 
.A1(n_982),
.A2(n_320),
.B(n_121),
.Y(n_1090)
);

AO21x2_ASAP7_75t_L g1091 ( 
.A1(n_1017),
.A2(n_118),
.B(n_122),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1023),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1092),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1039),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1054),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_1065),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1041),
.A2(n_1001),
.B(n_1014),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1044),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1052),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_1082),
.Y(n_1100)
);

AOI211xp5_ASAP7_75t_L g1101 ( 
.A1(n_1037),
.A2(n_1011),
.B(n_1007),
.C(n_992),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1058),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1070),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1085),
.B(n_990),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1087),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1070),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_1071),
.B(n_1023),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1088),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1071),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1060),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1090),
.A2(n_998),
.B(n_1015),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1055),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_1049),
.B(n_1015),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1084),
.A2(n_998),
.B(n_1029),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1055),
.Y(n_1115)
);

AO22x1_ASAP7_75t_L g1116 ( 
.A1(n_1080),
.A2(n_990),
.B1(n_126),
.B2(n_127),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1064),
.A2(n_124),
.B(n_131),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1063),
.A2(n_1074),
.B(n_1066),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1067),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1069),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1041),
.A2(n_1059),
.B(n_1062),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1051),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1047),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1067),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1075),
.B(n_1059),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1083),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1047),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1083),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1076),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1068),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1050),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1068),
.B(n_1038),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1040),
.A2(n_132),
.B(n_137),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1045),
.B(n_317),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1089),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_1086),
.B(n_140),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1089),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1091),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1056),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1091),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1078),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_1038),
.Y(n_1142)
);

OAI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1048),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1078),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1078),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1045),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1057),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1053),
.B(n_145),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1079),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_1056),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1036),
.A2(n_1042),
.B1(n_1061),
.B2(n_1037),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1057),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1043),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1104),
.B(n_1110),
.Y(n_1154)
);

XNOR2xp5_ASAP7_75t_L g1155 ( 
.A(n_1139),
.B(n_1073),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_R g1156 ( 
.A(n_1130),
.B(n_1072),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1122),
.B(n_1038),
.Y(n_1157)
);

XNOR2xp5_ASAP7_75t_L g1158 ( 
.A(n_1149),
.B(n_1081),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_R g1159 ( 
.A(n_1130),
.B(n_1135),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1122),
.B(n_1038),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1123),
.B(n_1073),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_R g1162 ( 
.A(n_1130),
.B(n_1077),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1132),
.B(n_1149),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1127),
.B(n_1053),
.Y(n_1164)
);

NAND2xp33_ASAP7_75t_SL g1165 ( 
.A(n_1148),
.B(n_1137),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1104),
.B(n_1081),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_R g1167 ( 
.A(n_1132),
.B(n_1081),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_R g1168 ( 
.A(n_1142),
.B(n_1077),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1103),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1132),
.B(n_1061),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1106),
.B(n_1046),
.Y(n_1171)
);

XOR2x2_ASAP7_75t_SL g1172 ( 
.A(n_1151),
.B(n_1080),
.Y(n_1172)
);

XNOR2xp5_ASAP7_75t_L g1173 ( 
.A(n_1148),
.B(n_1042),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_R g1174 ( 
.A(n_1142),
.B(n_1077),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1098),
.B(n_150),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_R g1176 ( 
.A(n_1131),
.B(n_152),
.Y(n_1176)
);

NAND2xp33_ASAP7_75t_R g1177 ( 
.A(n_1145),
.B(n_1125),
.Y(n_1177)
);

BUFx5_ASAP7_75t_L g1178 ( 
.A(n_1141),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1150),
.B(n_159),
.Y(n_1179)
);

BUFx8_ASAP7_75t_L g1180 ( 
.A(n_1147),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1120),
.B(n_162),
.Y(n_1181)
);

NAND2xp33_ASAP7_75t_R g1182 ( 
.A(n_1145),
.B(n_1125),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_R g1183 ( 
.A(n_1136),
.B(n_1112),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1152),
.B(n_163),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1120),
.B(n_166),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1095),
.B(n_167),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_R g1187 ( 
.A(n_1115),
.B(n_1144),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1095),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_R g1189 ( 
.A(n_1102),
.B(n_168),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_R g1190 ( 
.A(n_1136),
.B(n_1134),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1094),
.B(n_171),
.Y(n_1191)
);

INVxp33_ASAP7_75t_L g1192 ( 
.A(n_1099),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_1136),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1136),
.B(n_173),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1128),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_R g1196 ( 
.A(n_1107),
.B(n_316),
.Y(n_1196)
);

CKINVDCx8_ASAP7_75t_R g1197 ( 
.A(n_1113),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1121),
.B(n_174),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1126),
.B(n_1109),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1105),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1093),
.Y(n_1201)
);

NAND2xp33_ASAP7_75t_R g1202 ( 
.A(n_1134),
.B(n_175),
.Y(n_1202)
);

NAND2xp33_ASAP7_75t_R g1203 ( 
.A(n_1107),
.B(n_176),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1093),
.Y(n_1204)
);

NAND2xp33_ASAP7_75t_R g1205 ( 
.A(n_1129),
.B(n_177),
.Y(n_1205)
);

XNOR2xp5_ASAP7_75t_L g1206 ( 
.A(n_1101),
.B(n_178),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1126),
.B(n_179),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1105),
.B(n_182),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1108),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1116),
.B(n_186),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1194),
.B(n_1138),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1199),
.B(n_1108),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1154),
.B(n_1146),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1201),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1204),
.Y(n_1215)
);

NOR2xp67_ASAP7_75t_L g1216 ( 
.A(n_1195),
.B(n_1138),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1169),
.B(n_1153),
.Y(n_1217)
);

CKINVDCx14_ASAP7_75t_R g1218 ( 
.A(n_1158),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1188),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1166),
.B(n_1153),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1192),
.B(n_1173),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1200),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1209),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1173),
.B(n_1140),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1178),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1165),
.B(n_1146),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1178),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1161),
.B(n_1140),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1178),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1157),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1164),
.B(n_1097),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1178),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1163),
.B(n_1113),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1187),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1155),
.B(n_1116),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1171),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1160),
.B(n_1096),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1170),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1193),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1155),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1197),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1159),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1198),
.B(n_1119),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_1177),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1210),
.B(n_1119),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1183),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1181),
.B(n_1207),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1172),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1206),
.A2(n_1143),
.B1(n_1113),
.B2(n_1096),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1186),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1208),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1196),
.B(n_1124),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1179),
.B(n_1113),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1185),
.B(n_1124),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1214),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1234),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1218),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_R g1258 ( 
.A(n_1230),
.B(n_1205),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1215),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1239),
.B(n_1096),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1224),
.B(n_1100),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1236),
.B(n_1100),
.Y(n_1262)
);

NAND2x1p5_ASAP7_75t_L g1263 ( 
.A(n_1216),
.B(n_1133),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1244),
.B(n_1100),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1219),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1244),
.B(n_1133),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1222),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1227),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1223),
.Y(n_1269)
);

INVx5_ASAP7_75t_SL g1270 ( 
.A(n_1217),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1220),
.B(n_1118),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1217),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1248),
.A2(n_1206),
.B(n_1175),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1219),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1212),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1231),
.B(n_1180),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1221),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1212),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1220),
.B(n_1118),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1228),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1253),
.B(n_1182),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1213),
.B(n_1191),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1245),
.B(n_1189),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1255),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1255),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1259),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1281),
.B(n_1246),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1260),
.B(n_1225),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1275),
.B(n_1229),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1267),
.Y(n_1291)
);

NAND2x1_ASAP7_75t_L g1292 ( 
.A(n_1260),
.B(n_1232),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1267),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1265),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1268),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1284),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1274),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1281),
.B(n_1233),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1269),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1269),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1261),
.B(n_1230),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1278),
.B(n_1226),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_SL g1303 ( 
.A(n_1258),
.B(n_1203),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1296),
.A2(n_1235),
.B1(n_1202),
.B2(n_1190),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1303),
.A2(n_1167),
.B1(n_1235),
.B2(n_1241),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1290),
.Y(n_1306)
);

NAND2xp33_ASAP7_75t_R g1307 ( 
.A(n_1288),
.B(n_1257),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1302),
.B(n_1284),
.Y(n_1308)
);

AND2x4_ASAP7_75t_SL g1309 ( 
.A(n_1298),
.B(n_1242),
.Y(n_1309)
);

AO221x2_ASAP7_75t_L g1310 ( 
.A1(n_1302),
.A2(n_1240),
.B1(n_1276),
.B2(n_1273),
.C(n_1283),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1289),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1287),
.Y(n_1312)
);

CKINVDCx8_ASAP7_75t_R g1313 ( 
.A(n_1289),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_R g1314 ( 
.A(n_1294),
.B(n_1257),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1301),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1296),
.B(n_1280),
.Y(n_1316)
);

CKINVDCx16_ASAP7_75t_R g1317 ( 
.A(n_1307),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1315),
.B(n_1256),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1310),
.A2(n_1176),
.B1(n_1266),
.B2(n_1277),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_L g1320 ( 
.A(n_1305),
.B(n_1266),
.C(n_1297),
.Y(n_1320)
);

AOI22x1_ASAP7_75t_L g1321 ( 
.A1(n_1311),
.A2(n_1306),
.B1(n_1312),
.B2(n_1314),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1309),
.B(n_1256),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1308),
.B(n_1290),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1316),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1313),
.B(n_1292),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1304),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1311),
.B(n_1238),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1316),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1314),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1316),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1318),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1329),
.B(n_1299),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1322),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1317),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1321),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1319),
.A2(n_1260),
.B1(n_1261),
.B2(n_1264),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1319),
.A2(n_1249),
.B1(n_1270),
.B2(n_1211),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1324),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1326),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1338),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1334),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1331),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1339),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1335),
.B(n_1328),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_R g1345 ( 
.A(n_1332),
.B(n_1325),
.Y(n_1345)
);

INVxp33_ASAP7_75t_SL g1346 ( 
.A(n_1343),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1343),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1341),
.Y(n_1348)
);

INVxp33_ASAP7_75t_SL g1349 ( 
.A(n_1345),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1340),
.Y(n_1350)
);

INVx5_ASAP7_75t_SL g1351 ( 
.A(n_1342),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_1347),
.Y(n_1352)
);

NOR3xp33_ASAP7_75t_SL g1353 ( 
.A(n_1350),
.B(n_1344),
.C(n_1337),
.Y(n_1353)
);

OAI221xp5_ASAP7_75t_L g1354 ( 
.A1(n_1348),
.A2(n_1336),
.B1(n_1333),
.B2(n_1320),
.C(n_1325),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1346),
.B(n_1330),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1351),
.B(n_1323),
.Y(n_1356)
);

NOR4xp25_ASAP7_75t_L g1357 ( 
.A(n_1349),
.B(n_1300),
.C(n_1327),
.D(n_1293),
.Y(n_1357)
);

NAND4xp25_ASAP7_75t_L g1358 ( 
.A(n_1351),
.B(n_1252),
.C(n_1264),
.D(n_1247),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1347),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1356),
.Y(n_1360)
);

OAI211xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1353),
.A2(n_1250),
.B(n_1291),
.C(n_1252),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1352),
.A2(n_1184),
.B(n_1286),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1354),
.A2(n_1295),
.B(n_1285),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1357),
.A2(n_1268),
.B1(n_1262),
.B2(n_1174),
.C(n_1168),
.Y(n_1364)
);

OAI22x1_ASAP7_75t_L g1365 ( 
.A1(n_1359),
.A2(n_1211),
.B1(n_1263),
.B2(n_1251),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1355),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1366),
.B(n_1117),
.Y(n_1367)
);

AOI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1360),
.A2(n_1358),
.B1(n_1262),
.B2(n_1237),
.Y(n_1368)
);

NOR2x1_ASAP7_75t_L g1369 ( 
.A(n_1361),
.B(n_1282),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_1363),
.Y(n_1370)
);

NAND2xp33_ASAP7_75t_L g1371 ( 
.A(n_1364),
.B(n_1162),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1362),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1365),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1370),
.B(n_1282),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_R g1375 ( 
.A(n_1371),
.B(n_187),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1373),
.B(n_1272),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1372),
.B(n_1272),
.Y(n_1377)
);

XNOR2xp5_ASAP7_75t_L g1378 ( 
.A(n_1368),
.B(n_1263),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_R g1379 ( 
.A(n_1369),
.B(n_189),
.Y(n_1379)
);

NAND3xp33_ASAP7_75t_L g1380 ( 
.A(n_1367),
.B(n_1279),
.C(n_1271),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1370),
.B(n_1271),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1373),
.B(n_1156),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1373),
.B(n_1263),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1382),
.A2(n_1279),
.B1(n_1270),
.B2(n_1243),
.Y(n_1384)
);

AO22x2_ASAP7_75t_L g1385 ( 
.A1(n_1374),
.A2(n_1254),
.B1(n_1270),
.B2(n_194),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1375),
.Y(n_1386)
);

OA22x2_ASAP7_75t_L g1387 ( 
.A1(n_1383),
.A2(n_1117),
.B1(n_1114),
.B2(n_1270),
.Y(n_1387)
);

AOI221xp5_ASAP7_75t_L g1388 ( 
.A1(n_1379),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.C(n_196),
.Y(n_1388)
);

NAND2xp33_ASAP7_75t_SL g1389 ( 
.A(n_1376),
.B(n_198),
.Y(n_1389)
);

OAI221xp5_ASAP7_75t_L g1390 ( 
.A1(n_1381),
.A2(n_1111),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1377),
.A2(n_1114),
.B1(n_206),
.B2(n_208),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_SL g1392 ( 
.A(n_1380),
.B(n_199),
.C(n_210),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1378),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1393),
.A2(n_1111),
.B1(n_239),
.B2(n_240),
.Y(n_1394)
);

NAND4xp75_ASAP7_75t_L g1395 ( 
.A(n_1388),
.B(n_231),
.C(n_242),
.D(n_243),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1385),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1392),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_1397)
);

NAND4xp25_ASAP7_75t_L g1398 ( 
.A(n_1389),
.B(n_248),
.C(n_249),
.D(n_250),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1386),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_SL g1400 ( 
.A1(n_1384),
.A2(n_251),
.B(n_256),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1390),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1399),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1401),
.A2(n_1391),
.B1(n_1387),
.B2(n_259),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1396),
.A2(n_257),
.B(n_258),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1402),
.A2(n_1400),
.B1(n_1394),
.B2(n_1398),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1403),
.A2(n_1397),
.B1(n_1404),
.B2(n_1395),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1405),
.A2(n_261),
.B1(n_263),
.B2(n_265),
.Y(n_1407)
);

OAI322xp33_ASAP7_75t_L g1408 ( 
.A1(n_1406),
.A2(n_267),
.A3(n_268),
.B1(n_272),
.B2(n_275),
.C1(n_277),
.C2(n_278),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1407),
.A2(n_279),
.B(n_281),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1408),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1407),
.A2(n_285),
.B1(n_288),
.B2(n_290),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1409),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1412),
.A2(n_1410),
.B1(n_1411),
.B2(n_294),
.C(n_295),
.Y(n_1413)
);

AOI211xp5_ASAP7_75t_L g1414 ( 
.A1(n_1413),
.A2(n_292),
.B(n_293),
.C(n_297),
.Y(n_1414)
);


endmodule