module fake_jpeg_15108_n_269 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_38),
.B(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_33),
.B1(n_26),
.B2(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_44),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_22),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_9),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_49),
.B(n_66),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_0),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_56),
.B(n_57),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_43),
.B1(n_36),
.B2(n_19),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_25),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_28),
.B1(n_24),
.B2(n_30),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_58),
.B1(n_62),
.B2(n_24),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_26),
.B1(n_19),
.B2(n_37),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_78),
.B1(n_79),
.B2(n_30),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_52),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_26),
.B1(n_39),
.B2(n_31),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_27),
.B1(n_32),
.B2(n_20),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_22),
.B(n_18),
.C(n_25),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_81),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_20),
.B1(n_22),
.B2(n_18),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_84),
.B1(n_92),
.B2(n_55),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_27),
.B1(n_20),
.B2(n_28),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_22),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_0),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_47),
.B(n_2),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_65),
.B1(n_64),
.B2(n_24),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_47),
.A2(n_24),
.B1(n_28),
.B2(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_96),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_59),
.B1(n_53),
.B2(n_54),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_85),
.B1(n_101),
.B2(n_106),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_52),
.A3(n_69),
.B1(n_51),
.B2(n_60),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_21),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_114),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_81),
.B(n_79),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_62),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_109),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_108),
.B1(n_110),
.B2(n_89),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_58),
.B1(n_63),
.B2(n_61),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_113),
.B1(n_93),
.B2(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_63),
.B1(n_28),
.B2(n_30),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_115),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_72),
.A2(n_63),
.B1(n_21),
.B2(n_30),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_76),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_129),
.B1(n_130),
.B2(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_87),
.C(n_86),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_108),
.C(n_30),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_143),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_87),
.B1(n_85),
.B2(n_81),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_136),
.B(n_23),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_82),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_108),
.B1(n_95),
.B2(n_105),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_93),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_107),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_97),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_146),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_111),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_121),
.B(n_130),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_156),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_108),
.B1(n_112),
.B2(n_99),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_125),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_108),
.B1(n_80),
.B2(n_70),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_126),
.C(n_137),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_160),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_70),
.B1(n_21),
.B2(n_2),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_167),
.B1(n_164),
.B2(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_2),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_70),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_140),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_176),
.B(n_169),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_187),
.C(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_149),
.B(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_146),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_192),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_189),
.B(n_168),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_132),
.B1(n_135),
.B2(n_134),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_185),
.A2(n_190),
.B1(n_153),
.B2(n_156),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_119),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_132),
.C(n_142),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_124),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_145),
.B1(n_157),
.B2(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_173),
.B1(n_7),
.B2(n_8),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_191),
.B(n_179),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_204),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_161),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_173),
.Y(n_223)
);

AOI321xp33_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_160),
.A3(n_159),
.B1(n_162),
.B2(n_139),
.C(n_144),
.Y(n_200)
);

OA21x2_ASAP7_75t_SL g217 ( 
.A1(n_200),
.A2(n_210),
.B(n_175),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_188),
.C(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_207),
.C(n_212),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_180),
.Y(n_218)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_206),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_191),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_148),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_183),
.B(n_179),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_23),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_211),
.Y(n_228)
);

XOR2x2_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_3),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_172),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_6),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_229)
);

OAI322xp33_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_170),
.A3(n_192),
.B1(n_184),
.B2(n_174),
.C1(n_186),
.C2(n_183),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_214),
.A2(n_223),
.B1(n_205),
.B2(n_203),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_180),
.B(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_218),
.B(n_202),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_182),
.B(n_184),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_224),
.B1(n_226),
.B2(n_223),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_6),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_207),
.B(n_194),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_232),
.C(n_235),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_197),
.C(n_212),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_197),
.C(n_200),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_198),
.C(n_7),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_238),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_7),
.C(n_8),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_9),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_240),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_9),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_224),
.B1(n_213),
.B2(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_245),
.C(n_247),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_219),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_11),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_226),
.B1(n_228),
.B2(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_232),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_255),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_254),
.B(n_243),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_11),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_16),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_12),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_259),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_244),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_260),
.B(n_253),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_264),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_13),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_261),
.A2(n_14),
.B(n_15),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_261),
.C(n_263),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_262),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_267),
.Y(n_269)
);


endmodule