module real_jpeg_9378_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_346, n_347, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_346;
input n_347;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_24),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_62),
.B1(n_72),
.B2(n_75),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_62),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_3),
.A2(n_72),
.B1(n_75),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_3),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_163),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_163),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_163),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_4),
.A2(n_36),
.B1(n_72),
.B2(n_75),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_5),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_5),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_5),
.A2(n_135),
.B(n_161),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_10),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_72),
.B1(n_75),
.B2(n_97),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_97),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_97),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_11),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_11),
.A2(n_72),
.B1(n_75),
.B2(n_109),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_109),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_11),
.A2(n_24),
.B1(n_26),
.B2(n_109),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_12),
.A2(n_72),
.B1(n_75),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_12),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_114),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_114),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_114),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_14),
.A2(n_55),
.B(n_67),
.C(n_94),
.D(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_14),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_53),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_14),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_14),
.A2(n_115),
.B(n_117),
.Y(n_137)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_14),
.A2(n_33),
.B(n_49),
.C(n_151),
.D(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_14),
.B(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_14),
.B(n_37),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_14),
.A2(n_30),
.B(n_34),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_14),
.A2(n_24),
.B1(n_26),
.B2(n_132),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_15),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_15),
.A2(n_23),
.B1(n_72),
.B2(n_75),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_15),
.A2(n_23),
.B1(n_54),
.B2(n_55),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_16),
.A2(n_24),
.B1(n_26),
.B2(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_16),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_16),
.A2(n_64),
.B1(n_72),
.B2(n_75),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_16),
.A2(n_54),
.B1(n_55),
.B2(n_64),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_64),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_21),
.B(n_43),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_22),
.A2(n_27),
.B1(n_37),
.B2(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_29),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_24),
.A2(n_29),
.B(n_132),
.C(n_194),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_35),
.B(n_37),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_27),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_27),
.B(n_213),
.Y(n_222)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_28),
.A2(n_32),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_28),
.A2(n_32),
.B1(n_221),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_28),
.A2(n_212),
.B(n_250),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_28),
.A2(n_32),
.B1(n_61),
.B2(n_294),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_32),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_32),
.A2(n_222),
.B(n_294),
.Y(n_293)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_37),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_83),
.B(n_344),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_78),
.C(n_80),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_44),
.A2(n_45),
.B1(n_339),
.B2(n_341),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_59),
.C(n_65),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_46),
.A2(n_47),
.B1(n_65),
.B2(n_319),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_48),
.A2(n_57),
.B1(n_172),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_48),
.A2(n_207),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_48),
.A2(n_56),
.B1(n_57),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_53),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_49),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_49),
.A2(n_53),
.B1(n_247),
.B2(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_49),
.A2(n_53),
.B1(n_266),
.B2(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_51),
.B(n_54),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_52),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_68),
.B(n_70),
.C(n_71),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_68),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_55),
.A2(n_151),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_57),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_57),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_57),
.A2(n_173),
.B(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_59),
.A2(n_60),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_65),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_65),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_76),
.B(n_77),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_66),
.A2(n_76),
.B1(n_108),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_66),
.A2(n_149),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_66),
.A2(n_76),
.B1(n_204),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_66),
.A2(n_76),
.B1(n_232),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_66),
.A2(n_76),
.B1(n_241),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_67),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_67),
.A2(n_71),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_75),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_75),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_72),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_116),
.Y(n_115)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_75),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_108),
.B(n_110),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_76),
.B(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_76),
.A2(n_110),
.B(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_77),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_340),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_78),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_337),
.B(n_343),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_310),
.A3(n_330),
.B1(n_335),
.B2(n_336),
.C(n_346),
.Y(n_84)
);

AOI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_258),
.A3(n_298),
.B1(n_304),
.B2(n_309),
.C(n_347),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_215),
.C(n_254),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_187),
.B(n_214),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_166),
.B(n_186),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_143),
.B(n_165),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_120),
.B(n_142),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_92),
.B(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_93),
.A2(n_98),
.B1(n_99),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_107),
.C(n_112),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_115),
.B(n_117),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_119),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_115),
.A2(n_116),
.B1(n_162),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_115),
.A2(n_116),
.B1(n_177),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_115),
.A2(n_116),
.B1(n_197),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_115),
.A2(n_116),
.B1(n_230),
.B2(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_115),
.A2(n_116),
.B(n_239),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_124),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_132),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_129),
.B(n_141),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_127),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_136),
.B(n_140),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_133),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_145),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_156),
.B2(n_164),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_150),
.B1(n_154),
.B2(n_155),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_155),
.C(n_164),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_156),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_160),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_168),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_182),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_183),
.C(n_184),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_181),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_178),
.C(n_179),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_176),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_178),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_188),
.B(n_189),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_201),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_191),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_191),
.B(n_200),
.C(n_201),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_196),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_203),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_208),
.C(n_209),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_216),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_234),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_217),
.B(n_234),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_228),
.C(n_233),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_227),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_233),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_231),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_252),
.B2(n_253),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_242),
.C(n_253),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_240),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_248),
.C(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_248),
.B1(n_249),
.B2(n_251),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_245),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_256),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_276),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_259),
.B(n_276),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_269),
.C(n_275),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_260),
.A2(n_261),
.B1(n_269),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_265),
.C(n_267),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_269),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_271),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_270),
.A2(n_289),
.B(n_293),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_272),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_272),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_296),
.B2(n_297),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_287),
.B2(n_288),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_288),
.C(n_297),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_284),
.B(n_286),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_284),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_285),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_286),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_286),
.A2(n_312),
.B1(n_321),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_295),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_291),
.Y(n_295)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_296),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_305),
.B(n_308),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_301),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_323),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_323),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_321),
.C(n_322),
.Y(n_311)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_313),
.A2(n_314),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_319),
.C(n_320),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_325),
.C(n_329),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_317),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_333),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_331),
.B(n_332),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_342),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_339),
.Y(n_341)
);


endmodule