module fake_jpeg_7322_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_20),
.B1(n_18),
.B2(n_35),
.Y(n_58)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx2_ASAP7_75t_SL g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_45),
.B1(n_29),
.B2(n_31),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_17),
.C(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_18),
.B1(n_35),
.B2(n_24),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_32),
.B1(n_29),
.B2(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_87),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_57),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_74),
.A2(n_29),
.B1(n_19),
.B2(n_22),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_42),
.B1(n_18),
.B2(n_31),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_42),
.B1(n_46),
.B2(n_38),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_92),
.Y(n_108)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_44),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_62),
.Y(n_100)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_94),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_64),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_28),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_22),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_76),
.Y(n_117)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_61),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_125),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_110),
.B1(n_28),
.B2(n_33),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_40),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

AO21x2_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_70),
.B(n_97),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_127),
.A2(n_21),
.B1(n_118),
.B2(n_82),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_80),
.B(n_77),
.C(n_71),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_129),
.A2(n_133),
.B(n_141),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_104),
.B(n_98),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_32),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_150),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_40),
.C(n_44),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_148),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_46),
.B1(n_59),
.B2(n_77),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_151),
.B1(n_103),
.B2(n_126),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_32),
.B(n_25),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_33),
.B1(n_21),
.B2(n_38),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_146),
.B(n_149),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_59),
.B1(n_95),
.B2(n_79),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_145),
.A2(n_153),
.B1(n_56),
.B2(n_82),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_105),
.B(n_101),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_41),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_56),
.B1(n_79),
.B2(n_49),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_93),
.B1(n_89),
.B2(n_49),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_112),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_162),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_99),
.B1(n_107),
.B2(n_116),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_165),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_157),
.B(n_164),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_146),
.B1(n_135),
.B2(n_144),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_44),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_163),
.B(n_182),
.Y(n_193)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_120),
.B1(n_114),
.B2(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_104),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_167),
.A2(n_170),
.B1(n_172),
.B2(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_168),
.B(n_173),
.Y(n_204)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_169),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_178),
.B1(n_180),
.B2(n_154),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_27),
.B1(n_24),
.B2(n_23),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_98),
.B1(n_41),
.B2(n_30),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_174),
.A2(n_170),
.B1(n_173),
.B2(n_169),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_131),
.A2(n_98),
.B1(n_14),
.B2(n_15),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_24),
.A3(n_27),
.B1(n_23),
.B2(n_30),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_41),
.B1(n_30),
.B2(n_23),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_132),
.B1(n_138),
.B2(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_26),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_183),
.A2(n_141),
.B(n_151),
.Y(n_187)
);

BUFx24_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_181),
.B1(n_180),
.B2(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_195),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_194),
.B(n_207),
.Y(n_227)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_197),
.A2(n_199),
.B(n_200),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_171),
.B1(n_164),
.B2(n_168),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_210),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_184),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_148),
.B(n_149),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_213),
.B(n_211),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_149),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_208),
.C(n_213),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_211),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_154),
.B(n_147),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_155),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_218),
.B(n_221),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_226),
.B1(n_237),
.B2(n_190),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_174),
.B1(n_179),
.B2(n_183),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_230),
.B1(n_232),
.B2(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_223),
.B(n_235),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_162),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_225),
.C(n_231),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_159),
.C(n_136),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_130),
.B1(n_30),
.B2(n_27),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_228),
.B(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_200),
.A2(n_26),
.B1(n_40),
.B2(n_44),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_26),
.C(n_34),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_188),
.A2(n_26),
.B1(n_34),
.B2(n_2),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_34),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_190),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_186),
.A2(n_0),
.B(n_1),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_191),
.B(n_186),
.C(n_192),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_34),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_191),
.C(n_188),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_236),
.B(n_216),
.Y(n_268)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_196),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_233),
.C(n_222),
.Y(n_267)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_225),
.B(n_197),
.CI(n_206),
.CON(n_248),
.SN(n_248)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_256),
.Y(n_264)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_202),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_253),
.Y(n_277)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_210),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_212),
.B1(n_9),
.B2(n_10),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_259),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_263),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_260),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_7),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_270),
.C(n_275),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_239),
.C(n_231),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_230),
.B1(n_236),
.B2(n_219),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_240),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_247),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_238),
.C(n_232),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_237),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_243),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_7),
.B(n_14),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_254),
.C(n_245),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_267),
.C(n_266),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_285),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_269),
.Y(n_299)
);

OAI21x1_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_263),
.B(n_241),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_271),
.B(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_289),
.C(n_11),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_241),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_260),
.B1(n_246),
.B2(n_241),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_262),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_292),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_16),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_295),
.B(n_265),
.Y(n_297)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_11),
.B(n_12),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_301),
.Y(n_313)
);

NOR4xp25_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_269),
.C(n_275),
.D(n_277),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_300),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_306),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_282),
.C(n_288),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_293),
.A2(n_277),
.B1(n_272),
.B2(n_10),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_305),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_304),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_11),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_308),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_282),
.B(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_4),
.B(n_5),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_6),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_289),
.C(n_13),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_13),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_4),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_303),
.B(n_304),
.Y(n_320)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_325),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_327),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

AOI211xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_313),
.B(n_310),
.C(n_6),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_318),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_324),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_326),
.B(n_328),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_323),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_331),
.B(n_332),
.Y(n_338)
);


endmodule