module fake_netlist_6_2462_n_692 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_692);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_692;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_647;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_594;
wire n_565;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_655;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_688;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_15),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_85),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_93),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_L g141 ( 
.A(n_42),
.B(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_39),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_14),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_63),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_12),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_46),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g151 ( 
.A(n_60),
.B(n_29),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_68),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_58),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_83),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_48),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_43),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_92),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_32),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_16),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_53),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_25),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_41),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_14),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_28),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_2),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_15),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_64),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_102),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_101),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_132),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_27),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_76),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_70),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_100),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_22),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_0),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_145),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_21),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_146),
.B(n_3),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_23),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_6),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_6),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_170),
.Y(n_209)
);

OAI22x1_ASAP7_75t_SL g210 ( 
.A1(n_167),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_161),
.A2(n_170),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_135),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_144),
.A2(n_10),
.B(n_11),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_147),
.B(n_10),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_163),
.B(n_11),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_135),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

BUFx8_ASAP7_75t_SL g221 ( 
.A(n_140),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_165),
.A2(n_13),
.B(n_18),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_172),
.A2(n_18),
.B(n_19),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_156),
.B(n_19),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_195),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_211),
.B(n_140),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_195),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_192),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_134),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_166),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_216),
.B(n_166),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_168),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_225),
.B(n_168),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_190),
.B(n_137),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_225),
.B(n_141),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_202),
.A2(n_151),
.B(n_183),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_198),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_202),
.B(n_151),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_198),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_221),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_212),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_184),
.C(n_182),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_202),
.B(n_208),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_190),
.B(n_180),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_143),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_192),
.B(n_179),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_152),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_178),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_214),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_188),
.B(n_175),
.C(n_173),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_200),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_253),
.B(n_201),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_219),
.B1(n_189),
.B2(n_187),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_259),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_223),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_224),
.B(n_203),
.C(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_228),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_233),
.B(n_252),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_238),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_229),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_193),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_204),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_204),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_194),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_194),
.B1(n_199),
.B2(n_206),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_204),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_231),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_251),
.B(n_153),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_217),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_247),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_248),
.A2(n_244),
.B1(n_264),
.B2(n_274),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_217),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_199),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_231),
.B(n_196),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_197),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_217),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_249),
.Y(n_315)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_240),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_249),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_232),
.B(n_220),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_232),
.Y(n_320)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_236),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_154),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_254),
.B(n_155),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_230),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_273),
.B(n_159),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_235),
.A2(n_222),
.B1(n_215),
.B2(n_224),
.Y(n_327)
);

NAND2xp33_ASAP7_75t_L g328 ( 
.A(n_258),
.B(n_197),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_236),
.A2(n_197),
.B1(n_210),
.B2(n_215),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_258),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_254),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_301),
.A2(n_314),
.B(n_308),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_215),
.B(n_222),
.C(n_263),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_260),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_255),
.B(n_275),
.Y(n_335)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_255),
.B(n_271),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_260),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_271),
.B(n_256),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

NAND2xp33_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_197),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_256),
.B(n_246),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_289),
.A2(n_256),
.B(n_246),
.C(n_245),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_236),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_282),
.B(n_236),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_289),
.B(n_245),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_321),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_221),
.Y(n_349)
);

O2A1O1Ixp5_ASAP7_75t_L g350 ( 
.A1(n_277),
.A2(n_245),
.B(n_24),
.C(n_26),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_277),
.A2(n_245),
.B1(n_30),
.B2(n_33),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_288),
.B(n_297),
.Y(n_352)
);

A2O1A1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_323),
.A2(n_20),
.B(n_34),
.C(n_35),
.Y(n_353)
);

AOI21x1_ASAP7_75t_L g354 ( 
.A1(n_290),
.A2(n_88),
.B(n_36),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_280),
.A2(n_327),
.B1(n_323),
.B2(n_325),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_280),
.A2(n_89),
.B(n_37),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_293),
.B(n_20),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_38),
.Y(n_358)
);

NOR2x1_ASAP7_75t_L g359 ( 
.A(n_293),
.B(n_40),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_287),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_44),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g364 ( 
.A1(n_279),
.A2(n_45),
.B(n_47),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_278),
.B(n_52),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_284),
.B(n_55),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_56),
.B(n_57),
.Y(n_368)
);

A2O1A1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_283),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_310),
.B(n_320),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_287),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_309),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_69),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_296),
.B(n_71),
.Y(n_374)
);

AND2x6_ASAP7_75t_SL g375 ( 
.A(n_281),
.B(n_73),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_329),
.A2(n_74),
.B1(n_77),
.B2(n_79),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_316),
.B(n_80),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_316),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_81),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_316),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_294),
.B(n_87),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_300),
.A2(n_90),
.B1(n_91),
.B2(n_94),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_305),
.B(n_95),
.Y(n_383)
);

NOR3xp33_ASAP7_75t_L g384 ( 
.A(n_315),
.B(n_317),
.C(n_298),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_292),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_292),
.B(n_97),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_298),
.B(n_98),
.Y(n_387)
);

O2A1O1Ixp33_ASAP7_75t_L g388 ( 
.A1(n_302),
.A2(n_106),
.B(n_107),
.C(n_109),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_332),
.A2(n_342),
.B(n_339),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_341),
.A2(n_303),
.B(n_318),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_303),
.Y(n_391)
);

OAI21x1_ASAP7_75t_L g392 ( 
.A1(n_335),
.A2(n_322),
.B(n_318),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_371),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_355),
.A2(n_345),
.B(n_360),
.Y(n_394)
);

AO21x1_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_322),
.B(n_312),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_331),
.A2(n_312),
.B1(n_311),
.B2(n_306),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_311),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_344),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_306),
.B(n_304),
.C(n_110),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_304),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g401 ( 
.A1(n_337),
.A2(n_111),
.B(n_112),
.Y(n_401)
);

AO31x2_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_116),
.A3(n_117),
.B(n_118),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_336),
.A2(n_119),
.B(n_121),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_336),
.A2(n_360),
.B(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_361),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_362),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_340),
.B(n_128),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g409 ( 
.A(n_359),
.B(n_129),
.Y(n_409)
);

NAND2x1_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_130),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_349),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

AO32x2_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_131),
.A3(n_351),
.B1(n_380),
.B2(n_382),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_352),
.Y(n_414)
);

BUFx4f_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_346),
.B(n_384),
.Y(n_416)
);

NOR4xp25_ASAP7_75t_L g417 ( 
.A(n_357),
.B(n_353),
.C(n_372),
.D(n_388),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_333),
.A2(n_343),
.B(n_350),
.Y(n_418)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_366),
.A2(n_383),
.B(n_374),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_346),
.B(n_378),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_385),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_348),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_348),
.B(n_379),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_381),
.B(n_358),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g425 ( 
.A1(n_367),
.A2(n_387),
.B(n_386),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_368),
.A2(n_363),
.B(n_356),
.Y(n_426)
);

NAND2x1p5_ASAP7_75t_L g427 ( 
.A(n_354),
.B(n_375),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_332),
.A2(n_342),
.B(n_339),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_331),
.B(n_230),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g430 ( 
.A1(n_332),
.A2(n_342),
.B(n_339),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_334),
.B(n_286),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_334),
.B(n_286),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_355),
.A2(n_331),
.B1(n_248),
.B2(n_257),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_431),
.B(n_432),
.Y(n_435)
);

INVx3_ASAP7_75t_SL g436 ( 
.A(n_414),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_408),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_433),
.A2(n_424),
.B1(n_429),
.B2(n_398),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_412),
.Y(n_439)
);

OAI21x1_ASAP7_75t_SL g440 ( 
.A1(n_395),
.A2(n_394),
.B(n_418),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_411),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_393),
.B(n_420),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_389),
.A2(n_430),
.B(n_428),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_405),
.A2(n_427),
.B1(n_407),
.B2(n_409),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_391),
.B(n_423),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_397),
.B(n_434),
.Y(n_446)
);

BUFx4f_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_434),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_415),
.A2(n_434),
.B1(n_399),
.B2(n_422),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_415),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_426),
.A2(n_390),
.B(n_401),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_400),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_404),
.A2(n_396),
.B(n_409),
.Y(n_455)
);

AO21x2_ASAP7_75t_L g456 ( 
.A1(n_417),
.A2(n_403),
.B(n_406),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_417),
.A2(n_402),
.B(n_413),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_402),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_419),
.A2(n_433),
.B1(n_429),
.B2(n_253),
.Y(n_459)
);

AOI221xp5_ASAP7_75t_L g460 ( 
.A1(n_402),
.A2(n_279),
.B1(n_257),
.B2(n_273),
.C(n_433),
.Y(n_460)
);

NAND2x1p5_ASAP7_75t_L g461 ( 
.A(n_419),
.B(n_425),
.Y(n_461)
);

OAI221xp5_ASAP7_75t_L g462 ( 
.A1(n_429),
.A2(n_257),
.B1(n_248),
.B2(n_253),
.C(n_244),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_393),
.Y(n_464)
);

O2A1O1Ixp33_ASAP7_75t_SL g465 ( 
.A1(n_424),
.A2(n_364),
.B(n_369),
.C(n_398),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_432),
.Y(n_466)
);

AOI21xp33_ASAP7_75t_SL g467 ( 
.A1(n_429),
.A2(n_257),
.B(n_273),
.Y(n_467)
);

AO31x2_ASAP7_75t_L g468 ( 
.A1(n_395),
.A2(n_433),
.A3(n_283),
.B(n_355),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_326),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_408),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_471),
.A2(n_466),
.B1(n_459),
.B2(n_438),
.Y(n_475)
);

NAND2x1_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_449),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_474),
.Y(n_477)
);

AO21x2_ASAP7_75t_L g478 ( 
.A1(n_440),
.A2(n_452),
.B(n_443),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_474),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_438),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_473),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_469),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_470),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_472),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_437),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

BUFx5_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_442),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_435),
.B(n_445),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_454),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_439),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_437),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_454),
.Y(n_498)
);

AND4x1_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_444),
.C(n_462),
.D(n_441),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_463),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_446),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_468),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_446),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_448),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_468),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_468),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_483),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_458),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_496),
.B(n_467),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_457),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_491),
.Y(n_514)
);

NAND2x1_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_450),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_458),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_441),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_457),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_502),
.B(n_457),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_436),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_504),
.B(n_436),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_479),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_492),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_476),
.Y(n_524)
);

AND2x4_ASAP7_75t_SL g525 ( 
.A(n_501),
.B(n_437),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_479),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_475),
.A2(n_456),
.B1(n_436),
.B2(n_453),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_491),
.B(n_457),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_482),
.B(n_456),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_491),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_463),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_483),
.A2(n_456),
.B1(n_500),
.B2(n_501),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_506),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_500),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_480),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_491),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_484),
.B(n_450),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_478),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_484),
.B(n_455),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_499),
.B(n_451),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_485),
.B(n_461),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_491),
.B(n_461),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_480),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_485),
.B(n_461),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_489),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_486),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_522),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_522),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_528),
.B(n_506),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_526),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_526),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_535),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_513),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_514),
.B(n_486),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_510),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_513),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_518),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_511),
.B(n_516),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_512),
.B(n_495),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_SL g560 ( 
.A1(n_517),
.A2(n_491),
.B1(n_501),
.B2(n_477),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_511),
.B(n_491),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_520),
.B(n_495),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_516),
.B(n_509),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_519),
.B(n_508),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_518),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_533),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_533),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_540),
.A2(n_490),
.B1(n_488),
.B2(n_487),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_521),
.A2(n_451),
.B1(n_455),
.B2(n_490),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_519),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_529),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_529),
.B(n_508),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_514),
.B(n_497),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_542),
.B(n_507),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_542),
.B(n_503),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_535),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_523),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_561),
.B(n_536),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_562),
.B(n_534),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_561),
.B(n_539),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_571),
.B(n_539),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_547),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_571),
.B(n_539),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_576),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_527),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_578),
.B(n_515),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_566),
.B(n_524),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_555),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_547),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_548),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_566),
.B(n_539),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_576),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_578),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_558),
.B(n_515),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_538),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_558),
.B(n_541),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_548),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_567),
.B(n_570),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_570),
.B(n_538),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_563),
.B(n_541),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_572),
.B(n_564),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_553),
.B(n_538),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_563),
.B(n_544),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_577),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_550),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_551),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_580),
.B(n_554),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_585),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_585),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_593),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_588),
.B(n_577),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_581),
.B(n_557),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_594),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_605),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_583),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_593),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_607),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_581),
.B(n_602),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_586),
.A2(n_560),
.B1(n_568),
.B2(n_532),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_597),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_607),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_SL g623 ( 
.A(n_587),
.B(n_537),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_606),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_599),
.B(n_557),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_606),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_579),
.B(n_595),
.Y(n_628)
);

OAI32xp33_ASAP7_75t_L g629 ( 
.A1(n_623),
.A2(n_589),
.A3(n_596),
.B1(n_604),
.B2(n_601),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_620),
.A2(n_569),
.B1(n_555),
.B2(n_579),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_621),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_608),
.A2(n_592),
.B(n_582),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_615),
.B(n_619),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_628),
.A2(n_575),
.B1(n_574),
.B2(n_549),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_618),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_622),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_609),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_531),
.C(n_537),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_616),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_609),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_619),
.B(n_602),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_610),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_642),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_635),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_636),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_630),
.A2(n_614),
.B1(n_592),
.B2(n_627),
.Y(n_646)
);

AOI322xp5_ASAP7_75t_L g647 ( 
.A1(n_638),
.A2(n_613),
.A3(n_611),
.B1(n_617),
.B2(n_626),
.C1(n_624),
.C2(n_584),
.Y(n_647)
);

AOI221xp5_ASAP7_75t_L g648 ( 
.A1(n_629),
.A2(n_614),
.B1(n_613),
.B2(n_616),
.C(n_588),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_646),
.B(n_631),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g650 ( 
.A1(n_648),
.A2(n_632),
.B(n_633),
.Y(n_650)
);

AOI222xp33_ASAP7_75t_L g651 ( 
.A1(n_643),
.A2(n_634),
.B1(n_639),
.B2(n_641),
.C1(n_637),
.C2(n_640),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_647),
.B(n_612),
.Y(n_652)
);

OAI222xp33_ASAP7_75t_L g653 ( 
.A1(n_644),
.A2(n_612),
.B1(n_639),
.B2(n_625),
.C1(n_582),
.C2(n_584),
.Y(n_653)
);

AOI221x1_ASAP7_75t_L g654 ( 
.A1(n_645),
.A2(n_598),
.B1(n_588),
.B2(n_591),
.C(n_590),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_651),
.B(n_591),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_650),
.B(n_590),
.Y(n_656)
);

NAND4xp25_ASAP7_75t_L g657 ( 
.A(n_652),
.B(n_552),
.C(n_596),
.D(n_573),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_649),
.B(n_583),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_SL g659 ( 
.A(n_657),
.B(n_653),
.C(n_543),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_SL g660 ( 
.A(n_656),
.B(n_654),
.C(n_543),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_L g661 ( 
.A(n_658),
.B(n_545),
.C(n_465),
.Y(n_661)
);

NOR2x1_ASAP7_75t_SL g662 ( 
.A(n_660),
.B(n_655),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_659),
.B(n_573),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_661),
.B(n_600),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_R g665 ( 
.A(n_659),
.B(n_497),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_662),
.B(n_600),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_665),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_663),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_664),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_662),
.B(n_525),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_662),
.B(n_525),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_664),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_667),
.B(n_525),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_669),
.B(n_603),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_670),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_668),
.B(n_554),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_672),
.B(n_556),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_675),
.A2(n_666),
.B1(n_671),
.B2(n_603),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_677),
.Y(n_679)
);

AOI221xp5_ASAP7_75t_SL g680 ( 
.A1(n_674),
.A2(n_666),
.B1(n_546),
.B2(n_556),
.C(n_553),
.Y(n_680)
);

OA22x2_ASAP7_75t_L g681 ( 
.A1(n_676),
.A2(n_545),
.B1(n_546),
.B2(n_573),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_679),
.Y(n_682)
);

AOI22x1_ASAP7_75t_L g683 ( 
.A1(n_678),
.A2(n_673),
.B1(n_489),
.B2(n_497),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_681),
.A2(n_680),
.B1(n_447),
.B2(n_565),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_682),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_683),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_684),
.A2(n_447),
.B1(n_565),
.B2(n_549),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_685),
.B(n_554),
.Y(n_688)
);

OA21x2_ASAP7_75t_L g689 ( 
.A1(n_686),
.A2(n_447),
.B(n_498),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_688),
.B(n_687),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_690),
.B(n_689),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_691),
.A2(n_689),
.B1(n_489),
.B2(n_545),
.Y(n_692)
);


endmodule