module fake_jpeg_15949_n_291 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_291);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_291;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_20;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_44),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_49),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_39),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_47),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_28),
.Y(n_49)
);

BUFx2_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_51),
.B(n_52),
.Y(n_92)
);

NOR2xp67_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_65),
.Y(n_78)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_33),
.B1(n_26),
.B2(n_42),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_61),
.B1(n_39),
.B2(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_33),
.B1(n_29),
.B2(n_23),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_35),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_22),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_75),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_80),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_44),
.C(n_27),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_74),
.C(n_64),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_43),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_60),
.Y(n_110)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_29),
.B1(n_23),
.B2(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_23),
.B1(n_34),
.B2(n_25),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_34),
.B1(n_25),
.B2(n_17),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_55),
.B1(n_39),
.B2(n_57),
.Y(n_104)
);

NAND2x1_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_47),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_99),
.B(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_48),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_57),
.B1(n_60),
.B2(n_19),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_110),
.B1(n_111),
.B2(n_74),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_91),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_64),
.B(n_25),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_115),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_92),
.B1(n_84),
.B2(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_72),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_60),
.B1(n_42),
.B2(n_55),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_78),
.B1(n_71),
.B2(n_42),
.Y(n_128)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_122),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_98),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_74),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_24),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_94),
.B1(n_110),
.B2(n_116),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_131),
.C(n_137),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_69),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_132),
.A2(n_135),
.B(n_102),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_95),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_141),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_17),
.B(n_31),
.C(n_30),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_24),
.B(n_30),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_72),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_168),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_146),
.A2(n_169),
.B1(n_31),
.B2(n_21),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_138),
.C(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_101),
.Y(n_157)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_105),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_160),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_163),
.B(n_17),
.Y(n_179)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_162),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_113),
.B(n_112),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_32),
.B(n_20),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_97),
.B1(n_114),
.B2(n_118),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_123),
.B1(n_135),
.B2(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_58),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_117),
.B1(n_80),
.B2(n_31),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_183),
.C(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_171),
.B(n_153),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_134),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_178),
.B1(n_180),
.B2(n_193),
.Y(n_203)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_140),
.B1(n_139),
.B2(n_58),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_188),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_130),
.B1(n_80),
.B2(n_139),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_149),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_139),
.B1(n_124),
.B2(n_125),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_125),
.B1(n_124),
.B2(n_32),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_169),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_27),
.C(n_72),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_160),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_157),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_196),
.C(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_168),
.C(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_147),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_202),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_147),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_144),
.C(n_150),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_175),
.C(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_155),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_179),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_212),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_149),
.B1(n_167),
.B2(n_151),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_181),
.B1(n_189),
.B2(n_156),
.Y(n_232)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_190),
.B1(n_177),
.B2(n_186),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_225),
.B1(n_229),
.B2(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_194),
.C(n_18),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_203),
.B1(n_206),
.B2(n_201),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_204),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_192),
.B1(n_176),
.B2(n_145),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_176),
.B1(n_162),
.B2(n_154),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_178),
.B1(n_181),
.B2(n_166),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_224),
.A2(n_208),
.B(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_195),
.C(n_202),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_241),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_242),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_240),
.C(n_247),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_22),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_18),
.C(n_20),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_18),
.C(n_16),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_15),
.C(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_246),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_0),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_226),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_216),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_233),
.B(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_227),
.C(n_1),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_223),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_222),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_268),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_245),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_264),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_237),
.B1(n_236),
.B2(n_240),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_256),
.C(n_253),
.Y(n_269)
);

XNOR2x2_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_2),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_257),
.B(n_253),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_3),
.B(n_4),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_11),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_270),
.C(n_8),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_256),
.C(n_1),
.Y(n_270)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_276),
.B(n_6),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_259),
.B(n_264),
.Y(n_277)
);

AOI221xp5_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_278),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_271),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_282),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_7),
.B(n_8),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_8),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_284),
.B(n_9),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_9),
.B(n_10),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_286),
.B(n_10),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_10),
.Y(n_291)
);


endmodule