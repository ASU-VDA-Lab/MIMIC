module fake_jpeg_14598_n_25 (n_3, n_2, n_1, n_0, n_4, n_25);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_25;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g5 ( 
.A(n_0),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_0),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_6),
.B(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_6),
.B(n_3),
.Y(n_10)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_10),
.A2(n_11),
.B(n_12),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_12),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_8),
.Y(n_17)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_18),
.B(n_15),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_13),
.A2(n_8),
.B1(n_1),
.B2(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_1),
.B1(n_18),
.B2(n_20),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_23),
.A2(n_22),
.B(n_1),
.Y(n_24)
);

BUFx24_ASAP7_75t_SL g25 ( 
.A(n_24),
.Y(n_25)
);


endmodule