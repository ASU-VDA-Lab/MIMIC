module fake_netlist_6_887_n_2061 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2061);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2061;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_93),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_75),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_127),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_106),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_69),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_86),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_123),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_101),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_49),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_35),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_163),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_87),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_11),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_82),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_74),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_114),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_80),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_107),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_25),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_56),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_14),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_6),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_95),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_2),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_71),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_138),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_63),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_188),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_206),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_119),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_115),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_24),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_158),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_112),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_108),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_10),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_110),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_176),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_161),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_116),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_98),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_85),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_96),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_118),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_32),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_57),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_49),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_23),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_11),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_92),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_105),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_21),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_121),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_168),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_194),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_20),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_26),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_26),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_0),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_31),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_73),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_130),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_160),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_42),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_62),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_144),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_13),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_88),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_113),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_16),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_37),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_69),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_9),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_3),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_68),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_66),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_181),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_157),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_14),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_23),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_124),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_36),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_68),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_43),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_182),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_136),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_149),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_191),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_141),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_198),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_117),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_137),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_21),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_97),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_1),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_24),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_43),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_64),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_142),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_145),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_60),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_156),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_18),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_7),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_53),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_111),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_162),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_27),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_36),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_104),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_79),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_125),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_193),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_170),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_37),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_2),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_56),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_100),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_166),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_169),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_8),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_19),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_65),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_102),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_71),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_73),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_53),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_143),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_6),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_60),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_18),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_131),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_77),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_50),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_186),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_29),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_147),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_1),
.Y(n_357)
);

CKINVDCx11_ASAP7_75t_R g358 ( 
.A(n_184),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_195),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_173),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_9),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_29),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_154),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_75),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_61),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_128),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_27),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_201),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_72),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_13),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_54),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_19),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_81),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_135),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_164),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_89),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_84),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_171),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_196),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_40),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_208),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_55),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_77),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_65),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_129),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_205),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_210),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_51),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_148),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_59),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_34),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_15),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_16),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_46),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_197),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_146),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_99),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_177),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_20),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_0),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_58),
.Y(n_401)
);

BUFx2_ASAP7_75t_SL g402 ( 
.A(n_32),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_48),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_79),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_103),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_66),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_4),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_57),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_47),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_183),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_109),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_134),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_4),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_58),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_3),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_64),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_31),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_45),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_277),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_358),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_277),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_213),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_277),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_214),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_233),
.B(n_5),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_277),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_211),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_277),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_245),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_300),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_217),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_387),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_218),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_396),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_277),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_R g436 ( 
.A(n_274),
.B(n_83),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_398),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_277),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_277),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_231),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_220),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_224),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_386),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_277),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_342),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_342),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_342),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_225),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_248),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_342),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_342),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_230),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_405),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_248),
.B(n_7),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_219),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_230),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_275),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_233),
.B(n_8),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_333),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_275),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_300),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_292),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_292),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_280),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_300),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_333),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_395),
.B(n_412),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_293),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_280),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_395),
.B(n_10),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_412),
.B(n_12),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_293),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_226),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_238),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_219),
.B(n_12),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_413),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_243),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_246),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_247),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_249),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_400),
.Y(n_482)
);

BUFx2_ASAP7_75t_SL g483 ( 
.A(n_341),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_413),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_250),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_400),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_417),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_263),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_417),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_253),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_216),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_286),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_240),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_240),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_240),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_244),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_254),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_222),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_244),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_244),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_323),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_255),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_323),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_258),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_323),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_350),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_259),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_261),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_281),
.B(n_15),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_286),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_350),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_269),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_272),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_223),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_212),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_227),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_R g519 ( 
.A(n_273),
.B(n_209),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_350),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_287),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_296),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_391),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_391),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_391),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_445),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_445),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_495),
.B(n_215),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_460),
.A2(n_315),
.B1(n_344),
.B2(n_278),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_456),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_446),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_430),
.B(n_304),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_447),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_425),
.A2(n_355),
.B1(n_382),
.B2(n_367),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_447),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_428),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_430),
.B(n_306),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_215),
.Y(n_540)
);

OA21x2_ASAP7_75t_L g541 ( 
.A1(n_448),
.A2(n_232),
.B(n_212),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_221),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_448),
.B(n_281),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_486),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_491),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_421),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_474),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_451),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_430),
.B(n_308),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_451),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_456),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_421),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_456),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_452),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_478),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_423),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_452),
.Y(n_560)
);

AND3x2_ASAP7_75t_L g561 ( 
.A(n_455),
.B(n_471),
.C(n_472),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_456),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_512),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_426),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_435),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_435),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_489),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_438),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_499),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_439),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_439),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_516),
.Y(n_577)
);

AND2x6_ASAP7_75t_L g578 ( 
.A(n_444),
.B(n_297),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_444),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_453),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_457),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_457),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_518),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_458),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_R g586 ( 
.A(n_482),
.B(n_234),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_458),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_461),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_462),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_461),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_463),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_468),
.B(n_326),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_459),
.B(n_368),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_463),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_464),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_464),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_469),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_469),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_473),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_473),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_477),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_477),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_467),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_494),
.B(n_221),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_484),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_484),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_487),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_487),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_494),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_610),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_589),
.B(n_422),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_593),
.B(n_564),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_531),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_593),
.B(n_424),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_594),
.B(n_431),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_594),
.B(n_433),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_528),
.B(n_455),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_531),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_528),
.A2(n_482),
.B1(n_443),
.B2(n_440),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_578),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_533),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_610),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_576),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_546),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_528),
.B(n_297),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_546),
.Y(n_627)
);

BUFx4f_ASAP7_75t_L g628 ( 
.A(n_541),
.Y(n_628)
);

INVx6_ASAP7_75t_L g629 ( 
.A(n_589),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_531),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_576),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_534),
.B(n_493),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_576),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_564),
.B(n_441),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_575),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_575),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_540),
.A2(n_511),
.B1(n_476),
.B2(n_488),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_536),
.A2(n_481),
.B1(n_485),
.B2(n_479),
.Y(n_638)
);

AO21x2_ASAP7_75t_L g639 ( 
.A1(n_534),
.A2(n_436),
.B(n_229),
.Y(n_639)
);

INVxp33_ASAP7_75t_L g640 ( 
.A(n_547),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_533),
.Y(n_641)
);

AND3x2_ASAP7_75t_L g642 ( 
.A(n_547),
.B(n_312),
.C(n_360),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_533),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_578),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_540),
.A2(n_465),
.B1(n_470),
.B2(n_450),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_531),
.Y(n_646)
);

OAI21xp33_ASAP7_75t_SL g647 ( 
.A1(n_540),
.A2(n_237),
.B(n_232),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g648 ( 
.A1(n_566),
.A2(n_229),
.B(n_228),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_531),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_579),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_538),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_589),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_531),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_579),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_589),
.B(n_442),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_530),
.A2(n_493),
.B1(n_429),
.B2(n_432),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_590),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_L g658 ( 
.A1(n_536),
.A2(n_393),
.B1(n_365),
.B2(n_235),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_586),
.A2(n_505),
.B1(n_492),
.B2(n_236),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_590),
.B(n_449),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_590),
.B(n_475),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_566),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_538),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_586),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_590),
.B(n_480),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_538),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_566),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_SL g668 ( 
.A(n_574),
.B(n_490),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_576),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_538),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_577),
.B(n_498),
.Y(n_671)
);

BUFx8_ASAP7_75t_SL g672 ( 
.A(n_604),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_577),
.B(n_503),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_584),
.B(n_506),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_542),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_568),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_544),
.A2(n_414),
.B1(n_341),
.B2(n_462),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_584),
.B(n_509),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_539),
.B(n_510),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_531),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_542),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_549),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_568),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_539),
.B(n_515),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_542),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_576),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_551),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_542),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_544),
.B(n_360),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_549),
.B(n_420),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_558),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_551),
.B(n_521),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_578),
.B(n_389),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_543),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_568),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_543),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_569),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_569),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_531),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_574),
.B(n_522),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_569),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_605),
.B(n_466),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_541),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_544),
.A2(n_252),
.B1(n_260),
.B2(n_239),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_543),
.Y(n_705)
);

AND2x2_ASAP7_75t_SL g706 ( 
.A(n_541),
.B(n_389),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_570),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_543),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_605),
.B(n_545),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_553),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_548),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_570),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_553),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_548),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_561),
.A2(n_266),
.B1(n_267),
.B2(n_265),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_561),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_570),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_548),
.Y(n_718)
);

INVx6_ASAP7_75t_L g719 ( 
.A(n_576),
.Y(n_719)
);

INVx6_ASAP7_75t_L g720 ( 
.A(n_576),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_558),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_567),
.B(n_466),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_548),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_605),
.B(n_514),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_567),
.B(n_483),
.Y(n_725)
);

BUFx8_ASAP7_75t_SL g726 ( 
.A(n_604),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_553),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_567),
.B(n_466),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_604),
.B(n_483),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_567),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_530),
.B(n_519),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_553),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_597),
.B(n_525),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_567),
.B(n_496),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_554),
.B(n_228),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_553),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_554),
.B(n_496),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_554),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_554),
.B(n_497),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_545),
.B(n_497),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_559),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_545),
.B(n_282),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_559),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_576),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_559),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_581),
.B(n_500),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_545),
.B(n_282),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_541),
.Y(n_748)
);

BUFx4f_ASAP7_75t_L g749 ( 
.A(n_541),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_559),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_565),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_545),
.B(n_282),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_565),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_541),
.B(n_414),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_545),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_553),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_565),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_SL g758 ( 
.A(n_581),
.B(n_427),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_565),
.B(n_500),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_553),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_573),
.B(n_501),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_573),
.A2(n_330),
.B1(n_364),
.B2(n_361),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_627),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_687),
.B(n_573),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_625),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_625),
.B(n_434),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_706),
.A2(n_242),
.B1(n_262),
.B2(n_237),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_687),
.B(n_573),
.Y(n_768)
);

INVx8_ASAP7_75t_L g769 ( 
.A(n_729),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_733),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_684),
.B(n_532),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_692),
.B(n_532),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_733),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_725),
.B(n_535),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_616),
.B(n_617),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_611),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_664),
.B(n_437),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_702),
.B(n_535),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_628),
.A2(n_251),
.B(n_256),
.C(n_241),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_632),
.Y(n_780)
);

AO221x1_ASAP7_75t_L g781 ( 
.A1(n_658),
.A2(n_353),
.B1(n_357),
.B2(n_362),
.C(n_346),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_702),
.B(n_537),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_716),
.B(n_517),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_702),
.B(n_537),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_611),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_622),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_623),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_618),
.B(n_550),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_618),
.B(n_550),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_628),
.B(n_553),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_618),
.B(n_582),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_618),
.B(n_582),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_622),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_716),
.B(n_251),
.C(n_241),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_706),
.A2(n_262),
.B1(n_264),
.B2(n_242),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_637),
.A2(n_454),
.B1(n_257),
.B2(n_268),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_618),
.B(n_582),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_618),
.B(n_582),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_657),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_706),
.A2(n_271),
.B1(n_276),
.B2(n_264),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_618),
.B(n_582),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_746),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_626),
.A2(n_310),
.B1(n_313),
.B2(n_309),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_623),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_632),
.B(n_319),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_628),
.B(n_749),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_635),
.B(n_583),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_635),
.B(n_583),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_729),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_SL g810 ( 
.A(n_690),
.B(n_282),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_636),
.B(n_583),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_749),
.B(n_555),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_740),
.B(n_657),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_749),
.B(n_555),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_740),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_709),
.B(n_555),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_636),
.B(n_583),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_709),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_650),
.B(n_583),
.Y(n_819)
);

INVx8_ASAP7_75t_L g820 ( 
.A(n_729),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_615),
.B(n_279),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_650),
.B(n_587),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_703),
.Y(n_823)
);

AOI221xp5_ASAP7_75t_L g824 ( 
.A1(n_704),
.A2(n_362),
.B1(n_357),
.B2(n_353),
.C(n_370),
.Y(n_824)
);

BUFx5_ASAP7_75t_L g825 ( 
.A(n_703),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_626),
.A2(n_325),
.B1(n_329),
.B2(n_321),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_729),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_641),
.Y(n_828)
);

OR2x6_ASAP7_75t_SL g829 ( 
.A(n_638),
.B(n_283),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_709),
.B(n_555),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_668),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_626),
.B(n_332),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_629),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_643),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_643),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_679),
.B(n_673),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_626),
.A2(n_689),
.B1(n_709),
.B2(n_758),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_652),
.A2(n_556),
.B(n_555),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_674),
.B(n_284),
.Y(n_839)
);

INVx8_ASAP7_75t_L g840 ( 
.A(n_626),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_651),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_626),
.B(n_337),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_755),
.B(n_748),
.Y(n_843)
);

OAI221xp5_ASAP7_75t_L g844 ( 
.A1(n_647),
.A2(n_346),
.B1(n_369),
.B2(n_370),
.C(n_271),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_626),
.A2(n_327),
.B1(n_324),
.B2(n_320),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_620),
.B(n_294),
.C(n_289),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_654),
.B(n_587),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_651),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_663),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_659),
.B(n_295),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_SL g851 ( 
.A(n_721),
.B(n_286),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_724),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_755),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_654),
.B(n_587),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_652),
.B(n_587),
.Y(n_855)
);

AOI22x1_ASAP7_75t_L g856 ( 
.A1(n_748),
.A2(n_256),
.B1(n_339),
.B2(n_359),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_662),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_659),
.B(n_338),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_663),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_689),
.A2(n_335),
.B1(n_324),
.B2(n_320),
.Y(n_860)
);

BUFx8_ASAP7_75t_L g861 ( 
.A(n_672),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_667),
.B(n_555),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_SL g863 ( 
.A(n_721),
.B(n_286),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_667),
.B(n_587),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_726),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_645),
.B(n_640),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_671),
.B(n_501),
.Y(n_867)
);

BUFx4_ASAP7_75t_L g868 ( 
.A(n_682),
.Y(n_868)
);

BUFx5_ASAP7_75t_L g869 ( 
.A(n_730),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_676),
.B(n_555),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_629),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_676),
.B(n_600),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_629),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_678),
.B(n_502),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_689),
.A2(n_335),
.B1(n_303),
.B2(n_291),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_612),
.B(n_502),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_629),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_754),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_683),
.B(n_600),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_621),
.B(n_257),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_683),
.B(n_695),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_695),
.B(n_600),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_666),
.Y(n_883)
);

INVx5_ASAP7_75t_L g884 ( 
.A(n_754),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_697),
.B(n_555),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_697),
.B(n_600),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_691),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_642),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_698),
.B(n_556),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_698),
.B(n_556),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_754),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_613),
.B(n_298),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_701),
.B(n_600),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_666),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_701),
.B(n_578),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_670),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_707),
.B(n_578),
.Y(n_897)
);

INVx8_ASAP7_75t_L g898 ( 
.A(n_689),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_754),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_655),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_707),
.B(n_578),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_712),
.B(n_717),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_737),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_660),
.B(n_299),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_730),
.B(n_556),
.Y(n_905)
);

AOI221xp5_ASAP7_75t_L g906 ( 
.A1(n_647),
.A2(n_336),
.B1(n_340),
.B2(n_327),
.C(n_303),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_661),
.A2(n_339),
.B1(n_318),
.B2(n_311),
.Y(n_907)
);

BUFx5_ASAP7_75t_L g908 ( 
.A(n_689),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_722),
.B(n_728),
.Y(n_909)
);

NOR2x1p5_ASAP7_75t_L g910 ( 
.A(n_665),
.B(n_301),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_677),
.B(n_504),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_715),
.B(n_556),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_689),
.B(n_578),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_715),
.B(n_556),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_734),
.B(n_556),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_689),
.B(n_578),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_739),
.A2(n_268),
.B(n_270),
.C(n_397),
.Y(n_917)
);

AO221x1_ASAP7_75t_L g918 ( 
.A1(n_762),
.A2(n_340),
.B1(n_276),
.B2(n_291),
.C(n_336),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_634),
.B(n_504),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_639),
.B(n_578),
.Y(n_920)
);

NAND2xp33_ASAP7_75t_L g921 ( 
.A(n_735),
.B(n_343),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_670),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_639),
.A2(n_742),
.B1(n_752),
.B2(n_747),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_759),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_639),
.B(n_578),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_614),
.B(n_578),
.Y(n_926)
);

NOR2xp67_ASAP7_75t_L g927 ( 
.A(n_700),
.B(n_507),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_731),
.B(n_507),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_763),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_790),
.A2(n_631),
.B(n_624),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_790),
.A2(n_631),
.B(n_624),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_775),
.B(n_656),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_767),
.A2(n_761),
.B1(n_285),
.B2(n_288),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_L g934 ( 
.A(n_825),
.B(n_735),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_836),
.B(n_738),
.Y(n_935)
);

AO21x1_ASAP7_75t_L g936 ( 
.A1(n_912),
.A2(n_648),
.B(n_285),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_812),
.A2(n_631),
.B(n_624),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_836),
.B(n_738),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_771),
.B(n_743),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_772),
.B(n_743),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_802),
.B(n_745),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_852),
.B(n_508),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_857),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_767),
.A2(n_288),
.B1(n_305),
.B2(n_270),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_802),
.B(n_745),
.Y(n_945)
);

AOI21x1_ASAP7_75t_L g946 ( 
.A1(n_812),
.A2(n_751),
.B(n_750),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_920),
.A2(n_751),
.B(n_750),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_852),
.B(n_633),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_823),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_887),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_876),
.B(n_675),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_839),
.A2(n_720),
.B1(n_719),
.B2(n_693),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_765),
.B(n_508),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_876),
.B(n_675),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_900),
.B(n_681),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_814),
.A2(n_685),
.B(n_681),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_925),
.A2(n_688),
.B(n_685),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_814),
.A2(n_806),
.B(n_909),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_839),
.B(n_688),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_867),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_903),
.B(n_924),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_904),
.B(n_694),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_904),
.B(n_694),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_806),
.A2(n_669),
.B(n_633),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_909),
.A2(n_669),
.B(n_633),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_843),
.A2(n_686),
.B(n_669),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_780),
.B(n_686),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_843),
.A2(n_744),
.B(n_686),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_818),
.A2(n_719),
.B1(n_720),
.B2(n_693),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_766),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_816),
.A2(n_744),
.B(n_649),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_765),
.B(n_520),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_868),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_795),
.A2(n_375),
.B1(n_305),
.B2(n_307),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_796),
.A2(n_696),
.B(n_757),
.C(n_705),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_825),
.B(n_823),
.Y(n_976)
);

AO21x1_ASAP7_75t_L g977 ( 
.A1(n_912),
.A2(n_648),
.B(n_311),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_795),
.B(n_696),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_800),
.A2(n_409),
.B(n_369),
.C(n_380),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_800),
.B(n_705),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_L g981 ( 
.A(n_821),
.B(n_520),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_823),
.Y(n_982)
);

OR2x6_ASAP7_75t_L g983 ( 
.A(n_769),
.B(n_307),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_777),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_816),
.A2(n_744),
.B(n_649),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_830),
.A2(n_792),
.B(n_791),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_823),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_866),
.B(n_708),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_830),
.A2(n_649),
.B(n_646),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_850),
.B(n_858),
.C(n_824),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_797),
.A2(n_649),
.B(n_646),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_853),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_798),
.A2(n_801),
.B(n_789),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_788),
.A2(n_649),
.B(n_646),
.Y(n_994)
);

BUFx4f_ASAP7_75t_L g995 ( 
.A(n_769),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_768),
.B(n_708),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_825),
.B(n_646),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_837),
.A2(n_374),
.B1(n_318),
.B2(n_331),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_844),
.A2(n_711),
.B(n_757),
.C(n_714),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_815),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_855),
.A2(n_736),
.B(n_646),
.Y(n_1001)
);

OR2x2_ASAP7_75t_L g1002 ( 
.A(n_783),
.B(n_523),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_776),
.B(n_711),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_840),
.A2(n_736),
.B(n_619),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_874),
.B(n_523),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_915),
.A2(n_718),
.B(n_714),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_892),
.B(n_525),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_881),
.A2(n_723),
.B(n_718),
.C(n_753),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_785),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_915),
.A2(n_741),
.B(n_723),
.Y(n_1010)
);

CKINVDCx10_ASAP7_75t_R g1011 ( 
.A(n_861),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_878),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_813),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_892),
.B(n_290),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_787),
.B(n_741),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_804),
.B(n_753),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_813),
.B(n_585),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_840),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_850),
.A2(n_314),
.B(n_302),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_764),
.A2(n_619),
.B(n_614),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_884),
.A2(n_891),
.B1(n_899),
.B2(n_923),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_770),
.B(n_614),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_773),
.B(n_619),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_840),
.A2(n_736),
.B(n_653),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_764),
.B(n_630),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_898),
.A2(n_736),
.B(n_653),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_778),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_898),
.A2(n_736),
.B(n_653),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_928),
.B(n_719),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_898),
.A2(n_680),
.B(n_630),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_786),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_774),
.B(n_630),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_782),
.A2(n_784),
.B(n_832),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_825),
.B(n_680),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_884),
.A2(n_359),
.B1(n_331),
.B2(n_351),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_799),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_884),
.A2(n_363),
.B1(n_351),
.B2(n_366),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_809),
.B(n_585),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_928),
.B(n_719),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_825),
.B(n_680),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_906),
.A2(n_821),
.B(n_860),
.C(n_845),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_799),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_842),
.A2(n_710),
.B(n_699),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_902),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_845),
.A2(n_409),
.B(n_418),
.C(n_416),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_825),
.B(n_699),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_833),
.A2(n_710),
.B(n_699),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_881),
.B(n_710),
.Y(n_1048)
);

BUFx12f_ASAP7_75t_L g1049 ( 
.A(n_861),
.Y(n_1049)
);

NOR2xp67_ASAP7_75t_L g1050 ( 
.A(n_827),
.B(n_592),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_914),
.A2(n_366),
.B(n_397),
.C(n_363),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_914),
.A2(n_727),
.B(n_713),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_860),
.A2(n_418),
.B(n_416),
.C(n_406),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_793),
.Y(n_1054)
);

OAI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_810),
.A2(n_863),
.B1(n_851),
.B2(n_783),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_799),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_878),
.A2(n_385),
.B(n_374),
.C(n_375),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_907),
.A2(n_385),
.B(n_377),
.C(n_527),
.Y(n_1058)
);

NOR2xp67_ASAP7_75t_L g1059 ( 
.A(n_846),
.B(n_592),
.Y(n_1059)
);

AOI21x1_ASAP7_75t_L g1060 ( 
.A1(n_905),
.A2(n_527),
.B(n_526),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_783),
.B(n_720),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_833),
.A2(n_877),
.B(n_871),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_807),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_891),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_911),
.A2(n_317),
.B(n_316),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_871),
.A2(n_727),
.B(n_713),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_877),
.A2(n_884),
.B(n_926),
.Y(n_1067)
);

AOI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_805),
.A2(n_377),
.B(n_328),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_808),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_779),
.A2(n_529),
.B(n_552),
.C(n_557),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_799),
.B(n_713),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_873),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_913),
.A2(n_732),
.B(n_727),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_869),
.B(n_732),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_864),
.A2(n_756),
.B(n_732),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_916),
.A2(n_760),
.B(n_756),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_872),
.A2(n_760),
.B(n_756),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_919),
.B(n_595),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_838),
.A2(n_760),
.B(n_562),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_908),
.B(n_621),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_811),
.A2(n_562),
.B(n_563),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_828),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_917),
.A2(n_529),
.B(n_526),
.C(n_527),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_817),
.A2(n_562),
.B(n_563),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_879),
.A2(n_552),
.B(n_557),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_819),
.A2(n_847),
.B(n_822),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_869),
.B(n_720),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_910),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_882),
.A2(n_735),
.B(n_644),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_899),
.A2(n_735),
.B1(n_410),
.B2(n_381),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_L g1091 ( 
.A(n_908),
.B(n_735),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_854),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_886),
.A2(n_563),
.B(n_556),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_834),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_SL g1095 ( 
.A(n_865),
.B(n_290),
.Y(n_1095)
);

INVx11_ASAP7_75t_L g1096 ( 
.A(n_927),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_869),
.B(n_735),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_893),
.A2(n_563),
.B(n_562),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_L g1099 ( 
.A(n_831),
.B(n_404),
.C(n_348),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_869),
.B(n_875),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_794),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_895),
.A2(n_735),
.B(n_644),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_794),
.A2(n_529),
.B(n_526),
.C(n_552),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_888),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_873),
.A2(n_563),
.B(n_562),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_L g1106 ( 
.A(n_769),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_820),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_869),
.B(n_557),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_875),
.A2(n_803),
.B1(n_826),
.B2(n_873),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_873),
.B(n_595),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_897),
.A2(n_563),
.B(n_562),
.Y(n_1111)
);

AOI33xp33_ASAP7_75t_L g1112 ( 
.A1(n_829),
.A2(n_388),
.A3(n_380),
.B1(n_390),
.B2(n_406),
.B3(n_403),
.Y(n_1112)
);

NOR2xp67_ASAP7_75t_L g1113 ( 
.A(n_901),
.B(n_596),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_905),
.A2(n_560),
.B(n_571),
.Y(n_1114)
);

AO21x1_ASAP7_75t_L g1115 ( 
.A1(n_862),
.A2(n_885),
.B(n_870),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_949),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_932),
.B(n_820),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_935),
.B(n_938),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1009),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_932),
.B(n_820),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_960),
.B(n_869),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_990),
.A2(n_1055),
.B(n_1041),
.C(n_1101),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_961),
.B(n_862),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_950),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_935),
.B(n_781),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1055),
.B(n_908),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_990),
.B(n_908),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_938),
.A2(n_856),
.B1(n_849),
.B2(n_896),
.Y(n_1128)
);

OA22x2_ASAP7_75t_L g1129 ( 
.A1(n_1101),
.A2(n_918),
.B1(n_388),
.B2(n_390),
.Y(n_1129)
);

BUFx8_ASAP7_75t_SL g1130 ( 
.A(n_1049),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_949),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_960),
.B(n_870),
.Y(n_1132)
);

OAI21xp33_ASAP7_75t_SL g1133 ( 
.A1(n_1100),
.A2(n_885),
.B(n_889),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_934),
.A2(n_908),
.B(n_921),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_949),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_1014),
.B(n_415),
.C(n_322),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_929),
.B(n_908),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_984),
.A2(n_411),
.B1(n_379),
.B2(n_347),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_929),
.B(n_835),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1044),
.B(n_841),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1107),
.B(n_848),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_970),
.B(n_889),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_949),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1013),
.B(n_859),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1011),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1007),
.B(n_883),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1041),
.A2(n_922),
.B(n_894),
.C(n_890),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_982),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1027),
.A2(n_890),
.B(n_403),
.C(n_596),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1072),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_956),
.A2(n_880),
.B(n_560),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_943),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_944),
.A2(n_290),
.B1(n_392),
.B2(n_345),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1099),
.A2(n_1029),
.B1(n_1039),
.B2(n_981),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_974),
.A2(n_290),
.B1(n_392),
.B2(n_349),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_988),
.B(n_1005),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_988),
.B(n_597),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_993),
.A2(n_880),
.B(n_562),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_986),
.A2(n_373),
.B(n_376),
.C(n_378),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_941),
.B(n_597),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_1056),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1019),
.B(n_334),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1029),
.A2(n_356),
.B1(n_354),
.B2(n_352),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1018),
.B(n_621),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1033),
.A2(n_562),
.B(n_563),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_945),
.B(n_598),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1000),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1012),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_SL g1169 ( 
.A(n_1065),
.B(n_371),
.C(n_372),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_1012),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_948),
.B(n_598),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1068),
.A2(n_958),
.B(n_948),
.C(n_1039),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_R g1173 ( 
.A(n_995),
.B(n_383),
.Y(n_1173)
);

AOI21x1_ASAP7_75t_L g1174 ( 
.A1(n_946),
.A2(n_560),
.B(n_599),
.Y(n_1174)
);

INVxp67_ASAP7_75t_SL g1175 ( 
.A(n_982),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_939),
.B(n_598),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1104),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1056),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_940),
.B(n_601),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_SL g1180 ( 
.A(n_1018),
.B(n_621),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_953),
.B(n_384),
.Y(n_1181)
);

O2A1O1Ixp5_ASAP7_75t_L g1182 ( 
.A1(n_936),
.A2(n_606),
.B(n_601),
.C(n_607),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1013),
.B(n_601),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1056),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1091),
.A2(n_563),
.B(n_621),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_976),
.A2(n_644),
.B(n_621),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_978),
.A2(n_980),
.B1(n_1018),
.B2(n_959),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1057),
.A2(n_607),
.B(n_606),
.C(n_572),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1051),
.A2(n_606),
.B(n_607),
.C(n_407),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1064),
.Y(n_1190)
);

CKINVDCx16_ASAP7_75t_R g1191 ( 
.A(n_1095),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_972),
.B(n_392),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1064),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_976),
.A2(n_644),
.B(n_609),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_L g1195 ( 
.A(n_1088),
.B(n_90),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_987),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1040),
.A2(n_644),
.B(n_609),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1003),
.Y(n_1198)
);

AOI21xp33_ASAP7_75t_L g1199 ( 
.A1(n_998),
.A2(n_394),
.B(n_399),
.Y(n_1199)
);

NAND2x1_ASAP7_75t_L g1200 ( 
.A(n_1036),
.B(n_580),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1018),
.A2(n_401),
.B1(n_408),
.B2(n_571),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1099),
.A2(n_572),
.B(n_599),
.C(n_580),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_997),
.A2(n_644),
.B(n_609),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1056),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_933),
.A2(n_392),
.B1(n_608),
.B2(n_602),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1031),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1021),
.A2(n_609),
.B1(n_608),
.B2(n_580),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_997),
.A2(n_602),
.B(n_599),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_973),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1072),
.Y(n_1210)
);

AOI21x1_ASAP7_75t_L g1211 ( 
.A1(n_962),
.A2(n_608),
.B(n_602),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1054),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1017),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1063),
.B(n_580),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_SL g1215 ( 
.A(n_1112),
.B(n_588),
.Y(n_1215)
);

AO21x1_ASAP7_75t_L g1216 ( 
.A1(n_963),
.A2(n_608),
.B(n_602),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1015),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_942),
.B(n_1017),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1016),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1038),
.B(n_591),
.Y(n_1220)
);

AO21x2_ASAP7_75t_L g1221 ( 
.A1(n_947),
.A2(n_599),
.B(n_591),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1074),
.A2(n_591),
.B(n_588),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1069),
.B(n_591),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1082),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1094),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1038),
.B(n_172),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1022),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_992),
.B(n_17),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_951),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1092),
.B(n_603),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1034),
.A2(n_588),
.B(n_603),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1002),
.B(n_955),
.Y(n_1232)
);

NOR2x1_ASAP7_75t_R g1233 ( 
.A(n_1036),
.B(n_603),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1078),
.B(n_603),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1034),
.A2(n_588),
.B(n_603),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1060),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_983),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1046),
.A2(n_588),
.B(n_603),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1059),
.A2(n_603),
.B(n_588),
.C(n_25),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1046),
.A2(n_603),
.B(n_588),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_954),
.A2(n_588),
.B1(n_207),
.B2(n_204),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1109),
.A2(n_17),
.B1(n_22),
.B2(n_28),
.Y(n_1242)
);

AOI221x1_ASAP7_75t_L g1243 ( 
.A1(n_1035),
.A2(n_22),
.B1(n_28),
.B2(n_30),
.C(n_33),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_967),
.B(n_30),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_967),
.B(n_33),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_979),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1061),
.B(n_38),
.Y(n_1247)
);

CKINVDCx8_ASAP7_75t_R g1248 ( 
.A(n_983),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1032),
.B(n_39),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1078),
.B(n_91),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1023),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1061),
.B(n_39),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_930),
.A2(n_94),
.B(n_202),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_995),
.B(n_203),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1096),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_931),
.A2(n_190),
.B(n_189),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_937),
.A2(n_187),
.B(n_185),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1072),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_952),
.A2(n_180),
.B1(n_178),
.B2(n_175),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_979),
.B(n_40),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1110),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1114),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1106),
.B(n_174),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_983),
.B(n_41),
.Y(n_1264)
);

OR2x6_ASAP7_75t_L g1265 ( 
.A(n_1042),
.B(n_167),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_996),
.B(n_41),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_994),
.A2(n_159),
.B(n_153),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1050),
.B(n_1042),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1037),
.A2(n_42),
.A3(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1086),
.A2(n_152),
.B(n_150),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1110),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1087),
.A2(n_140),
.B(n_139),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_999),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_991),
.A2(n_133),
.B(n_132),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1048),
.B(n_44),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1122),
.A2(n_1058),
.B(n_1113),
.C(n_975),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1118),
.B(n_1045),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1168),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1162),
.A2(n_1090),
.B(n_1106),
.C(n_1067),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1136),
.A2(n_1045),
.B(n_1053),
.C(n_1103),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1165),
.A2(n_1085),
.B(n_1043),
.Y(n_1281)
);

NOR2xp67_ASAP7_75t_L g1282 ( 
.A(n_1120),
.B(n_1071),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1156),
.A2(n_969),
.B1(n_1108),
.B2(n_1097),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1247),
.A2(n_1115),
.B1(n_977),
.B2(n_1072),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1232),
.B(n_1053),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1125),
.A2(n_1070),
.B(n_1083),
.C(n_1025),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1213),
.B(n_1020),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1116),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1116),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1232),
.B(n_957),
.Y(n_1290)
);

AOI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1211),
.A2(n_965),
.B(n_1079),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1134),
.A2(n_964),
.B(n_1028),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1229),
.B(n_1076),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1191),
.B(n_1052),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1117),
.B(n_971),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1229),
.B(n_1073),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1124),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1145),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1120),
.A2(n_1077),
.B1(n_1075),
.B2(n_1102),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1244),
.A2(n_1008),
.B(n_985),
.C(n_968),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1177),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1242),
.A2(n_1089),
.B(n_1062),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1192),
.B(n_1006),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1130),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1216),
.A2(n_966),
.A3(n_1001),
.B(n_1084),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1172),
.A2(n_1010),
.B(n_1080),
.C(n_989),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1247),
.A2(n_1080),
.B1(n_1111),
.B2(n_1066),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1182),
.A2(n_1081),
.B(n_1098),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1275),
.A2(n_1093),
.B(n_1047),
.C(n_1030),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1127),
.A2(n_1026),
.B(n_1024),
.Y(n_1310)
);

AOI221x1_ASAP7_75t_L g1311 ( 
.A1(n_1270),
.A2(n_1105),
.B1(n_1004),
.B2(n_50),
.C(n_51),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1154),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1174),
.A2(n_126),
.B(n_122),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1170),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1167),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1209),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1187),
.A2(n_1126),
.B(n_1158),
.Y(n_1317)
);

O2A1O1Ixp5_ASAP7_75t_SL g1318 ( 
.A1(n_1207),
.A2(n_52),
.B(n_54),
.C(n_55),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1116),
.Y(n_1319)
);

AOI221x1_ASAP7_75t_L g1320 ( 
.A1(n_1252),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.C(n_63),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1151),
.A2(n_120),
.B(n_70),
.Y(n_1321)
);

AO32x2_ASAP7_75t_L g1322 ( 
.A1(n_1128),
.A2(n_67),
.A3(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1133),
.A2(n_67),
.B(n_76),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1198),
.B(n_78),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1189),
.A2(n_78),
.A3(n_80),
.B(n_1147),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1170),
.Y(n_1326)
);

AOI221x1_ASAP7_75t_L g1327 ( 
.A1(n_1245),
.A2(n_1259),
.B1(n_1275),
.B2(n_1159),
.C(n_1239),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1242),
.A2(n_1181),
.B1(n_1228),
.B2(n_1142),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1255),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1222),
.A2(n_1208),
.B(n_1240),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1236),
.A2(n_1243),
.A3(n_1262),
.B(n_1273),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1231),
.A2(n_1235),
.B(n_1238),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1213),
.B(n_1218),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1197),
.A2(n_1194),
.B(n_1203),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1171),
.A2(n_1121),
.A3(n_1241),
.B(n_1149),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_1173),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1146),
.A2(n_1157),
.B(n_1179),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1169),
.B(n_1199),
.C(n_1155),
.Y(n_1338)
);

BUFx8_ASAP7_75t_L g1339 ( 
.A(n_1237),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1249),
.A2(n_1266),
.B(n_1230),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1217),
.B(n_1219),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1176),
.A2(n_1123),
.B(n_1160),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1248),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1185),
.A2(n_1253),
.B(n_1256),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1261),
.B(n_1227),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1166),
.A2(n_1137),
.B(n_1223),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1169),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1221),
.A2(n_1257),
.B(n_1214),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1261),
.B(n_1251),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1140),
.B(n_1132),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1221),
.A2(n_1135),
.B(n_1121),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1135),
.A2(n_1234),
.B(n_1164),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1132),
.A2(n_1274),
.A3(n_1267),
.B(n_1228),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_1129),
.B2(n_1271),
.Y(n_1354)
);

BUFx12f_ASAP7_75t_L g1355 ( 
.A(n_1264),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1246),
.A2(n_1152),
.B(n_1226),
.C(n_1225),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1175),
.B(n_1148),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1164),
.A2(n_1233),
.B(n_1250),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1200),
.A2(n_1186),
.B(n_1144),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1272),
.A2(n_1202),
.B(n_1150),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1260),
.A2(n_1155),
.B(n_1153),
.C(n_1220),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1148),
.B(n_1193),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1153),
.A2(n_1220),
.B1(n_1163),
.B2(n_1206),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1141),
.B(n_1138),
.Y(n_1364)
);

CKINVDCx14_ASAP7_75t_R g1365 ( 
.A(n_1265),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1190),
.B(n_1193),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1183),
.A2(n_1224),
.B(n_1212),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1141),
.B(n_1268),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1150),
.A2(n_1258),
.B(n_1210),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1190),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1175),
.A2(n_1263),
.B(n_1254),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_L g1372 ( 
.A(n_1188),
.B(n_1201),
.C(n_1139),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_SL g1373 ( 
.A1(n_1204),
.A2(n_1196),
.B(n_1258),
.C(n_1210),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1268),
.B(n_1204),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1180),
.A2(n_1265),
.B(n_1178),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1161),
.B(n_1265),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1205),
.B(n_1195),
.C(n_1161),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1131),
.A2(n_1143),
.B(n_1178),
.Y(n_1378)
);

CKINVDCx16_ASAP7_75t_R g1379 ( 
.A(n_1131),
.Y(n_1379)
);

INVxp67_ASAP7_75t_SL g1380 ( 
.A(n_1131),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1205),
.A2(n_1129),
.B(n_1269),
.C(n_1143),
.Y(n_1381)
);

OR2x6_ASAP7_75t_L g1382 ( 
.A(n_1131),
.B(n_1143),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1269),
.A2(n_1143),
.A3(n_1178),
.B(n_1184),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1178),
.Y(n_1384)
);

AOI211x1_ASAP7_75t_L g1385 ( 
.A1(n_1269),
.A2(n_1118),
.B(n_1125),
.C(n_844),
.Y(n_1385)
);

AO21x2_ASAP7_75t_L g1386 ( 
.A1(n_1269),
.A2(n_1216),
.B(n_1172),
.Y(n_1386)
);

AOI221x1_ASAP7_75t_L g1387 ( 
.A1(n_1184),
.A2(n_990),
.B1(n_1118),
.B2(n_1270),
.C(n_1172),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1184),
.A2(n_1134),
.B(n_934),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1184),
.B(n_1055),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1116),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1168),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_SL g1392 ( 
.A1(n_1118),
.A2(n_1041),
.B(n_1126),
.C(n_775),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1134),
.A2(n_934),
.B(n_898),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1118),
.A2(n_810),
.B1(n_863),
.B2(n_851),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1117),
.B(n_775),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1216),
.A2(n_977),
.A3(n_936),
.B(n_1187),
.Y(n_1396)
);

AOI221x1_ASAP7_75t_L g1397 ( 
.A1(n_1118),
.A2(n_990),
.B1(n_1270),
.B2(n_1172),
.C(n_1187),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1165),
.A2(n_1174),
.B(n_1151),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1192),
.B(n_777),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1168),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1216),
.A2(n_977),
.A3(n_936),
.B(n_1187),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1165),
.A2(n_1174),
.B(n_1151),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1118),
.B(n_836),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1213),
.B(n_627),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1191),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1119),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1134),
.A2(n_934),
.B(n_898),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1213),
.B(n_1107),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1165),
.A2(n_1174),
.B(n_1151),
.Y(n_1409)
);

AO32x2_ASAP7_75t_L g1410 ( 
.A1(n_1187),
.A2(n_974),
.A3(n_944),
.B1(n_796),
.B2(n_998),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1168),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1118),
.B(n_836),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1165),
.A2(n_1174),
.B(n_1151),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1133),
.A2(n_1122),
.B(n_1118),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1265),
.B(n_769),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1116),
.Y(n_1416)
);

OAI22x1_ASAP7_75t_L g1417 ( 
.A1(n_1120),
.A2(n_932),
.B1(n_775),
.B2(n_1117),
.Y(n_1417)
);

BUFx2_ASAP7_75t_SL g1418 ( 
.A(n_1124),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_SL g1419 ( 
.A1(n_1118),
.A2(n_1041),
.B(n_1126),
.C(n_775),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1116),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1165),
.A2(n_1174),
.B(n_1151),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1216),
.A2(n_977),
.A3(n_936),
.B(n_1187),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1119),
.Y(n_1423)
);

AOI211x1_ASAP7_75t_L g1424 ( 
.A1(n_1118),
.A2(n_1125),
.B(n_844),
.C(n_961),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1134),
.A2(n_934),
.B(n_898),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1216),
.A2(n_1182),
.B(n_1172),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1134),
.A2(n_934),
.B(n_898),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1119),
.Y(n_1428)
);

AOI211x1_ASAP7_75t_L g1429 ( 
.A1(n_1118),
.A2(n_1125),
.B(n_844),
.C(n_961),
.Y(n_1429)
);

OR2x6_ASAP7_75t_L g1430 ( 
.A(n_1265),
.B(n_769),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1168),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1134),
.A2(n_934),
.B(n_898),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1213),
.B(n_1107),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1119),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1172),
.A2(n_775),
.B(n_836),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1119),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1118),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1119),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1117),
.B(n_775),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1118),
.A2(n_775),
.B1(n_836),
.B2(n_1156),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1122),
.A2(n_836),
.B(n_990),
.C(n_932),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1328),
.A2(n_1403),
.B1(n_1412),
.B2(n_1437),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1382),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1362),
.B(n_1391),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1298),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1301),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1328),
.A2(n_1437),
.B1(n_1320),
.B2(n_1338),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1406),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1338),
.A2(n_1394),
.B(n_1441),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1440),
.A2(n_1385),
.B1(n_1395),
.B2(n_1439),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1428),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1417),
.A2(n_1312),
.B1(n_1435),
.B2(n_1399),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1329),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1434),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1414),
.A2(n_1323),
.B1(n_1347),
.B2(n_1389),
.Y(n_1455)
);

NAND2x1p5_ASAP7_75t_L g1456 ( 
.A(n_1366),
.B(n_1370),
.Y(n_1456)
);

CKINVDCx11_ASAP7_75t_R g1457 ( 
.A(n_1336),
.Y(n_1457)
);

BUFx4f_ASAP7_75t_SL g1458 ( 
.A(n_1297),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_1304),
.Y(n_1459)
);

INVx6_ASAP7_75t_L g1460 ( 
.A(n_1379),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1405),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1288),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1311),
.A2(n_1323),
.B1(n_1341),
.B2(n_1414),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1357),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_SL g1465 ( 
.A1(n_1365),
.A2(n_1303),
.B1(n_1285),
.B2(n_1377),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1333),
.A2(n_1418),
.B1(n_1343),
.B2(n_1376),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_1339),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1339),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1377),
.A2(n_1405),
.B1(n_1430),
.B2(n_1415),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1324),
.A2(n_1350),
.B1(n_1277),
.B2(n_1397),
.Y(n_1470)
);

INVx6_ASAP7_75t_L g1471 ( 
.A(n_1368),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1294),
.A2(n_1372),
.B1(n_1364),
.B2(n_1287),
.Y(n_1472)
);

INVx4_ASAP7_75t_L g1473 ( 
.A(n_1382),
.Y(n_1473)
);

INVx6_ASAP7_75t_L g1474 ( 
.A(n_1368),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1282),
.A2(n_1415),
.B1(n_1430),
.B2(n_1355),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1288),
.Y(n_1476)
);

BUFx12f_ASAP7_75t_L g1477 ( 
.A(n_1404),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1415),
.A2(n_1430),
.B1(n_1290),
.B2(n_1322),
.Y(n_1478)
);

BUFx10_ASAP7_75t_L g1479 ( 
.A(n_1408),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1315),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1374),
.Y(n_1481)
);

INVx8_ASAP7_75t_L g1482 ( 
.A(n_1382),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1282),
.A2(n_1363),
.B1(n_1361),
.B2(n_1372),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1322),
.A2(n_1386),
.B1(n_1342),
.B2(n_1436),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1431),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1316),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1278),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1322),
.A2(n_1386),
.B1(n_1438),
.B2(n_1423),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1287),
.A2(n_1411),
.B1(n_1400),
.B2(n_1371),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1314),
.Y(n_1490)
);

CKINVDCx6p67_ASAP7_75t_R g1491 ( 
.A(n_1431),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1385),
.A2(n_1429),
.B1(n_1424),
.B2(n_1381),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1354),
.A2(n_1345),
.B1(n_1349),
.B2(n_1387),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1354),
.A2(n_1295),
.B1(n_1296),
.B2(n_1293),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1319),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1326),
.A2(n_1433),
.B1(n_1408),
.B2(n_1284),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1367),
.Y(n_1497)
);

INVx6_ASAP7_75t_L g1498 ( 
.A(n_1374),
.Y(n_1498)
);

BUFx10_ASAP7_75t_L g1499 ( 
.A(n_1433),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1392),
.A2(n_1419),
.B1(n_1283),
.B2(n_1337),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1319),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1340),
.A2(n_1317),
.B1(n_1299),
.B2(n_1346),
.Y(n_1502)
);

INVx6_ASAP7_75t_L g1503 ( 
.A(n_1319),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1327),
.A2(n_1299),
.B1(n_1302),
.B2(n_1307),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1424),
.A2(n_1429),
.B1(n_1356),
.B2(n_1276),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1340),
.A2(n_1358),
.B1(n_1426),
.B2(n_1307),
.Y(n_1506)
);

OAI21xp33_ASAP7_75t_L g1507 ( 
.A1(n_1280),
.A2(n_1279),
.B(n_1302),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1384),
.B(n_1380),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1331),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1384),
.B(n_1420),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1331),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1375),
.A2(n_1300),
.B1(n_1351),
.B2(n_1352),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1390),
.Y(n_1513)
);

INVx8_ASAP7_75t_L g1514 ( 
.A(n_1390),
.Y(n_1514)
);

BUFx8_ASAP7_75t_L g1515 ( 
.A(n_1390),
.Y(n_1515)
);

CKINVDCx14_ASAP7_75t_R g1516 ( 
.A(n_1289),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1373),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1416),
.A2(n_1420),
.B1(n_1310),
.B2(n_1426),
.Y(n_1518)
);

CKINVDCx6p67_ASAP7_75t_R g1519 ( 
.A(n_1416),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1348),
.A2(n_1360),
.B1(n_1321),
.B2(n_1308),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1369),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1348),
.A2(n_1308),
.B1(n_1388),
.B2(n_1359),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1378),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1313),
.B(n_1344),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1410),
.A2(n_1383),
.B1(n_1318),
.B2(n_1432),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1334),
.A2(n_1292),
.B1(n_1330),
.B2(n_1332),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1398),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1383),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1393),
.A2(n_1425),
.B1(n_1407),
.B2(n_1427),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1325),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1402),
.A2(n_1409),
.B1(n_1413),
.B2(n_1421),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1306),
.Y(n_1532)
);

INVx6_ASAP7_75t_L g1533 ( 
.A(n_1286),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1281),
.A2(n_1410),
.B1(n_1353),
.B2(n_1335),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1383),
.A2(n_1353),
.B1(n_1335),
.B2(n_1309),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1353),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1291),
.A2(n_1335),
.B1(n_1396),
.B2(n_1401),
.Y(n_1537)
);

INVx6_ASAP7_75t_L g1538 ( 
.A(n_1396),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1396),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1422),
.A2(n_1305),
.B1(n_1401),
.B2(n_546),
.Y(n_1540)
);

INVx6_ASAP7_75t_L g1541 ( 
.A(n_1401),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1422),
.A2(n_990),
.B1(n_1338),
.B2(n_932),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1422),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1305),
.A2(n_990),
.B1(n_1338),
.B2(n_932),
.Y(n_1544)
);

INVx6_ASAP7_75t_L g1545 ( 
.A(n_1379),
.Y(n_1545)
);

BUFx12f_ASAP7_75t_L g1546 ( 
.A(n_1304),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1406),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1338),
.A2(n_546),
.B1(n_810),
.B2(n_851),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1552)
);

BUFx2_ASAP7_75t_SL g1553 ( 
.A(n_1316),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1301),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1328),
.A2(n_1437),
.B1(n_1118),
.B2(n_1320),
.Y(n_1556)
);

CKINVDCx6p67_ASAP7_75t_R g1557 ( 
.A(n_1298),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1406),
.Y(n_1558)
);

INVx8_ASAP7_75t_L g1559 ( 
.A(n_1382),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1301),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1406),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1328),
.A2(n_1118),
.B1(n_1242),
.B2(n_1403),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1338),
.A2(n_546),
.B1(n_810),
.B2(n_851),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1379),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1336),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1328),
.A2(n_1118),
.B1(n_1242),
.B2(n_1403),
.Y(n_1567)
);

INVx8_ASAP7_75t_L g1568 ( 
.A(n_1382),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1569)
);

OAI22x1_ASAP7_75t_L g1570 ( 
.A1(n_1328),
.A2(n_1437),
.B1(n_1338),
.B2(n_1395),
.Y(n_1570)
);

BUFx4f_ASAP7_75t_L g1571 ( 
.A(n_1298),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1406),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1399),
.B(n_777),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1304),
.Y(n_1574)
);

OAI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1328),
.A2(n_1437),
.B1(n_1118),
.B2(n_1320),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1406),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1406),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1379),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1406),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1406),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1405),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1582)
);

BUFx12f_ASAP7_75t_L g1583 ( 
.A(n_1304),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1406),
.Y(n_1584)
);

BUFx12f_ASAP7_75t_L g1585 ( 
.A(n_1304),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1301),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1338),
.A2(n_990),
.B1(n_932),
.B2(n_775),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_SL g1588 ( 
.A1(n_1336),
.A2(n_1191),
.B1(n_656),
.B2(n_932),
.Y(n_1588)
);

BUFx4f_ASAP7_75t_SL g1589 ( 
.A(n_1329),
.Y(n_1589)
);

BUFx10_ASAP7_75t_L g1590 ( 
.A(n_1304),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1406),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1406),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1406),
.Y(n_1593)
);

NAND2x1p5_ASAP7_75t_L g1594 ( 
.A(n_1443),
.B(n_1517),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1509),
.Y(n_1595)
);

AOI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1570),
.A2(n_1512),
.B(n_1530),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1443),
.Y(n_1597)
);

NAND2x1p5_ASAP7_75t_L g1598 ( 
.A(n_1443),
.B(n_1518),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1511),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1527),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1528),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1536),
.Y(n_1602)
);

NAND2x1_ASAP7_75t_L g1603 ( 
.A(n_1533),
.B(n_1521),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1543),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1544),
.B(n_1542),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1524),
.A2(n_1531),
.B(n_1522),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1475),
.B(n_1443),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1540),
.B(n_1478),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1527),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1540),
.B(n_1478),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1549),
.B(n_1550),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1538),
.Y(n_1612)
);

NAND2x1p5_ASAP7_75t_L g1613 ( 
.A(n_1483),
.B(n_1473),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1456),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1541),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1534),
.A2(n_1507),
.B(n_1506),
.Y(n_1616)
);

AO21x2_ASAP7_75t_L g1617 ( 
.A1(n_1537),
.A2(n_1504),
.B(n_1463),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1532),
.B(n_1473),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1541),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1539),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1488),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1488),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1532),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1457),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1551),
.B(n_1552),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1492),
.B(n_1484),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1554),
.A2(n_1569),
.B(n_1565),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1524),
.A2(n_1529),
.B(n_1512),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1485),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1477),
.B(n_1588),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1464),
.B(n_1480),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1484),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1444),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1548),
.A2(n_1563),
.B1(n_1455),
.B2(n_1587),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1497),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1537),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1535),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1508),
.Y(n_1638)
);

AO22x1_ASAP7_75t_L g1639 ( 
.A1(n_1450),
.A2(n_1567),
.B1(n_1562),
.B2(n_1442),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1535),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1505),
.Y(n_1641)
);

AO21x2_ASAP7_75t_L g1642 ( 
.A1(n_1504),
.A2(n_1463),
.B(n_1447),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1482),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1505),
.Y(n_1644)
);

NOR2xp67_ASAP7_75t_R g1645 ( 
.A(n_1533),
.B(n_1468),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1548),
.A2(n_1563),
.B(n_1449),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1533),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_SL g1648 ( 
.A1(n_1562),
.A2(n_1567),
.B1(n_1442),
.B2(n_1466),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1593),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1582),
.B(n_1470),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1592),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1547),
.Y(n_1653)
);

AO21x2_ASAP7_75t_L g1654 ( 
.A1(n_1447),
.A2(n_1556),
.B(n_1575),
.Y(n_1654)
);

INVx5_ASAP7_75t_SL g1655 ( 
.A(n_1491),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1520),
.A2(n_1526),
.B(n_1502),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1591),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1558),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1561),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1523),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1494),
.B(n_1465),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1460),
.A2(n_1545),
.B1(n_1564),
.B2(n_1578),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1573),
.B(n_1486),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1559),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1572),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1490),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1576),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1510),
.Y(n_1668)
);

AO21x1_ASAP7_75t_L g1669 ( 
.A1(n_1556),
.A2(n_1575),
.B(n_1470),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1577),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1580),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1584),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1472),
.A2(n_1452),
.B(n_1489),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1465),
.B(n_1525),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1525),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1500),
.A2(n_1493),
.B(n_1469),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1448),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1579),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1487),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1446),
.B(n_1586),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1568),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1568),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1500),
.A2(n_1493),
.B(n_1469),
.Y(n_1683)
);

AOI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1513),
.A2(n_1581),
.B(n_1461),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1496),
.B(n_1578),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1476),
.A2(n_1519),
.B(n_1515),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1471),
.A2(n_1474),
.B1(n_1555),
.B2(n_1560),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1462),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1515),
.A2(n_1516),
.B(n_1514),
.Y(n_1689)
);

AO21x1_ASAP7_75t_SL g1690 ( 
.A1(n_1514),
.A2(n_1503),
.B(n_1481),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1471),
.A2(n_1474),
.B1(n_1545),
.B2(n_1460),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1481),
.B(n_1498),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1481),
.B(n_1498),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1498),
.B(n_1474),
.Y(n_1694)
);

NAND2x1p5_ASAP7_75t_L g1695 ( 
.A(n_1495),
.B(n_1501),
.Y(n_1695)
);

BUFx2_ASAP7_75t_SL g1696 ( 
.A(n_1479),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1479),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1503),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1514),
.A2(n_1503),
.B(n_1499),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1471),
.B(n_1553),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1458),
.A2(n_1566),
.B1(n_1467),
.B2(n_1589),
.Y(n_1701)
);

OAI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1646),
.A2(n_1453),
.B(n_1445),
.C(n_1459),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1638),
.B(n_1557),
.Y(n_1703)
);

AO21x1_ASAP7_75t_L g1704 ( 
.A1(n_1683),
.A2(n_1571),
.B(n_1590),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1668),
.B(n_1571),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1676),
.A2(n_1590),
.B(n_1574),
.C(n_1583),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1633),
.B(n_1546),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1685),
.B(n_1585),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1689),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1634),
.A2(n_1648),
.B1(n_1625),
.B2(n_1611),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1637),
.B(n_1640),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1598),
.B(n_1639),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1620),
.B(n_1631),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1647),
.B(n_1650),
.Y(n_1714)
);

OA21x2_ASAP7_75t_L g1715 ( 
.A1(n_1628),
.A2(n_1656),
.B(n_1669),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1660),
.B(n_1629),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1669),
.A2(n_1627),
.B1(n_1654),
.B2(n_1642),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1661),
.A2(n_1673),
.B(n_1605),
.C(n_1674),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1640),
.B(n_1632),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1673),
.A2(n_1661),
.B(n_1605),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1639),
.A2(n_1642),
.B1(n_1654),
.B2(n_1674),
.C(n_1621),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1654),
.A2(n_1642),
.B(n_1647),
.C(n_1613),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1647),
.B(n_1613),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1647),
.B(n_1613),
.Y(n_1724)
);

OA21x2_ASAP7_75t_L g1725 ( 
.A1(n_1628),
.A2(n_1656),
.B(n_1606),
.Y(n_1725)
);

NAND4xp25_ASAP7_75t_L g1726 ( 
.A(n_1630),
.B(n_1641),
.C(n_1644),
.D(n_1687),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1621),
.A2(n_1622),
.B1(n_1608),
.B2(n_1610),
.C(n_1632),
.Y(n_1727)
);

AO32x2_ASAP7_75t_L g1728 ( 
.A1(n_1614),
.A2(n_1691),
.A3(n_1597),
.B1(n_1617),
.B2(n_1622),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1617),
.A2(n_1596),
.B(n_1636),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1595),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1662),
.A2(n_1655),
.B1(n_1679),
.B2(n_1641),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_SL g1732 ( 
.A(n_1623),
.B(n_1690),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1655),
.A2(n_1679),
.B1(n_1644),
.B2(n_1666),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1663),
.A2(n_1684),
.B(n_1623),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1618),
.B(n_1684),
.Y(n_1735)
);

OA21x2_ASAP7_75t_L g1736 ( 
.A1(n_1636),
.A2(n_1599),
.B(n_1595),
.Y(n_1736)
);

NAND4xp25_ASAP7_75t_L g1737 ( 
.A(n_1675),
.B(n_1651),
.C(n_1672),
.D(n_1671),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1626),
.B(n_1608),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1607),
.B(n_1612),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1635),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1607),
.B(n_1612),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_R g1742 ( 
.A(n_1624),
.B(n_1645),
.Y(n_1742)
);

OAI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1610),
.A2(n_1675),
.B(n_1626),
.C(n_1616),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1653),
.B(n_1667),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1616),
.B(n_1667),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1603),
.A2(n_1643),
.B(n_1664),
.C(n_1686),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1700),
.A2(n_1686),
.B(n_1598),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1599),
.A2(n_1602),
.B(n_1601),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1615),
.B(n_1619),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1677),
.B(n_1671),
.C(n_1652),
.Y(n_1750)
);

BUFx4f_ASAP7_75t_SL g1751 ( 
.A(n_1688),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1616),
.B(n_1635),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1649),
.B(n_1652),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1649),
.B(n_1657),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1658),
.B(n_1670),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1643),
.A2(n_1664),
.B(n_1689),
.C(n_1699),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1747),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1704),
.B(n_1697),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1748),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1750),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1748),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1707),
.B(n_1680),
.Y(n_1762)
);

NAND2xp33_ASAP7_75t_SL g1763 ( 
.A(n_1710),
.B(n_1708),
.Y(n_1763)
);

OAI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1717),
.A2(n_1701),
.B1(n_1692),
.B2(n_1693),
.C(n_1598),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1709),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1719),
.B(n_1665),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1745),
.Y(n_1767)
);

NOR2x1_ASAP7_75t_SL g1768 ( 
.A(n_1712),
.B(n_1743),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1720),
.A2(n_1682),
.B1(n_1681),
.B2(n_1694),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1711),
.B(n_1659),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1730),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1745),
.B(n_1604),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1739),
.B(n_1615),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1730),
.Y(n_1774)
);

INVx4_ASAP7_75t_L g1775 ( 
.A(n_1751),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1713),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1721),
.A2(n_1655),
.B1(n_1594),
.B2(n_1677),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1739),
.B(n_1741),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1741),
.B(n_1604),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1740),
.Y(n_1780)
);

OR2x2_ASAP7_75t_L g1781 ( 
.A(n_1752),
.B(n_1609),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1734),
.B(n_1697),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1753),
.B(n_1678),
.Y(n_1783)
);

NAND2x1_ASAP7_75t_L g1784 ( 
.A(n_1712),
.B(n_1597),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1735),
.Y(n_1785)
);

INVx4_ASAP7_75t_L g1786 ( 
.A(n_1751),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1756),
.B(n_1600),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1763),
.A2(n_1727),
.B1(n_1718),
.B2(n_1738),
.C(n_1722),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1760),
.B(n_1716),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1765),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1767),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1761),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1761),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1778),
.B(n_1728),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1771),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1785),
.B(n_1728),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1777),
.A2(n_1718),
.B1(n_1738),
.B2(n_1706),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1761),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1785),
.B(n_1728),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_SL g1800 ( 
.A(n_1775),
.B(n_1742),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1757),
.B(n_1702),
.C(n_1706),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1757),
.A2(n_1714),
.B1(n_1726),
.B2(n_1737),
.C(n_1735),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1774),
.B(n_1729),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1774),
.B(n_1754),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1780),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1785),
.B(n_1728),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_L g1807 ( 
.A(n_1782),
.B(n_1714),
.C(n_1715),
.Y(n_1807)
);

NAND4xp25_ASAP7_75t_SL g1808 ( 
.A(n_1769),
.B(n_1746),
.C(n_1756),
.D(n_1705),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1776),
.Y(n_1809)
);

NAND5xp2_ASAP7_75t_L g1810 ( 
.A(n_1764),
.B(n_1746),
.C(n_1723),
.D(n_1724),
.E(n_1594),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1766),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1787),
.B(n_1749),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1767),
.B(n_1736),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1777),
.A2(n_1731),
.B(n_1724),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1787),
.B(n_1765),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1767),
.B(n_1736),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1762),
.B(n_1703),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1780),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1780),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1781),
.B(n_1736),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1768),
.A2(n_1712),
.B(n_1732),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1758),
.A2(n_1715),
.B(n_1723),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1773),
.B(n_1715),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1784),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1781),
.B(n_1744),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1783),
.B(n_1755),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1813),
.B(n_1759),
.Y(n_1827)
);

NAND2x1p5_ASAP7_75t_L g1828 ( 
.A(n_1824),
.B(n_1784),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1813),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1794),
.B(n_1759),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1790),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1790),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1805),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1794),
.B(n_1787),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1811),
.B(n_1795),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1795),
.B(n_1766),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1796),
.B(n_1725),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1805),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1816),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1816),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1792),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1788),
.B(n_1733),
.Y(n_1842)
);

NAND2xp67_ASAP7_75t_L g1843 ( 
.A(n_1803),
.B(n_1694),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1796),
.B(n_1725),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1799),
.B(n_1725),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1799),
.B(n_1779),
.Y(n_1846)
);

BUFx2_ASAP7_75t_SL g1847 ( 
.A(n_1824),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1792),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1806),
.B(n_1768),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1824),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1793),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1818),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1793),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1818),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1820),
.B(n_1772),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1793),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1791),
.B(n_1823),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1819),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1803),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1826),
.B(n_1770),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1826),
.B(n_1770),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1819),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1798),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1789),
.Y(n_1864)
);

INVx2_ASAP7_75t_SL g1865 ( 
.A(n_1824),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1841),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1841),
.Y(n_1867)
);

OAI32xp33_ASAP7_75t_L g1868 ( 
.A1(n_1842),
.A2(n_1801),
.A3(n_1797),
.B1(n_1807),
.B2(n_1822),
.Y(n_1868)
);

INVxp33_ASAP7_75t_L g1869 ( 
.A(n_1842),
.Y(n_1869)
);

INVxp67_ASAP7_75t_L g1870 ( 
.A(n_1831),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1849),
.B(n_1815),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1849),
.B(n_1815),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1850),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1833),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1849),
.B(n_1815),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1849),
.B(n_1834),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1834),
.B(n_1815),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1835),
.B(n_1820),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1834),
.B(n_1812),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1841),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1833),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1831),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1833),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1835),
.B(n_1831),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1838),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1838),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1828),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1838),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1836),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1841),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1852),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_L g1892 ( 
.A(n_1864),
.B(n_1801),
.C(n_1807),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1832),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1852),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1834),
.B(n_1812),
.Y(n_1895)
);

AOI22x1_ASAP7_75t_L g1896 ( 
.A1(n_1847),
.A2(n_1822),
.B1(n_1824),
.B2(n_1800),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1848),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1852),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1846),
.B(n_1812),
.Y(n_1899)
);

OAI21xp33_ASAP7_75t_L g1900 ( 
.A1(n_1843),
.A2(n_1808),
.B(n_1810),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1854),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1832),
.B(n_1804),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1864),
.B(n_1809),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1848),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1859),
.B(n_1823),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1832),
.B(n_1804),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1855),
.B(n_1825),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1836),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1854),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1859),
.B(n_1802),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1848),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1876),
.B(n_1850),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1876),
.B(n_1877),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_SL g1914 ( 
.A1(n_1868),
.A2(n_1896),
.B1(n_1892),
.B2(n_1910),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1877),
.B(n_1850),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1879),
.B(n_1847),
.Y(n_1916)
);

NOR2x1_ASAP7_75t_L g1917 ( 
.A(n_1892),
.B(n_1910),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1874),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1874),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1870),
.B(n_1859),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1881),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1884),
.B(n_1855),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1870),
.B(n_1893),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1881),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1903),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1883),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1884),
.B(n_1855),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1879),
.B(n_1847),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1883),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1893),
.B(n_1830),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1895),
.B(n_1865),
.Y(n_1931)
);

AOI221x1_ASAP7_75t_L g1932 ( 
.A1(n_1900),
.A2(n_1797),
.B1(n_1810),
.B2(n_1869),
.C(n_1903),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1895),
.B(n_1865),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1871),
.B(n_1865),
.Y(n_1934)
);

OAI21xp33_ASAP7_75t_L g1935 ( 
.A1(n_1868),
.A2(n_1814),
.B(n_1843),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1871),
.B(n_1865),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1873),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1885),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1872),
.B(n_1830),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1872),
.B(n_1830),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1875),
.B(n_1830),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1873),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1885),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1875),
.B(n_1857),
.Y(n_1944)
);

AOI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1900),
.A2(n_1821),
.B(n_1800),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1889),
.B(n_1908),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1899),
.B(n_1857),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1882),
.B(n_1860),
.Y(n_1948)
);

OAI21xp33_ASAP7_75t_L g1949 ( 
.A1(n_1914),
.A2(n_1843),
.B(n_1814),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1913),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1942),
.Y(n_1951)
);

NAND3xp33_ASAP7_75t_L g1952 ( 
.A(n_1917),
.B(n_1896),
.C(n_1878),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1925),
.B(n_1907),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1917),
.B(n_1882),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1935),
.B(n_1899),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1937),
.Y(n_1956)
);

AOI21xp33_ASAP7_75t_L g1957 ( 
.A1(n_1935),
.A2(n_1878),
.B(n_1902),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1937),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1937),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1945),
.A2(n_1887),
.B1(n_1824),
.B2(n_1828),
.Y(n_1960)
);

AOI322xp5_ASAP7_75t_L g1961 ( 
.A1(n_1923),
.A2(n_1930),
.A3(n_1946),
.B1(n_1920),
.B2(n_1932),
.C1(n_1948),
.C2(n_1941),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1923),
.B(n_1907),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1946),
.B(n_1860),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1913),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1918),
.Y(n_1965)
);

NAND4xp25_ASAP7_75t_SL g1966 ( 
.A(n_1932),
.B(n_1821),
.C(n_1928),
.D(n_1916),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_SL g1967 ( 
.A1(n_1920),
.A2(n_1828),
.B1(n_1817),
.B2(n_1887),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1948),
.B(n_1861),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1918),
.Y(n_1969)
);

AOI22xp33_ASAP7_75t_SL g1970 ( 
.A1(n_1916),
.A2(n_1887),
.B1(n_1828),
.B2(n_1655),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1930),
.A2(n_1906),
.B1(n_1902),
.B2(n_1905),
.Y(n_1971)
);

AOI211xp5_ASAP7_75t_L g1972 ( 
.A1(n_1928),
.A2(n_1887),
.B(n_1905),
.C(n_1906),
.Y(n_1972)
);

OAI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1912),
.A2(n_1828),
.B(n_1837),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1915),
.B(n_1886),
.Y(n_1974)
);

NOR2x1_ASAP7_75t_L g1975 ( 
.A(n_1919),
.B(n_1886),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1919),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1954),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1951),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1975),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1956),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1952),
.B(n_1933),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1949),
.B(n_1915),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1958),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1966),
.A2(n_1933),
.B1(n_1931),
.B2(n_1934),
.Y(n_1984)
);

OAI21xp5_ASAP7_75t_SL g1985 ( 
.A1(n_1957),
.A2(n_1912),
.B(n_1931),
.Y(n_1985)
);

AOI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1967),
.A2(n_1933),
.B1(n_1934),
.B2(n_1936),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1959),
.Y(n_1987)
);

INVxp67_ASAP7_75t_L g1988 ( 
.A(n_1955),
.Y(n_1988)
);

NOR3xp33_ASAP7_75t_SL g1989 ( 
.A(n_1957),
.B(n_1924),
.C(n_1921),
.Y(n_1989)
);

OAI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1960),
.A2(n_1927),
.B1(n_1922),
.B2(n_1943),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1965),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1950),
.A2(n_1933),
.B1(n_1944),
.B2(n_1947),
.Y(n_1992)
);

AOI21x1_ASAP7_75t_L g1993 ( 
.A1(n_1969),
.A2(n_1924),
.B(n_1921),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1976),
.Y(n_1994)
);

OAI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1961),
.A2(n_1936),
.B(n_1927),
.Y(n_1995)
);

OAI211xp5_ASAP7_75t_L g1996 ( 
.A1(n_1972),
.A2(n_1922),
.B(n_1926),
.C(n_1943),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1964),
.B(n_1939),
.Y(n_1997)
);

AOI32xp33_ASAP7_75t_L g1998 ( 
.A1(n_1968),
.A2(n_1944),
.A3(n_1947),
.B1(n_1941),
.B2(n_1940),
.Y(n_1998)
);

AOI21xp33_ASAP7_75t_L g1999 ( 
.A1(n_1982),
.A2(n_1953),
.B(n_1962),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1987),
.Y(n_2000)
);

NOR2x1_ASAP7_75t_L g2001 ( 
.A(n_1979),
.B(n_1974),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1982),
.B(n_1974),
.Y(n_2002)
);

INVx2_ASAP7_75t_SL g2003 ( 
.A(n_1997),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1977),
.B(n_1963),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1987),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1978),
.B(n_1971),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1981),
.Y(n_2007)
);

OAI21x1_ASAP7_75t_L g2008 ( 
.A1(n_1993),
.A2(n_1973),
.B(n_1971),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1980),
.B(n_1944),
.Y(n_2009)
);

AOI221xp5_ASAP7_75t_L g2010 ( 
.A1(n_1995),
.A2(n_1973),
.B1(n_1970),
.B2(n_1929),
.C(n_1938),
.Y(n_2010)
);

AOI222xp33_ASAP7_75t_L g2011 ( 
.A1(n_1988),
.A2(n_1938),
.B1(n_1926),
.B2(n_1929),
.C1(n_1939),
.C2(n_1940),
.Y(n_2011)
);

AOI222xp33_ASAP7_75t_L g2012 ( 
.A1(n_1985),
.A2(n_1990),
.B1(n_1996),
.B2(n_1989),
.C1(n_1983),
.C2(n_1994),
.Y(n_2012)
);

OAI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1986),
.A2(n_1944),
.B1(n_1947),
.B2(n_1855),
.Y(n_2013)
);

NOR2x1_ASAP7_75t_L g2014 ( 
.A(n_2000),
.B(n_1991),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_2012),
.B(n_1998),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_2007),
.B(n_1984),
.Y(n_2016)
);

NOR2xp67_ASAP7_75t_L g2017 ( 
.A(n_2005),
.B(n_1992),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_2006),
.B(n_1990),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2009),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2009),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_2001),
.Y(n_2021)
);

AOI221x1_ASAP7_75t_L g2022 ( 
.A1(n_1999),
.A2(n_2002),
.B1(n_2004),
.B2(n_2010),
.C(n_1898),
.Y(n_2022)
);

OAI211xp5_ASAP7_75t_SL g2023 ( 
.A1(n_2003),
.A2(n_1911),
.B(n_1880),
.C(n_1867),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_2011),
.B(n_2008),
.Y(n_2024)
);

AOI221xp5_ASAP7_75t_L g2025 ( 
.A1(n_2018),
.A2(n_2015),
.B1(n_2024),
.B2(n_2016),
.C(n_2013),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2019),
.B(n_1947),
.Y(n_2026)
);

O2A1O1Ixp33_ASAP7_75t_L g2027 ( 
.A1(n_2015),
.A2(n_1840),
.B(n_1839),
.C(n_1829),
.Y(n_2027)
);

OAI221xp5_ASAP7_75t_SL g2028 ( 
.A1(n_2021),
.A2(n_1911),
.B1(n_1897),
.B2(n_1904),
.C(n_1890),
.Y(n_2028)
);

O2A1O1Ixp5_ASAP7_75t_L g2029 ( 
.A1(n_2020),
.A2(n_1911),
.B(n_1866),
.C(n_1904),
.Y(n_2029)
);

INVxp67_ASAP7_75t_L g2030 ( 
.A(n_2017),
.Y(n_2030)
);

AOI211xp5_ASAP7_75t_SL g2031 ( 
.A1(n_2023),
.A2(n_1909),
.B(n_1891),
.C(n_1894),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_SL g2032 ( 
.A(n_2030),
.B(n_2026),
.Y(n_2032)
);

OAI221xp5_ASAP7_75t_SL g2033 ( 
.A1(n_2025),
.A2(n_2022),
.B1(n_2014),
.B2(n_1867),
.C(n_1904),
.Y(n_2033)
);

NOR2x1p5_ASAP7_75t_L g2034 ( 
.A(n_2027),
.B(n_1888),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_2028),
.A2(n_1880),
.B1(n_1866),
.B2(n_1867),
.C(n_1897),
.Y(n_2035)
);

OAI211xp5_ASAP7_75t_L g2036 ( 
.A1(n_2031),
.A2(n_1866),
.B(n_1880),
.C(n_1890),
.Y(n_2036)
);

AOI221xp5_ASAP7_75t_L g2037 ( 
.A1(n_2029),
.A2(n_1897),
.B1(n_1890),
.B2(n_1898),
.C(n_1888),
.Y(n_2037)
);

NOR4xp25_ASAP7_75t_L g2038 ( 
.A(n_2025),
.B(n_1909),
.C(n_1901),
.D(n_1894),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2025),
.A2(n_1901),
.B(n_1891),
.C(n_1829),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_2032),
.A2(n_2039),
.B1(n_2038),
.B2(n_2034),
.Y(n_2040)
);

NAND4xp75_ASAP7_75t_L g2041 ( 
.A(n_2033),
.B(n_1844),
.C(n_1837),
.D(n_1845),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_2036),
.A2(n_1655),
.B1(n_1839),
.B2(n_1840),
.Y(n_2042)
);

INVxp33_ASAP7_75t_L g2043 ( 
.A(n_2035),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2037),
.Y(n_2044)
);

NAND4xp75_ASAP7_75t_L g2045 ( 
.A(n_2032),
.B(n_1844),
.C(n_1845),
.D(n_1837),
.Y(n_2045)
);

OAI322xp33_ASAP7_75t_L g2046 ( 
.A1(n_2040),
.A2(n_1840),
.A3(n_1839),
.B1(n_1829),
.B2(n_1827),
.C1(n_1863),
.C2(n_1853),
.Y(n_2046)
);

NOR2x1_ASAP7_75t_L g2047 ( 
.A(n_2041),
.B(n_1827),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2044),
.B(n_1829),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_2047),
.A2(n_2043),
.B1(n_2042),
.B2(n_2045),
.Y(n_2049)
);

AO22x2_ASAP7_75t_L g2050 ( 
.A1(n_2049),
.A2(n_2048),
.B1(n_2046),
.B2(n_1840),
.Y(n_2050)
);

OAI21xp33_ASAP7_75t_SL g2051 ( 
.A1(n_2050),
.A2(n_1839),
.B(n_1827),
.Y(n_2051)
);

AOI311xp33_ASAP7_75t_L g2052 ( 
.A1(n_2050),
.A2(n_1858),
.A3(n_1862),
.B(n_1854),
.C(n_1698),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2051),
.Y(n_2053)
);

OAI22xp5_ASAP7_75t_SL g2054 ( 
.A1(n_2052),
.A2(n_1696),
.B1(n_1695),
.B2(n_1775),
.Y(n_2054)
);

NAND2x1_ASAP7_75t_SL g2055 ( 
.A(n_2053),
.B(n_1848),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_2054),
.A2(n_1845),
.B1(n_1844),
.B2(n_1837),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_SL g2057 ( 
.A1(n_2055),
.A2(n_1696),
.B1(n_1695),
.B2(n_1786),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2057),
.A2(n_2056),
.B(n_1851),
.Y(n_2058)
);

INVx4_ASAP7_75t_L g2059 ( 
.A(n_2058),
.Y(n_2059)
);

OAI221xp5_ASAP7_75t_R g2060 ( 
.A1(n_2059),
.A2(n_1827),
.B1(n_1863),
.B2(n_1856),
.C(n_1853),
.Y(n_2060)
);

AOI211xp5_ASAP7_75t_L g2061 ( 
.A1(n_2060),
.A2(n_1697),
.B(n_1851),
.C(n_1853),
.Y(n_2061)
);


endmodule