module real_jpeg_12321_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_202;
wire n_179;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_64),
.B1(n_70),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_4),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_4),
.A2(n_30),
.B1(n_64),
.B2(n_70),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_5),
.A2(n_34),
.B1(n_37),
.B2(n_41),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_5),
.A2(n_41),
.B1(n_64),
.B2(n_70),
.Y(n_154)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_7),
.A2(n_34),
.B1(n_37),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_7),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_7),
.A2(n_64),
.B1(n_70),
.B2(n_81),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_9),
.A2(n_64),
.B1(n_70),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_9),
.Y(n_114)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_12),
.A2(n_34),
.B1(n_37),
.B2(n_58),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_12),
.A2(n_58),
.B1(n_64),
.B2(n_70),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_13),
.A2(n_64),
.B1(n_70),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_13),
.A2(n_34),
.B1(n_37),
.B2(n_72),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_14),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_14),
.A2(n_46),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_14),
.B(n_59),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_14),
.B(n_28),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_14),
.A2(n_34),
.B1(n_37),
.B2(n_76),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_14),
.A2(n_37),
.B(n_85),
.C(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_14),
.B(n_42),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_14),
.B(n_67),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_14),
.B(n_98),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_14),
.A2(n_28),
.B(n_151),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_15),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_15),
.A2(n_34),
.B1(n_37),
.B2(n_49),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_15),
.A2(n_49),
.B1(n_64),
.B2(n_70),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_16),
.A2(n_64),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_16),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_16),
.A2(n_34),
.B1(n_37),
.B2(n_69),
.Y(n_88)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_129),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_128),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_104),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_22),
.B(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_77),
.C(n_94),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_23),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_60),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_43),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_25),
.B(n_43),
.C(n_60),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_39),
.B2(n_42),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_27),
.A2(n_32),
.B1(n_33),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_28),
.A2(n_29),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_28),
.B(n_53),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_28),
.A2(n_34),
.A3(n_36),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_29),
.A2(n_46),
.A3(n_54),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_31),
.A2(n_42),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_32),
.A2(n_33),
.B1(n_40),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_32),
.A2(n_33),
.B1(n_137),
.B2(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_34),
.A2(n_37),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_35),
.B(n_37),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_50),
.B1(n_56),
.B2(n_59),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_45),
.A2(n_51),
.B1(n_52),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_51),
.A2(n_52),
.B1(n_57),
.B2(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_73),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_61),
.A2(n_62),
.B1(n_73),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_67),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_63),
.A2(n_67),
.B1(n_142),
.B2(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_63),
.A2(n_67),
.B1(n_154),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_63),
.A2(n_67),
.B1(n_76),
.B2(n_194),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_63),
.A2(n_67),
.B1(n_187),
.B2(n_194),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_64),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_70),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_64),
.B(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_66),
.A2(n_90),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_70),
.A2(n_76),
.B(n_86),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_77),
.B(n_94),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_89),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_89),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_83),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_82),
.A2(n_87),
.B1(n_145),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_98),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_83),
.A2(n_97),
.B1(n_98),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_83),
.A2(n_98),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_83),
.A2(n_98),
.B1(n_173),
.B2(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_101),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_127),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_116),
.B1(n_125),
.B2(n_126),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_115),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_225),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_221),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_165),
.B(n_220),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_155),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_133),
.B(n_155),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_143),
.C(n_146),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_134),
.B(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_140),
.C(n_141),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_148),
.A2(n_149),
.B1(n_153),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_164),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_161),
.C(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_214),
.B(n_219),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_203),
.B(n_213),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_183),
.B(n_202),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_169),
.B(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_179),
.C(n_181),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_191),
.B(n_201),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_189),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_197),
.B(n_200),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_198),
.B(n_199),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_204),
.B(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);


endmodule