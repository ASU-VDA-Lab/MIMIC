module fake_jpeg_15871_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_21),
.B(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_21),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_48),
.B(n_17),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_17),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_24),
.B1(n_23),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_56),
.B1(n_59),
.B2(n_32),
.Y(n_94)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_23),
.B1(n_27),
.B2(n_18),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_23),
.B1(n_27),
.B2(n_22),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_60)
);

OA22x2_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_43),
.B1(n_41),
.B2(n_35),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_63),
.B(n_69),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_39),
.B1(n_42),
.B2(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_64),
.A2(n_88),
.B1(n_92),
.B2(n_96),
.Y(n_117)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_77),
.B(n_82),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_76),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_73),
.B(n_78),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_95),
.B(n_30),
.C(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_37),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_39),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_79),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_34),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_84),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_0),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_22),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_85),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_0),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_61),
.B1(n_49),
.B2(n_30),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_19),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_19),
.B1(n_32),
.B2(n_20),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_53),
.B1(n_51),
.B2(n_49),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_98),
.B1(n_61),
.B2(n_30),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_20),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_26),
.B1(n_30),
.B2(n_29),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_56),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_99),
.B1(n_53),
.B2(n_49),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_60),
.C(n_31),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_86),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_99),
.B1(n_66),
.B2(n_65),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_106),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_123),
.B1(n_79),
.B2(n_77),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_63),
.B1(n_96),
.B2(n_74),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_74),
.B1(n_72),
.B2(n_76),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_68),
.A2(n_25),
.B1(n_18),
.B2(n_16),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_125),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_129),
.B(n_156),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_137),
.B1(n_117),
.B2(n_106),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_140),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_82),
.B(n_86),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_133),
.A2(n_29),
.B(n_25),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_134),
.B(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_75),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_143),
.B1(n_146),
.B2(n_149),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_129),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_82),
.B1(n_75),
.B2(n_74),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_147),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_77),
.B1(n_94),
.B2(n_92),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_64),
.B1(n_65),
.B2(n_14),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_25),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_105),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_16),
.Y(n_155)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_30),
.C(n_29),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_127),
.B1(n_103),
.B2(n_125),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_179),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_113),
.B(n_126),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_113),
.B1(n_117),
.B2(n_105),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_163),
.A2(n_165),
.B1(n_174),
.B2(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_107),
.Y(n_168)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_156),
.C(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_31),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_104),
.B(n_109),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_153),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_107),
.B1(n_104),
.B2(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_18),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_180),
.B(n_0),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_136),
.A2(n_89),
.B1(n_67),
.B2(n_108),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_108),
.B1(n_89),
.B2(n_67),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_185),
.A2(n_186),
.B1(n_140),
.B2(n_31),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_133),
.A2(n_108),
.B1(n_25),
.B2(n_18),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_158),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_142),
.C(n_16),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_163),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_179),
.B(n_172),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_187),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_200),
.C(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_154),
.C(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_212),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_213),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_206),
.A2(n_209),
.B1(n_215),
.B2(n_172),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_1),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_164),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_165),
.A2(n_178),
.B1(n_185),
.B2(n_173),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_181),
.B(n_7),
.CI(n_13),
.CON(n_216),
.SN(n_216)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_218),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_15),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_170),
.B(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_223),
.B(n_1),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_161),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_225),
.C(n_227),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_197),
.C(n_217),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_174),
.B1(n_183),
.B2(n_162),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_240),
.B1(n_214),
.B2(n_196),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_159),
.C(n_167),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_230),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_186),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_166),
.B1(n_189),
.B2(n_175),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_223),
.Y(n_243)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_203),
.A2(n_207),
.B1(n_193),
.B2(n_210),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_192),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_237),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_176),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_169),
.C(n_184),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_214),
.C(n_204),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_207),
.A2(n_184),
.B1(n_190),
.B2(n_3),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_244),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_216),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_259),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_228),
.A2(n_201),
.B(n_204),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_254),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_229),
.B(n_216),
.CI(n_196),
.CON(n_247),
.SN(n_247)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_247),
.B(n_251),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_255),
.C(n_260),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_239),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_194),
.C(n_211),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_194),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_221),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_238),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_2),
.C(n_5),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_6),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_6),
.C(n_8),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_245),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_232),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_274),
.C(n_276),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_236),
.B(n_235),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_271),
.B(n_256),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_SL g270 ( 
.A1(n_247),
.A2(n_220),
.A3(n_226),
.B1(n_240),
.B2(n_230),
.C1(n_10),
.C2(n_11),
.Y(n_270)
);

OAI221xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.C(n_5),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_6),
.Y(n_273)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_2),
.C(n_5),
.Y(n_276)
);

BUFx12f_ASAP7_75t_SL g277 ( 
.A(n_252),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_250),
.B1(n_252),
.B2(n_243),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_288),
.C(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_259),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_268),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_299),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_281),
.A2(n_275),
.B(n_268),
.C(n_266),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_300),
.B(n_289),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_262),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_261),
.C(n_260),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_281),
.B(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_305),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_279),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_300),
.C(n_297),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_308),
.A2(n_301),
.B(n_293),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_292),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_310),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_309),
.Y(n_314)
);

OAI311xp33_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_313),
.A3(n_311),
.B1(n_307),
.C1(n_291),
.Y(n_315)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_8),
.B(n_10),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_5),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_317),
.Y(n_318)
);


endmodule