module fake_ariane_426_n_1845 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1845);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1845;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1660;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_129),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_65),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_6),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_86),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_170),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_66),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_26),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_136),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_184),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_104),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_53),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_84),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_96),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_148),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_56),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_50),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_69),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_142),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_110),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_42),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_109),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_89),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_87),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_73),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_20),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_103),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_165),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_176),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_53),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_75),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_34),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_83),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_92),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_91),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_128),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_143),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_138),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_68),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_108),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_150),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_29),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_130),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_161),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_137),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_71),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_112),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_181),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_121),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_134),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_125),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_95),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_169),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_133),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_33),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_17),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_80),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_21),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_78),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_93),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_106),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_45),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_100),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_107),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_172),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_28),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_182),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_61),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_3),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_119),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_29),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_22),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_2),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_19),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_22),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_126),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_21),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_23),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_27),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_57),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_62),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_162),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_19),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_120),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_127),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_7),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_64),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_32),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_15),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_74),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_41),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_147),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_55),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_159),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_3),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_4),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_61),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_114),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_16),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_101),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_77),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_26),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_118),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_81),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_90),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_15),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_70),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_145),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_117),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_178),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_183),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_5),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_160),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_173),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_115),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_179),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_64),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_14),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_46),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_111),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_37),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_9),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_174),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_65),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_132),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_46),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_10),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_13),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_32),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_116),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_76),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_39),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_50),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_58),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_188),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_124),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_139),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_16),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_149),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_102),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_98),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_57),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_47),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_56),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_18),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_141),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_8),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_30),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_52),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_25),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_164),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_14),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_155),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_85),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_13),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_47),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_4),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_25),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_49),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_62),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_36),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_167),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_99),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_187),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_140),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_52),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_88),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_42),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_18),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_144),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_63),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_39),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_36),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_6),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_49),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_292),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_280),
.B(n_0),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_267),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_278),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_292),
.B(n_0),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_253),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_295),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_377),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_293),
.B(n_1),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_201),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_205),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_295),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_213),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_295),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_215),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_294),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_295),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_203),
.B(n_1),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_296),
.Y(n_398)
);

INVxp33_ASAP7_75t_SL g399 ( 
.A(n_330),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_295),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_217),
.B(n_5),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_334),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_317),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_195),
.Y(n_405)
);

INVxp33_ASAP7_75t_SL g406 ( 
.A(n_353),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_318),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_371),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_210),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_300),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_257),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_259),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_263),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_222),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_326),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_227),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_326),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_351),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_271),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_274),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_230),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_231),
.B(n_233),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_212),
.B(n_8),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_275),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_360),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_195),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_249),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_281),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_360),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_270),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_282),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_284),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_289),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_303),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_306),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_360),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_219),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_310),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_316),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_273),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_321),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_363),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_354),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_238),
.B(n_9),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_373),
.B(n_10),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_373),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_249),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_194),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_306),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_291),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_301),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_208),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_234),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_234),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_288),
.B(n_11),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_252),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_192),
.B(n_206),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_209),
.B(n_11),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_252),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_194),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_198),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_198),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_354),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_327),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_390),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_410),
.B(n_211),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_457),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_405),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_409),
.Y(n_481)
);

CKINVDCx8_ASAP7_75t_R g482 ( 
.A(n_394),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_416),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_458),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_404),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_407),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_408),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_403),
.B(n_354),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_399),
.A2(n_376),
.B1(n_338),
.B2(n_193),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_434),
.B(n_229),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_382),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_402),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_418),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_381),
.B(n_219),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_385),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_411),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_427),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_389),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_385),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_392),
.Y(n_507)
);

NAND2xp33_ASAP7_75t_L g508 ( 
.A(n_381),
.B(n_190),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_438),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_434),
.B(n_232),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_403),
.B(n_249),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_435),
.B(n_314),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_421),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_411),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_385),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_395),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_449),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_415),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_385),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_417),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_385),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_383),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_398),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_461),
.B(n_314),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_428),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_413),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_459),
.Y(n_529)
);

NOR2x1_ASAP7_75t_L g530 ( 
.A(n_462),
.B(n_228),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_414),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_424),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_417),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_421),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_419),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_420),
.Y(n_537)
);

AND2x2_ASAP7_75t_SL g538 ( 
.A(n_435),
.B(n_327),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_426),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_456),
.B(n_314),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_430),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_420),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_422),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_456),
.B(n_340),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_422),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_460),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_445),
.B(n_236),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_538),
.B(n_436),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_544),
.Y(n_551)
);

NAND3xp33_ASAP7_75t_L g552 ( 
.A(n_508),
.B(n_440),
.C(n_439),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_538),
.B(n_441),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_538),
.B(n_442),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_501),
.B(n_466),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_544),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_501),
.B(n_446),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_524),
.B(n_452),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_544),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_480),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_543),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_474),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_524),
.B(n_470),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_480),
.B(n_448),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_515),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_474),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_479),
.A2(n_401),
.B1(n_406),
.B2(n_397),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_501),
.A2(n_464),
.B1(n_453),
.B2(n_429),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_543),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_536),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_543),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_476),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_476),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_540),
.B(n_401),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_482),
.B(n_387),
.Y(n_575)
);

BUFx4f_ASAP7_75t_L g576 ( 
.A(n_540),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_545),
.B(n_511),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_502),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_519),
.B(n_532),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_536),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_501),
.A2(n_467),
.B1(n_388),
.B2(n_454),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_481),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_494),
.B(n_471),
.Y(n_583)
);

INVx8_ASAP7_75t_L g584 ( 
.A(n_527),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_519),
.B(n_450),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_519),
.B(n_237),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_526),
.A2(n_472),
.B1(n_269),
.B2(n_362),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_484),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_519),
.B(n_532),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_484),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_545),
.B(n_447),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_485),
.B(n_384),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_532),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_497),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_511),
.B(n_447),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_485),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_483),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_548),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_502),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_543),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_543),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_526),
.B(n_380),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_491),
.B(n_451),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_478),
.B(n_380),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_494),
.B(n_528),
.Y(n_605)
);

NOR2x1p5_ASAP7_75t_L g606 ( 
.A(n_531),
.B(n_202),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_532),
.B(n_239),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_495),
.B(n_462),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_510),
.B(n_530),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_537),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_512),
.A2(n_283),
.B1(n_347),
.B2(n_336),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_489),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_549),
.B(n_455),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_539),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_541),
.B(n_455),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_477),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_489),
.B(n_344),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_490),
.B(n_463),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_490),
.A2(n_299),
.B1(n_297),
.B2(n_290),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_486),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_492),
.B(n_465),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_492),
.B(n_465),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_496),
.B(n_468),
.Y(n_624)
);

INVx4_ASAP7_75t_SL g625 ( 
.A(n_537),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_502),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_487),
.B(n_202),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_488),
.B(n_473),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_482),
.B(n_473),
.Y(n_629)
);

AND2x2_ASAP7_75t_SL g630 ( 
.A(n_498),
.B(n_344),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_498),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_493),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_515),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_505),
.B(n_507),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_537),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_499),
.A2(n_256),
.B1(n_379),
.B2(n_333),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_493),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_499),
.B(n_423),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_503),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_516),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_537),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_537),
.B(n_245),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_503),
.B(n_251),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_514),
.B(n_240),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_514),
.B(n_276),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_513),
.Y(n_646)
);

BUFx4f_ASAP7_75t_L g647 ( 
.A(n_518),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_502),
.Y(n_648)
);

INVxp33_ASAP7_75t_SL g649 ( 
.A(n_525),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_518),
.B(n_423),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_521),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_513),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_534),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_521),
.B(n_228),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_522),
.B(n_247),
.Y(n_655)
);

OAI21xp33_ASAP7_75t_SL g656 ( 
.A1(n_522),
.A2(n_286),
.B(n_277),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_533),
.A2(n_361),
.B1(n_375),
.B2(n_331),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_535),
.B(n_241),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_535),
.B(n_425),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_506),
.Y(n_660)
);

INVx6_ASAP7_75t_L g661 ( 
.A(n_506),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_506),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_542),
.A2(n_340),
.B1(n_258),
.B2(n_248),
.Y(n_663)
);

INVx5_ASAP7_75t_L g664 ( 
.A(n_515),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_542),
.B(n_546),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_546),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_534),
.B(n_241),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_500),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_523),
.B(n_262),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_523),
.A2(n_340),
.B1(n_214),
.B2(n_312),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_523),
.B(n_262),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_515),
.B(n_250),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_523),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_504),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_509),
.Y(n_675)
);

INVxp33_ASAP7_75t_L g676 ( 
.A(n_517),
.Y(n_676)
);

INVxp33_ASAP7_75t_L g677 ( 
.A(n_529),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_547),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_515),
.B(n_255),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_520),
.B(n_224),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_520),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_520),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_520),
.B(n_260),
.Y(n_683)
);

INVx5_ASAP7_75t_L g684 ( 
.A(n_515),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_475),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_665),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_630),
.B(n_265),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_598),
.B(n_218),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_L g689 ( 
.A(n_593),
.B(n_431),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_596),
.B(n_190),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_630),
.B(n_191),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_604),
.B(n_191),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_675),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_613),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_613),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_550),
.B(n_224),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_562),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_576),
.B(n_197),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_558),
.B(n_605),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_550),
.A2(n_196),
.B1(n_315),
.B2(n_207),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_553),
.A2(n_315),
.B1(n_207),
.B2(n_235),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_555),
.A2(n_342),
.B(n_332),
.C(n_328),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_592),
.B(n_199),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_553),
.B(n_554),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_567),
.B(n_342),
.C(n_332),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_592),
.B(n_199),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_566),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_572),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_582),
.B(n_322),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_554),
.B(n_322),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_592),
.B(n_200),
.Y(n_711)
);

NAND2x1_ASAP7_75t_L g712 ( 
.A(n_661),
.B(n_431),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_608),
.B(n_200),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_577),
.B(n_323),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_576),
.B(n_204),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_617),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_608),
.B(n_204),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_557),
.B(n_323),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_602),
.B(n_591),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_595),
.B(n_216),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_609),
.B(n_216),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_616),
.B(n_325),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_563),
.B(n_325),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_614),
.Y(n_724)
);

INVxp33_ASAP7_75t_L g725 ( 
.A(n_634),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_586),
.B(n_328),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_632),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_609),
.B(n_220),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_632),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_647),
.B(n_221),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_668),
.B(n_337),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_564),
.B(n_603),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_594),
.B(n_585),
.C(n_621),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_573),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_647),
.A2(n_590),
.B(n_588),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_656),
.A2(n_444),
.B(n_437),
.C(n_433),
.Y(n_736)
);

NOR3x1_ASAP7_75t_L g737 ( 
.A(n_627),
.B(n_378),
.C(n_372),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_564),
.B(n_221),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_568),
.A2(n_337),
.B1(n_346),
.B2(n_348),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_637),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_629),
.B(n_223),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_586),
.B(n_225),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_628),
.B(n_226),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_637),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_643),
.B(n_226),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_643),
.B(n_607),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_646),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_607),
.B(n_346),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_612),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_560),
.B(n_324),
.Y(n_751)
);

AND2x2_ASAP7_75t_SL g752 ( 
.A(n_583),
.B(n_266),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_597),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_644),
.B(n_324),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_644),
.B(n_329),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_631),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_569),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_615),
.B(n_348),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_584),
.B(n_235),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_644),
.B(n_329),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_621),
.B(n_364),
.C(n_349),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_644),
.B(n_645),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_614),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_639),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_646),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_651),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_645),
.B(n_335),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_552),
.B(n_349),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_652),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_569),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_652),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_585),
.B(n_352),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_615),
.B(n_352),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_653),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_574),
.A2(n_350),
.B1(n_358),
.B2(n_374),
.Y(n_775)
);

BUFx4f_ASAP7_75t_SL g776 ( 
.A(n_597),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_666),
.Y(n_777)
);

OAI221xp5_ASAP7_75t_L g778 ( 
.A1(n_581),
.A2(n_362),
.B1(n_356),
.B2(n_359),
.C(n_364),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_574),
.A2(n_350),
.B1(n_358),
.B2(n_374),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_618),
.A2(n_356),
.B1(n_359),
.B2(n_365),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_614),
.B(n_365),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_614),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_579),
.B(n_370),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_574),
.A2(n_335),
.B1(n_304),
.B2(n_308),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_574),
.A2(n_268),
.B1(n_339),
.B2(n_341),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_645),
.B(n_370),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_579),
.B(n_372),
.Y(n_787)
);

AO221x1_ASAP7_75t_L g788 ( 
.A1(n_561),
.A2(n_367),
.B1(n_357),
.B2(n_253),
.C(n_366),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_619),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_623),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_624),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_589),
.B(n_378),
.Y(n_792)
);

O2A1O1Ixp5_ASAP7_75t_L g793 ( 
.A1(n_635),
.A2(n_369),
.B(n_345),
.C(n_355),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_638),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_L g795 ( 
.A1(n_618),
.A2(n_368),
.B1(n_343),
.B2(n_433),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_570),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_645),
.B(n_242),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_570),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_650),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_658),
.B(n_243),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_658),
.B(n_551),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_674),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_587),
.B(n_589),
.C(n_685),
.Y(n_803)
);

OAI221xp5_ASAP7_75t_L g804 ( 
.A1(n_620),
.A2(n_444),
.B1(n_437),
.B2(n_432),
.C(n_305),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_580),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_611),
.A2(n_302),
.B1(n_246),
.B2(n_261),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_560),
.A2(n_307),
.B1(n_264),
.B2(n_272),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_560),
.Y(n_808)
);

INVx8_ASAP7_75t_L g809 ( 
.A(n_584),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_580),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_556),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_606),
.B(n_432),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_658),
.B(n_244),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_584),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_635),
.A2(n_641),
.B(n_571),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_659),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_640),
.B(n_12),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_618),
.A2(n_253),
.B1(n_357),
.B2(n_367),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_680),
.A2(n_309),
.B1(n_285),
.B2(n_320),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_559),
.B(n_12),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_680),
.A2(n_298),
.B1(n_319),
.B2(n_313),
.Y(n_821)
);

O2A1O1Ixp5_ASAP7_75t_L g822 ( 
.A1(n_635),
.A2(n_279),
.B(n_287),
.C(n_311),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_575),
.B(n_17),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_561),
.B(n_23),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_655),
.B(n_622),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_654),
.A2(n_254),
.B1(n_357),
.B2(n_253),
.Y(n_826)
);

BUFx4_ASAP7_75t_L g827 ( 
.A(n_649),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_584),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_676),
.B(n_24),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_655),
.B(n_254),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_622),
.B(n_254),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_667),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_663),
.A2(n_367),
.B1(n_253),
.B2(n_28),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_571),
.B(n_27),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_667),
.Y(n_835)
);

OR2x6_ASAP7_75t_SL g836 ( 
.A(n_739),
.B(n_649),
.Y(n_836)
);

OA22x2_ASAP7_75t_L g837 ( 
.A1(n_781),
.A2(n_642),
.B1(n_676),
.B2(n_677),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_809),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_699),
.B(n_725),
.Y(n_839)
);

NOR3xp33_ASAP7_75t_L g840 ( 
.A(n_772),
.B(n_600),
.C(n_642),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_687),
.A2(n_657),
.B1(n_636),
.B2(n_670),
.Y(n_841)
);

NOR2x1_ASAP7_75t_L g842 ( 
.A(n_828),
.B(n_578),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_686),
.B(n_654),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_697),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_802),
.B(n_677),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_707),
.Y(n_846)
);

INVx5_ASAP7_75t_L g847 ( 
.A(n_809),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_747),
.B(n_618),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_776),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_753),
.B(n_667),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_809),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_719),
.B(n_618),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_789),
.B(n_669),
.Y(n_853)
);

BUFx8_ASAP7_75t_L g854 ( 
.A(n_781),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_790),
.B(n_669),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_687),
.A2(n_713),
.B1(n_717),
.B2(n_746),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_776),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_763),
.B(n_569),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_791),
.B(n_669),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_688),
.B(n_671),
.Y(n_860)
);

AO21x1_ASAP7_75t_L g861 ( 
.A1(n_704),
.A2(n_830),
.B(n_738),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_752),
.B(n_662),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_828),
.Y(n_863)
);

AO21x1_ASAP7_75t_L g864 ( 
.A1(n_704),
.A2(n_683),
.B(n_679),
.Y(n_864)
);

OR2x6_ASAP7_75t_SL g865 ( 
.A(n_827),
.B(n_30),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_793),
.A2(n_683),
.B(n_679),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_718),
.B(n_794),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_723),
.B(n_671),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_782),
.B(n_601),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_831),
.A2(n_672),
.B(n_578),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_799),
.B(n_601),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_752),
.A2(n_601),
.B1(n_569),
.B2(n_672),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_696),
.A2(n_682),
.B(n_681),
.C(n_610),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_751),
.A2(n_648),
.B(n_626),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_691),
.A2(n_601),
.B1(n_610),
.B2(n_648),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_751),
.A2(n_660),
.B(n_626),
.Y(n_876)
);

OAI21xp33_ASAP7_75t_L g877 ( 
.A1(n_772),
.A2(n_749),
.B(n_726),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_762),
.B(n_610),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_816),
.B(n_741),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_730),
.A2(n_578),
.B(n_662),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_691),
.A2(n_610),
.B1(n_599),
.B2(n_673),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_696),
.A2(n_682),
.B(n_681),
.C(n_565),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_694),
.Y(n_883)
);

NOR2xp67_ASAP7_75t_L g884 ( 
.A(n_814),
.B(n_662),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_757),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_757),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_812),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_710),
.A2(n_749),
.B1(n_726),
.B2(n_833),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_690),
.B(n_722),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_708),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_734),
.B(n_625),
.Y(n_891)
);

BUFx4f_ASAP7_75t_L g892 ( 
.A(n_759),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_724),
.B(n_625),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_808),
.A2(n_715),
.B(n_698),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_724),
.B(n_684),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_824),
.A2(n_684),
.B(n_664),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_714),
.B(n_661),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_824),
.A2(n_664),
.B(n_633),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_757),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_693),
.Y(n_900)
);

AOI21xp33_ASAP7_75t_L g901 ( 
.A1(n_768),
.A2(n_31),
.B(n_33),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_745),
.B(n_803),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_705),
.A2(n_633),
.B1(n_565),
.B2(n_35),
.Y(n_903)
);

BUFx4f_ASAP7_75t_L g904 ( 
.A(n_759),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_750),
.A2(n_565),
.B(n_72),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_778),
.A2(n_31),
.B(n_34),
.C(n_35),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_694),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_756),
.A2(n_565),
.B(n_82),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_716),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_783),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_834),
.A2(n_38),
.B(n_40),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_764),
.A2(n_97),
.B(n_185),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_783),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_766),
.A2(n_94),
.B(n_171),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_757),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_777),
.A2(n_79),
.B(n_168),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_L g917 ( 
.A(n_733),
.B(n_43),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_702),
.A2(n_44),
.B(n_48),
.C(n_51),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_787),
.B(n_792),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_787),
.B(n_48),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_792),
.A2(n_51),
.B(n_54),
.C(n_55),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_801),
.A2(n_123),
.B(n_163),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_796),
.A2(n_113),
.B(n_158),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_798),
.A2(n_805),
.B(n_813),
.Y(n_924)
);

BUFx4f_ASAP7_75t_L g925 ( 
.A(n_759),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_758),
.Y(n_926)
);

AOI22x1_ASAP7_75t_L g927 ( 
.A1(n_811),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_770),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_780),
.B(n_59),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_834),
.A2(n_60),
.B(n_63),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_800),
.A2(n_135),
.B(n_67),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_770),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_716),
.A2(n_105),
.B(n_131),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_770),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_692),
.B(n_60),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_702),
.A2(n_146),
.B(n_152),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_820),
.A2(n_736),
.B(n_822),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_832),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_743),
.B(n_720),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_768),
.B(n_773),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_770),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_775),
.B(n_779),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_721),
.B(n_728),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_780),
.B(n_797),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_754),
.B(n_755),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_740),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_L g947 ( 
.A(n_761),
.B(n_742),
.C(n_786),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_760),
.B(n_767),
.Y(n_948)
);

OAI321xp33_ASAP7_75t_L g949 ( 
.A1(n_785),
.A2(n_784),
.A3(n_701),
.B1(n_700),
.B2(n_823),
.C(n_818),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_744),
.A2(n_774),
.B(n_765),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_744),
.A2(n_769),
.B(n_748),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_771),
.A2(n_774),
.B(n_810),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_712),
.Y(n_953)
);

NAND2x1_ASAP7_75t_L g954 ( 
.A(n_771),
.B(n_695),
.Y(n_954)
);

CKINVDCx10_ASAP7_75t_R g955 ( 
.A(n_737),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_742),
.A2(n_703),
.B(n_706),
.C(n_711),
.Y(n_956)
);

AOI21xp33_ASAP7_75t_L g957 ( 
.A1(n_709),
.A2(n_731),
.B(n_835),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_820),
.B(n_689),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_727),
.Y(n_959)
);

AO32x1_ASAP7_75t_L g960 ( 
.A1(n_729),
.A2(n_788),
.A3(n_817),
.B1(n_807),
.B2(n_806),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_812),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_819),
.B(n_821),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_818),
.A2(n_826),
.B(n_795),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_829),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_804),
.Y(n_965)
);

OR2x6_ASAP7_75t_SL g966 ( 
.A(n_795),
.B(n_621),
.Y(n_966)
);

CKINVDCx16_ASAP7_75t_R g967 ( 
.A(n_753),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_723),
.B(n_577),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_825),
.A2(n_815),
.B(n_735),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_694),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_793),
.A2(n_735),
.B(n_747),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_732),
.A2(n_825),
.B(n_739),
.C(n_747),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_825),
.A2(n_815),
.B(n_735),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_732),
.A2(n_825),
.B(n_739),
.C(n_747),
.Y(n_974)
);

NOR2x1_ASAP7_75t_L g975 ( 
.A(n_828),
.B(n_615),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_825),
.A2(n_815),
.B(n_735),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_697),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_732),
.B(n_576),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_732),
.B(n_596),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_694),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_757),
.Y(n_981)
);

O2A1O1Ixp5_ASAP7_75t_L g982 ( 
.A1(n_738),
.A2(n_825),
.B(n_751),
.C(n_730),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_732),
.B(n_596),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_825),
.A2(n_732),
.B1(n_687),
.B2(n_747),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_732),
.A2(n_825),
.B(n_739),
.C(n_747),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_687),
.A2(n_752),
.B1(n_577),
.B2(n_691),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_825),
.A2(n_815),
.B(n_735),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_825),
.A2(n_815),
.B(n_735),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_825),
.A2(n_815),
.B(n_735),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_776),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_825),
.A2(n_732),
.B1(n_687),
.B2(n_747),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_793),
.A2(n_735),
.B(n_747),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_732),
.A2(n_825),
.B(n_739),
.C(n_747),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_732),
.B(n_596),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_699),
.B(n_390),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_809),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_825),
.A2(n_732),
.B1(n_687),
.B2(n_747),
.Y(n_997)
);

NAND2x1_ASAP7_75t_L g998 ( 
.A(n_996),
.B(n_885),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_838),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_940),
.B(n_877),
.Y(n_1000)
);

AOI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_919),
.A2(n_888),
.B(n_856),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_849),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_967),
.B(n_995),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_900),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_839),
.B(n_968),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_987),
.A2(n_989),
.B(n_988),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_984),
.B(n_991),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_838),
.Y(n_1009)
);

O2A1O1Ixp5_ASAP7_75t_L g1010 ( 
.A1(n_920),
.A2(n_937),
.B(n_958),
.C(n_864),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_997),
.B(n_979),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_857),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_896),
.A2(n_898),
.B(n_867),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_844),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_942),
.A2(n_972),
.B(n_985),
.C(n_993),
.Y(n_1015)
);

BUFx12f_ASAP7_75t_L g1016 ( 
.A(n_990),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_971),
.A2(n_992),
.B(n_974),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_846),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_890),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_887),
.B(n_961),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_983),
.A2(n_994),
.B1(n_986),
.B2(n_962),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_911),
.A2(n_930),
.B(n_913),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_982),
.A2(n_956),
.B(n_943),
.C(n_879),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_939),
.B(n_862),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_950),
.A2(n_951),
.B(n_952),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_889),
.B(n_977),
.Y(n_1026)
);

AO31x2_ASAP7_75t_L g1027 ( 
.A1(n_861),
.A2(n_873),
.A3(n_882),
.B(n_924),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_838),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_896),
.A2(n_898),
.B(n_894),
.Y(n_1029)
);

BUFx4_ASAP7_75t_SL g1030 ( 
.A(n_863),
.Y(n_1030)
);

CKINVDCx16_ASAP7_75t_R g1031 ( 
.A(n_836),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_851),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_938),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_936),
.A2(n_945),
.B(n_948),
.C(n_902),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_961),
.B(n_926),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_911),
.A2(n_930),
.B(n_906),
.C(n_949),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_847),
.B(n_892),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_966),
.A2(n_935),
.B1(n_963),
.B2(n_903),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_949),
.A2(n_944),
.B(n_901),
.C(n_848),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_978),
.B(n_946),
.Y(n_1040)
);

NAND2x1p5_ASAP7_75t_L g1041 ( 
.A(n_847),
.B(n_996),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_847),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_917),
.A2(n_921),
.B(n_910),
.C(n_929),
.Y(n_1043)
);

NAND2x1_ASAP7_75t_L g1044 ( 
.A(n_885),
.B(n_886),
.Y(n_1044)
);

AO21x1_ASAP7_75t_L g1045 ( 
.A1(n_937),
.A2(n_866),
.B(n_843),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_866),
.A2(n_852),
.B(n_870),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_850),
.B(n_845),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_SL g1048 ( 
.A1(n_871),
.A2(n_931),
.B(n_918),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_959),
.Y(n_1049)
);

AO21x2_ASAP7_75t_L g1050 ( 
.A1(n_870),
.A2(n_875),
.B(n_840),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_874),
.A2(n_876),
.B(n_880),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_905),
.A2(n_908),
.B(n_954),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_975),
.B(n_851),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_922),
.A2(n_923),
.B(n_933),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_868),
.B(n_841),
.Y(n_1055)
);

AO31x2_ASAP7_75t_L g1056 ( 
.A1(n_907),
.A2(n_909),
.A3(n_980),
.B(n_970),
.Y(n_1056)
);

AND3x4_ASAP7_75t_L g1057 ( 
.A(n_947),
.B(n_955),
.C(n_865),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_L g1058 ( 
.A(n_927),
.B(n_841),
.C(n_897),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_965),
.B(n_860),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_853),
.A2(n_859),
.B(n_855),
.C(n_957),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_892),
.B(n_904),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_851),
.B(n_893),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_964),
.B(n_904),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_872),
.B(n_895),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_878),
.A2(n_914),
.B(n_916),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_891),
.A2(n_981),
.B(n_941),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_912),
.A2(n_981),
.B(n_886),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_960),
.A2(n_837),
.A3(n_881),
.B(n_858),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_925),
.B(n_837),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_941),
.B(n_934),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_899),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_869),
.A2(n_884),
.B(n_842),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_899),
.A2(n_932),
.B(n_915),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_925),
.A2(n_960),
.B(n_899),
.C(n_915),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_915),
.A2(n_928),
.B(n_932),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_928),
.A2(n_932),
.B(n_934),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_928),
.A2(n_934),
.B(n_960),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_953),
.A2(n_864),
.A3(n_861),
.B(n_873),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_854),
.A2(n_973),
.B(n_969),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_854),
.A2(n_973),
.B(n_969),
.Y(n_1080)
);

NOR2x1_ASAP7_75t_L g1081 ( 
.A(n_863),
.B(n_615),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_919),
.A2(n_984),
.B1(n_997),
.B2(n_991),
.Y(n_1082)
);

OA21x2_ASAP7_75t_L g1083 ( 
.A1(n_864),
.A2(n_973),
.B(n_969),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_979),
.B(n_983),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_883),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_L g1089 ( 
.A1(n_919),
.A2(n_920),
.B(n_856),
.C(n_738),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_883),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_847),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_900),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_849),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_847),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_877),
.A2(n_919),
.B(n_940),
.C(n_888),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_984),
.B(n_991),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_847),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_SL g1101 ( 
.A1(n_984),
.A2(n_997),
.B(n_991),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_961),
.B(n_828),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_877),
.A2(n_919),
.B(n_888),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_984),
.B(n_991),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_847),
.Y(n_1105)
);

NOR2xp67_ASAP7_75t_SL g1106 ( 
.A(n_847),
.B(n_615),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_838),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1110)
);

AOI21xp33_ASAP7_75t_L g1111 ( 
.A1(n_877),
.A2(n_919),
.B(n_888),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1112)
);

OAI222xp33_ASAP7_75t_L g1113 ( 
.A1(n_841),
.A2(n_494),
.B1(n_605),
.B2(n_583),
.C1(n_986),
.C2(n_427),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_847),
.B(n_996),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_984),
.B(n_991),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_877),
.B(n_649),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_877),
.A2(n_919),
.B(n_940),
.C(n_888),
.Y(n_1120)
);

AND2x2_ASAP7_75t_SL g1121 ( 
.A(n_942),
.B(n_687),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_942),
.A2(n_877),
.B1(n_621),
.B2(n_940),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_838),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_984),
.B(n_991),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_984),
.B(n_991),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_877),
.A2(n_919),
.B(n_940),
.C(n_888),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_984),
.B(n_991),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_849),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_883),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_877),
.A2(n_919),
.B(n_940),
.C(n_888),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_864),
.A2(n_861),
.A3(n_873),
.B(n_882),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_844),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_984),
.B(n_991),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_896),
.A2(n_898),
.B(n_825),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_969),
.A2(n_976),
.B(n_973),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1024),
.B(n_1122),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1094),
.A2(n_1117),
.B(n_1095),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_SL g1145 ( 
.A(n_1071),
.B(n_1042),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1078),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1121),
.B(n_1006),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1014),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1047),
.B(n_1093),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1061),
.B(n_1037),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1024),
.B(n_1026),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1042),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_1031),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1071),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1113),
.B(n_1118),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1018),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1085),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_L g1158 ( 
.A(n_1001),
.B(n_1022),
.C(n_1082),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1008),
.A2(n_1125),
.B1(n_1116),
.B2(n_1104),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1098),
.B(n_1127),
.C(n_1120),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1100),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1112),
.A2(n_1123),
.B(n_1115),
.Y(n_1162)
);

CKINVDCx6p67_ASAP7_75t_R g1163 ( 
.A(n_1016),
.Y(n_1163)
);

AND2x2_ASAP7_75t_SL g1164 ( 
.A(n_1008),
.B(n_1099),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_SL g1165 ( 
.A(n_1003),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1056),
.Y(n_1166)
);

BUFx8_ASAP7_75t_L g1167 ( 
.A(n_1129),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1102),
.B(n_1020),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1071),
.B(n_1009),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1026),
.B(n_1086),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1132),
.B(n_1001),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1102),
.B(n_1020),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1078),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1004),
.B(n_1106),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1000),
.B(n_1005),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1059),
.B(n_1035),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1020),
.B(n_1009),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1009),
.B(n_1053),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1011),
.A2(n_1021),
.B(n_1034),
.Y(n_1179)
);

OAI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1015),
.A2(n_1104),
.B(n_1128),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1069),
.B(n_1019),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1021),
.B(n_1011),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1103),
.A2(n_1111),
.B1(n_1038),
.B2(n_1055),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_999),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1137),
.B(n_1033),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1063),
.B(n_1103),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1078),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1133),
.Y(n_1188)
);

NAND2x1_ASAP7_75t_L g1189 ( 
.A(n_1100),
.B(n_1105),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1053),
.B(n_999),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1111),
.B(n_1099),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1134),
.A2(n_1139),
.B(n_1135),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1081),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1036),
.A2(n_1138),
.B(n_1116),
.C(n_1125),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1082),
.B(n_1126),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1087),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1101),
.B(n_1126),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1090),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1030),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1049),
.B(n_1096),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_999),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1013),
.A2(n_1128),
.B(n_1138),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1023),
.B(n_1012),
.Y(n_1203)
);

AOI21xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1057),
.A2(n_1038),
.B(n_1043),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1094),
.A2(n_1142),
.B(n_1119),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1079),
.B(n_1089),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1095),
.A2(n_1117),
.B(n_1131),
.Y(n_1207)
);

NOR2x1_ASAP7_75t_SL g1208 ( 
.A(n_1105),
.B(n_1064),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1040),
.B(n_1060),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1010),
.A2(n_1017),
.B(n_1058),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1130),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1028),
.Y(n_1212)
);

BUFx8_ASAP7_75t_L g1213 ( 
.A(n_1028),
.Y(n_1213)
);

CKINVDCx14_ASAP7_75t_R g1214 ( 
.A(n_1032),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_1032),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1032),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1119),
.A2(n_1017),
.B(n_1079),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_1070),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1040),
.Y(n_1219)
);

AND2x4_ASAP7_75t_SL g1220 ( 
.A(n_1107),
.B(n_1124),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1107),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1058),
.B(n_1046),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1062),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1046),
.B(n_1045),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1062),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1091),
.B(n_1097),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1039),
.B(n_1080),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1041),
.A2(n_1114),
.B1(n_998),
.B2(n_1029),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1075),
.Y(n_1229)
);

OAI21xp33_ASAP7_75t_L g1230 ( 
.A1(n_1044),
.A2(n_1077),
.B(n_1066),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1133),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_R g1232 ( 
.A(n_1072),
.B(n_1074),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1002),
.A2(n_1007),
.B(n_1140),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1073),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1068),
.B(n_1076),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1050),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1068),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1083),
.A2(n_1048),
.B1(n_1050),
.B2(n_1133),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1067),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1052),
.B(n_1065),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_1092),
.A2(n_1141),
.B(n_1136),
.C(n_1110),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1108),
.A2(n_1109),
.B(n_1054),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1051),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1071),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1003),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1093),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1093),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1024),
.B(n_1122),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1006),
.B(n_1004),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1121),
.B(n_722),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1014),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1061),
.B(n_1037),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1093),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1098),
.A2(n_919),
.B(n_877),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1121),
.B(n_722),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1061),
.B(n_1037),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1085),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1024),
.B(n_1122),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1121),
.B(n_722),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1014),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1121),
.B(n_722),
.Y(n_1262)
);

NAND2xp33_ASAP7_75t_L g1263 ( 
.A(n_1015),
.B(n_919),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1030),
.Y(n_1264)
);

BUFx12f_ASAP7_75t_L g1265 ( 
.A(n_1016),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1020),
.B(n_1061),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1121),
.B(n_722),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1003),
.Y(n_1268)
);

OAI22x1_ASAP7_75t_L g1269 ( 
.A1(n_1122),
.A2(n_1057),
.B1(n_986),
.B2(n_942),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1085),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1087),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1078),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_1020),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1042),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1098),
.A2(n_919),
.B(n_877),
.C(n_1120),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1085),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1093),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1024),
.B(n_1122),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1024),
.B(n_1122),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1121),
.B(n_722),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1122),
.A2(n_919),
.B1(n_942),
.B2(n_888),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1085),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1003),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1087),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1122),
.A2(n_919),
.B1(n_942),
.B2(n_888),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1084),
.A2(n_1088),
.B(n_1085),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1144),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1155),
.A2(n_1281),
.B1(n_1285),
.B2(n_1267),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1199),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1155),
.A2(n_1251),
.B1(n_1280),
.B2(n_1260),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1185),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_1149),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1264),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1153),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1269),
.A2(n_1256),
.B1(n_1262),
.B2(n_1164),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1148),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1156),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1164),
.A2(n_1197),
.B1(n_1147),
.B2(n_1160),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1204),
.B(n_1248),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1144),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1144),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1252),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1261),
.Y(n_1303)
);

AO22x1_ASAP7_75t_L g1304 ( 
.A1(n_1197),
.A2(n_1158),
.B1(n_1255),
.B2(n_1273),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1153),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1226),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1158),
.A2(n_1181),
.B1(n_1171),
.B2(n_1180),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1143),
.A2(n_1278),
.B1(n_1279),
.B2(n_1259),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1248),
.B(n_1247),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1173),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1159),
.A2(n_1194),
.B1(n_1195),
.B2(n_1183),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1173),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1187),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1187),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1213),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1272),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1272),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1194),
.A2(n_1195),
.B1(n_1183),
.B2(n_1182),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1249),
.A2(n_1191),
.B1(n_1203),
.B2(n_1179),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1265),
.Y(n_1320)
);

INVx6_ASAP7_75t_L g1321 ( 
.A(n_1213),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1171),
.A2(n_1263),
.B1(n_1186),
.B2(n_1170),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1154),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1254),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1174),
.A2(n_1253),
.B1(n_1150),
.B2(n_1257),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1246),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1266),
.B(n_1234),
.Y(n_1327)
);

OR2x6_ASAP7_75t_L g1328 ( 
.A(n_1266),
.B(n_1227),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1196),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1271),
.A2(n_1284),
.B1(n_1151),
.B2(n_1209),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1163),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1196),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1241),
.A2(n_1205),
.B(n_1207),
.Y(n_1333)
);

CKINVDCx11_ASAP7_75t_R g1334 ( 
.A(n_1246),
.Y(n_1334)
);

AO21x1_ASAP7_75t_L g1335 ( 
.A1(n_1275),
.A2(n_1206),
.B(n_1217),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1286),
.A2(n_1258),
.B(n_1270),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1157),
.A2(n_1192),
.B(n_1276),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1268),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1229),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1209),
.B(n_1219),
.Y(n_1340)
);

BUFx10_ASAP7_75t_L g1341 ( 
.A(n_1165),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1198),
.Y(n_1342)
);

AO21x1_ASAP7_75t_L g1343 ( 
.A1(n_1222),
.A2(n_1202),
.B(n_1238),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1211),
.A2(n_1250),
.B1(n_1176),
.B2(n_1237),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1235),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1188),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1226),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1277),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1218),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1167),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1150),
.A2(n_1253),
.B1(n_1257),
.B2(n_1193),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1218),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1210),
.B(n_1231),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1154),
.Y(n_1354)
);

CKINVDCx11_ASAP7_75t_R g1355 ( 
.A(n_1268),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1266),
.A2(n_1273),
.B1(n_1175),
.B2(n_1200),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1283),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1175),
.A2(n_1222),
.B(n_1282),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1214),
.A2(n_1224),
.B1(n_1162),
.B2(n_1236),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1243),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1168),
.A2(n_1172),
.B1(n_1165),
.B2(n_1223),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1177),
.B(n_1178),
.Y(n_1362)
);

AOI21xp33_ASAP7_75t_L g1363 ( 
.A1(n_1230),
.A2(n_1224),
.B(n_1225),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1244),
.A2(n_1228),
.B(n_1240),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1232),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1215),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1283),
.B(n_1167),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1184),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1190),
.A2(n_1216),
.B1(n_1212),
.B2(n_1201),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1208),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1220),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1245),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1239),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1221),
.B(n_1169),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1239),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1221),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1189),
.B(n_1152),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1145),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1152),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1161),
.Y(n_1380)
);

CKINVDCx11_ASAP7_75t_R g1381 ( 
.A(n_1161),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1240),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1274),
.A2(n_1233),
.B(n_1242),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1274),
.B(n_1273),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1164),
.B(n_1197),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1149),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1164),
.B(n_1197),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1164),
.B(n_1197),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1197),
.A2(n_1122),
.B1(n_942),
.B2(n_919),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1227),
.A2(n_1232),
.B(n_1206),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1155),
.A2(n_752),
.B1(n_1121),
.B2(n_687),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1273),
.B(n_1171),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1155),
.A2(n_1121),
.B1(n_752),
.B2(n_942),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1146),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1144),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1199),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1199),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1155),
.A2(n_966),
.B1(n_1122),
.B2(n_836),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1185),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1166),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1185),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1185),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1155),
.A2(n_1121),
.B1(n_942),
.B2(n_995),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1155),
.A2(n_1121),
.B1(n_752),
.B2(n_942),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1308),
.B(n_1340),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1353),
.B(n_1385),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1324),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1393),
.A2(n_1404),
.B1(n_1391),
.B2(n_1403),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1353),
.B(n_1385),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1387),
.B(n_1388),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1345),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1370),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1363),
.A2(n_1335),
.B(n_1343),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1320),
.Y(n_1414)
);

CKINVDCx6p67_ASAP7_75t_R g1415 ( 
.A(n_1320),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1289),
.B(n_1396),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1376),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1346),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1346),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1348),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1339),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1340),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1339),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1309),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1334),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1375),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1383),
.A2(n_1333),
.B(n_1300),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1292),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1328),
.B(n_1304),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1383),
.A2(n_1300),
.B(n_1287),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1287),
.A2(n_1300),
.B(n_1336),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1334),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1328),
.B(n_1304),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1375),
.Y(n_1434)
);

AOI21xp33_ASAP7_75t_L g1435 ( 
.A1(n_1389),
.A2(n_1398),
.B(n_1311),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1328),
.B(n_1327),
.Y(n_1436)
);

INVx4_ASAP7_75t_L g1437 ( 
.A(n_1377),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1310),
.Y(n_1438)
);

AO21x2_ASAP7_75t_L g1439 ( 
.A1(n_1390),
.A2(n_1359),
.B(n_1318),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1328),
.B(n_1327),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1360),
.B(n_1301),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1310),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1312),
.Y(n_1443)
);

AO31x2_ASAP7_75t_L g1444 ( 
.A1(n_1301),
.A2(n_1395),
.A3(n_1319),
.B(n_1400),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1287),
.A2(n_1336),
.B(n_1337),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1312),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1313),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1322),
.B(n_1291),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1313),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1395),
.B(n_1358),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1299),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1402),
.B(n_1399),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1401),
.B(n_1296),
.Y(n_1453)
);

AO21x1_ASAP7_75t_SL g1454 ( 
.A1(n_1307),
.A2(n_1298),
.B(n_1295),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1390),
.A2(n_1314),
.B(n_1394),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1314),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1350),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1316),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1373),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1316),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1326),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1317),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1373),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1355),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1317),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1366),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1336),
.A2(n_1337),
.B(n_1382),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1364),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1394),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1297),
.B(n_1302),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1365),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1349),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1303),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1329),
.Y(n_1474)
);

BUFx2_ASAP7_75t_SL g1475 ( 
.A(n_1326),
.Y(n_1475)
);

INVxp67_ASAP7_75t_L g1476 ( 
.A(n_1368),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1332),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1386),
.B(n_1352),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1355),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1288),
.B(n_1330),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1342),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1392),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1380),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1471),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1450),
.B(n_1344),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1451),
.B(n_1325),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1418),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1450),
.B(n_1347),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1418),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1422),
.B(n_1411),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1419),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1419),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1406),
.B(n_1347),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1408),
.A2(n_1290),
.B1(n_1294),
.B2(n_1305),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1454),
.A2(n_1294),
.B1(n_1305),
.B2(n_1351),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1406),
.B(n_1306),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1430),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1471),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1409),
.B(n_1306),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1421),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1421),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1430),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1409),
.B(n_1357),
.Y(n_1503)
);

NOR2x1_ASAP7_75t_L g1504 ( 
.A(n_1437),
.B(n_1357),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1441),
.B(n_1410),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1435),
.A2(n_1338),
.B1(n_1367),
.B2(n_1356),
.C(n_1361),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1445),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1455),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1454),
.A2(n_1327),
.B1(n_1321),
.B2(n_1362),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1410),
.B(n_1379),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1437),
.B(n_1384),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1480),
.A2(n_1327),
.B1(n_1321),
.B2(n_1362),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1411),
.B(n_1354),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1459),
.Y(n_1514)
);

AND2x2_ASAP7_75t_SL g1515 ( 
.A(n_1437),
.B(n_1376),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1431),
.B(n_1372),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1431),
.B(n_1444),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1444),
.B(n_1372),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1444),
.B(n_1354),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1455),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1439),
.A2(n_1374),
.B(n_1371),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1426),
.B(n_1434),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1444),
.B(n_1323),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1439),
.B(n_1323),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1455),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1459),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1439),
.B(n_1354),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1463),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1438),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1490),
.B(n_1407),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1495),
.A2(n_1424),
.B(n_1476),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_SL g1532 ( 
.A1(n_1495),
.A2(n_1432),
.B(n_1425),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1490),
.B(n_1420),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1505),
.B(n_1423),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1494),
.A2(n_1485),
.B1(n_1506),
.B2(n_1509),
.Y(n_1535)
);

NOR3xp33_ASAP7_75t_L g1536 ( 
.A(n_1506),
.B(n_1412),
.C(n_1461),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1501),
.B(n_1472),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1501),
.B(n_1478),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1505),
.B(n_1466),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1503),
.B(n_1464),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1494),
.A2(n_1405),
.B1(n_1448),
.B2(n_1452),
.C(n_1473),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1498),
.B(n_1453),
.Y(n_1542)
);

AOI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1486),
.A2(n_1473),
.B1(n_1453),
.B2(n_1470),
.C(n_1428),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1511),
.A2(n_1429),
.B(n_1433),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1488),
.B(n_1423),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1509),
.A2(n_1436),
.B1(n_1440),
.B2(n_1415),
.Y(n_1546)
);

OAI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1512),
.A2(n_1527),
.B1(n_1485),
.B2(n_1524),
.C(n_1521),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1498),
.B(n_1461),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1512),
.A2(n_1415),
.B1(n_1479),
.B2(n_1412),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1515),
.B(n_1417),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1488),
.B(n_1438),
.Y(n_1551)
);

AND2x2_ASAP7_75t_SL g1552 ( 
.A(n_1515),
.B(n_1468),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1514),
.Y(n_1553)
);

OAI21xp5_ASAP7_75t_SL g1554 ( 
.A1(n_1524),
.A2(n_1414),
.B(n_1483),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1524),
.A2(n_1483),
.B(n_1447),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1503),
.A2(n_1457),
.B1(n_1429),
.B2(n_1433),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1517),
.A2(n_1442),
.B1(n_1447),
.B2(n_1446),
.C(n_1449),
.Y(n_1557)
);

OA211x2_ASAP7_75t_L g1558 ( 
.A1(n_1513),
.A2(n_1416),
.B(n_1475),
.C(n_1378),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1529),
.B(n_1443),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1529),
.B(n_1446),
.Y(n_1560)
);

NOR3xp33_ASAP7_75t_L g1561 ( 
.A(n_1497),
.B(n_1460),
.C(n_1458),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1507),
.A2(n_1467),
.B(n_1427),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1484),
.B(n_1449),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1503),
.B(n_1350),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1517),
.B(n_1469),
.C(n_1465),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1484),
.B(n_1456),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1493),
.B(n_1456),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1514),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1517),
.A2(n_1462),
.B1(n_1458),
.B2(n_1469),
.C(n_1460),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1510),
.B(n_1289),
.Y(n_1570)
);

OAI221xp5_ASAP7_75t_L g1571 ( 
.A1(n_1527),
.A2(n_1369),
.B1(n_1482),
.B2(n_1462),
.C(n_1465),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1484),
.B(n_1475),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1508),
.A2(n_1413),
.B1(n_1474),
.B2(n_1477),
.C(n_1481),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1500),
.B(n_1413),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1500),
.B(n_1413),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1510),
.B(n_1396),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1510),
.B(n_1331),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1515),
.B(n_1417),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1496),
.B(n_1499),
.Y(n_1579)
);

NOR3xp33_ASAP7_75t_L g1580 ( 
.A(n_1497),
.B(n_1381),
.C(n_1434),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1552),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1553),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1568),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1562),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1565),
.B(n_1526),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1559),
.B(n_1487),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1560),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1562),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1579),
.B(n_1516),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1565),
.B(n_1487),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1557),
.B(n_1489),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1574),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1562),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1575),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1563),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1569),
.B(n_1489),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1562),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1551),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1566),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1561),
.B(n_1491),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1552),
.B(n_1504),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1567),
.B(n_1500),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1551),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1552),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1534),
.B(n_1518),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1550),
.B(n_1502),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1534),
.B(n_1518),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1537),
.Y(n_1608)
);

NAND2x1_ASAP7_75t_L g1609 ( 
.A(n_1544),
.B(n_1522),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1555),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1545),
.B(n_1518),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1572),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1539),
.B(n_1519),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1573),
.B(n_1491),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1542),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1530),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1604),
.B(n_1540),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1616),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1610),
.B(n_1533),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1604),
.B(n_1580),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1588),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1616),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1608),
.Y(n_1623)
);

NAND4xp75_ASAP7_75t_L g1624 ( 
.A(n_1614),
.B(n_1558),
.C(n_1541),
.D(n_1531),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1614),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1604),
.B(n_1564),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1588),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1582),
.Y(n_1628)
);

NAND2x1_ASAP7_75t_L g1629 ( 
.A(n_1581),
.B(n_1544),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1590),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1590),
.Y(n_1631)
);

NOR2xp67_ASAP7_75t_L g1632 ( 
.A(n_1581),
.B(n_1585),
.Y(n_1632)
);

OR2x6_ASAP7_75t_L g1633 ( 
.A(n_1609),
.B(n_1436),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_L g1634 ( 
.A(n_1585),
.B(n_1577),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1605),
.B(n_1607),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1608),
.B(n_1543),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1578),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1608),
.B(n_1538),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1610),
.B(n_1548),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1610),
.A2(n_1532),
.B1(n_1535),
.B2(n_1536),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1586),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1600),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1591),
.B(n_1526),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_SL g1644 ( 
.A(n_1585),
.B(n_1528),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1589),
.B(n_1522),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1586),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1607),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1595),
.B(n_1528),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1591),
.A2(n_1547),
.B1(n_1596),
.B2(n_1571),
.Y(n_1649)
);

OAI21xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1605),
.A2(n_1576),
.B(n_1570),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1595),
.B(n_1492),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_SL g1652 ( 
.A(n_1602),
.B(n_1554),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1600),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1607),
.B(n_1522),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1587),
.B(n_1492),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1599),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1612),
.B(n_1331),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1657),
.B(n_1596),
.Y(n_1658)
);

OR2x6_ASAP7_75t_L g1659 ( 
.A(n_1624),
.B(n_1532),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1635),
.B(n_1609),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1599),
.Y(n_1661)
);

NOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1634),
.B(n_1609),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1642),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1640),
.A2(n_1601),
.B1(n_1589),
.B2(n_1598),
.Y(n_1664)
);

OAI21xp33_ASAP7_75t_L g1665 ( 
.A1(n_1625),
.A2(n_1615),
.B(n_1587),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1621),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1653),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1651),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1655),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1615),
.Y(n_1670)
);

AND2x2_ASAP7_75t_SL g1671 ( 
.A(n_1649),
.B(n_1582),
.Y(n_1671)
);

OAI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1636),
.A2(n_1601),
.B1(n_1546),
.B2(n_1556),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_SL g1673 ( 
.A(n_1644),
.B(n_1601),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1618),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1644),
.A2(n_1549),
.B(n_1588),
.C(n_1584),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1652),
.B(n_1635),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1652),
.B(n_1647),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1626),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1622),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1619),
.B(n_1615),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1626),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1643),
.B(n_1603),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1621),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1643),
.B(n_1603),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1627),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1638),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1627),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1650),
.B(n_1599),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1623),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1628),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1647),
.B(n_1589),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1632),
.A2(n_1631),
.B(n_1630),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1639),
.B(n_1603),
.Y(n_1694)
);

O2A1O1Ixp5_ASAP7_75t_L g1695 ( 
.A1(n_1620),
.A2(n_1588),
.B(n_1606),
.C(n_1597),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1617),
.B(n_1589),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1630),
.B(n_1583),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1639),
.B(n_1631),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1617),
.B(n_1589),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1620),
.B(n_1645),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1648),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1641),
.B(n_1646),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1656),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1703),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1702),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1661),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1695),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1658),
.B(n_1293),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1702),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1661),
.A2(n_1597),
.B1(n_1593),
.B2(n_1584),
.C(n_1588),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1663),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1677),
.B(n_1700),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1659),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1671),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1671),
.Y(n_1717)
);

OAI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1659),
.A2(n_1629),
.B1(n_1597),
.B2(n_1584),
.C(n_1593),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1659),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1677),
.B(n_1654),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1681),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1687),
.B(n_1641),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1667),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1678),
.B(n_1646),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1659),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1675),
.B(n_1593),
.C(n_1584),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1698),
.B(n_1656),
.Y(n_1727)
);

OAI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1658),
.A2(n_1675),
.B1(n_1693),
.B2(n_1665),
.C(n_1662),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1690),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1691),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1690),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1660),
.B(n_1673),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1698),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1674),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1679),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1685),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1669),
.Y(n_1737)
);

AOI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1672),
.A2(n_1597),
.B1(n_1593),
.B2(n_1594),
.C(n_1592),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1668),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1666),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1706),
.B(n_1673),
.C(n_1689),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1714),
.B(n_1700),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1706),
.A2(n_1664),
.B1(n_1689),
.B2(n_1701),
.C(n_1594),
.Y(n_1743)
);

OAI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1728),
.A2(n_1629),
.B1(n_1633),
.B2(n_1601),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1721),
.B(n_1670),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1728),
.A2(n_1660),
.B1(n_1699),
.B2(n_1696),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1704),
.Y(n_1747)
);

NAND2x1p5_ASAP7_75t_L g1748 ( 
.A(n_1715),
.B(n_1315),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1717),
.A2(n_1697),
.B(n_1660),
.Y(n_1749)
);

INVxp67_ASAP7_75t_SL g1750 ( 
.A(n_1716),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1717),
.A2(n_1680),
.B1(n_1682),
.B2(n_1684),
.C(n_1633),
.Y(n_1751)
);

OAI32xp33_ASAP7_75t_L g1752 ( 
.A1(n_1716),
.A2(n_1699),
.A3(n_1696),
.B1(n_1694),
.B2(n_1601),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1707),
.A2(n_1692),
.B1(n_1637),
.B2(n_1589),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1704),
.Y(n_1754)
);

NAND2x1p5_ASAP7_75t_L g1755 ( 
.A(n_1715),
.B(n_1315),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1716),
.A2(n_1633),
.B1(n_1321),
.B2(n_1688),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1709),
.Y(n_1757)
);

AOI222xp33_ASAP7_75t_L g1758 ( 
.A1(n_1712),
.A2(n_1592),
.B1(n_1525),
.B2(n_1520),
.C1(n_1686),
.C2(n_1683),
.Y(n_1758)
);

OAI321xp33_ASAP7_75t_L g1759 ( 
.A1(n_1707),
.A2(n_1633),
.A3(n_1688),
.B1(n_1686),
.B2(n_1683),
.C(n_1666),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1734),
.B(n_1692),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1715),
.A2(n_1321),
.B1(n_1637),
.B2(n_1523),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1731),
.B(n_1613),
.Y(n_1762)
);

OAI31xp33_ASAP7_75t_L g1763 ( 
.A1(n_1707),
.A2(n_1637),
.A3(n_1520),
.B(n_1525),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1735),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1731),
.B(n_1613),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1735),
.Y(n_1766)
);

O2A1O1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1715),
.A2(n_1583),
.B(n_1611),
.C(n_1613),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1757),
.B(n_1709),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1764),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1757),
.B(n_1711),
.Y(n_1771)
);

AND2x4_ASAP7_75t_SL g1772 ( 
.A(n_1766),
.B(n_1730),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1741),
.B(n_1708),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1750),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1760),
.Y(n_1775)
);

INVx4_ASAP7_75t_L g1776 ( 
.A(n_1748),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1747),
.B(n_1711),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1749),
.B(n_1720),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1754),
.Y(n_1779)
);

OAI31xp33_ASAP7_75t_L g1780 ( 
.A1(n_1751),
.A2(n_1718),
.A3(n_1719),
.B(n_1725),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1759),
.A2(n_1712),
.B(n_1738),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1745),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1762),
.B(n_1733),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1755),
.Y(n_1784)
);

AND2x4_ASAP7_75t_SL g1785 ( 
.A(n_1761),
.B(n_1733),
.Y(n_1785)
);

NAND2xp33_ASAP7_75t_SL g1786 ( 
.A(n_1746),
.B(n_1732),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1765),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1753),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1774),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1781),
.A2(n_1726),
.B1(n_1743),
.B2(n_1763),
.C(n_1725),
.Y(n_1790)
);

AOI211xp5_ASAP7_75t_L g1791 ( 
.A1(n_1773),
.A2(n_1752),
.B(n_1744),
.C(n_1734),
.Y(n_1791)
);

OAI22xp33_ASAP7_75t_SL g1792 ( 
.A1(n_1774),
.A2(n_1718),
.B1(n_1725),
.B2(n_1719),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_SL g1793 ( 
.A1(n_1778),
.A2(n_1767),
.B(n_1736),
.Y(n_1793)
);

NAND3x1_ASAP7_75t_L g1794 ( 
.A(n_1782),
.B(n_1771),
.C(n_1769),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1780),
.B(n_1786),
.C(n_1775),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1785),
.A2(n_1738),
.B(n_1726),
.C(n_1719),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1778),
.A2(n_1736),
.B(n_1710),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1768),
.B(n_1720),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1768),
.B(n_1777),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1775),
.Y(n_1800)
);

NOR2x1_ASAP7_75t_L g1801 ( 
.A(n_1795),
.B(n_1770),
.Y(n_1801)
);

OAI322xp33_ASAP7_75t_L g1802 ( 
.A1(n_1800),
.A2(n_1782),
.A3(n_1770),
.B1(n_1787),
.B2(n_1775),
.C1(n_1788),
.C2(n_1783),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1798),
.B(n_1777),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1799),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1797),
.B(n_1777),
.Y(n_1805)
);

NOR3xp33_ASAP7_75t_L g1806 ( 
.A(n_1796),
.B(n_1776),
.C(n_1770),
.Y(n_1806)
);

NOR2x1p5_ASAP7_75t_L g1807 ( 
.A(n_1789),
.B(n_1776),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1793),
.B(n_1777),
.Y(n_1808)
);

NOR3xp33_ASAP7_75t_L g1809 ( 
.A(n_1790),
.B(n_1776),
.C(n_1784),
.Y(n_1809)
);

AND5x1_ASAP7_75t_L g1810 ( 
.A(n_1791),
.B(n_1756),
.C(n_1761),
.D(n_1785),
.E(n_1769),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1792),
.A2(n_1785),
.B1(n_1784),
.B2(n_1787),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_SL g1812 ( 
.A(n_1794),
.B(n_1776),
.C(n_1758),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1804),
.Y(n_1813)
);

NOR4xp25_ASAP7_75t_L g1814 ( 
.A(n_1802),
.B(n_1812),
.C(n_1808),
.D(n_1805),
.Y(n_1814)
);

OAI211xp5_ASAP7_75t_SL g1815 ( 
.A1(n_1801),
.A2(n_1779),
.B(n_1705),
.C(n_1710),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1803),
.B(n_1772),
.Y(n_1816)
);

OAI21xp33_ASAP7_75t_L g1817 ( 
.A1(n_1809),
.A2(n_1771),
.B(n_1772),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1806),
.B(n_1772),
.Y(n_1818)
);

NOR2xp67_ASAP7_75t_L g1819 ( 
.A(n_1811),
.B(n_1729),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1813),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1818),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1815),
.A2(n_1729),
.B1(n_1779),
.B2(n_1807),
.Y(n_1822)
);

NOR2xp67_ASAP7_75t_L g1823 ( 
.A(n_1816),
.B(n_1779),
.Y(n_1823)
);

INVxp67_ASAP7_75t_SL g1824 ( 
.A(n_1819),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1817),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1820),
.B(n_1814),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1823),
.B(n_1729),
.Y(n_1827)
);

OAI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1824),
.A2(n_1705),
.B(n_1739),
.Y(n_1828)
);

OAI211xp5_ASAP7_75t_L g1829 ( 
.A1(n_1822),
.A2(n_1293),
.B(n_1397),
.C(n_1810),
.Y(n_1829)
);

NOR2x1p5_ASAP7_75t_L g1830 ( 
.A(n_1824),
.B(n_1397),
.Y(n_1830)
);

XNOR2xp5_ASAP7_75t_L g1831 ( 
.A(n_1830),
.B(n_1821),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1826),
.B(n_1825),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1827),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1832),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1834),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1835),
.A2(n_1833),
.B1(n_1828),
.B2(n_1831),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1835),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1836),
.B(n_1829),
.Y(n_1838)
);

OA21x2_ASAP7_75t_L g1839 ( 
.A1(n_1837),
.A2(n_1723),
.B(n_1713),
.Y(n_1839)
);

AOI21xp33_ASAP7_75t_SL g1840 ( 
.A1(n_1838),
.A2(n_1740),
.B(n_1756),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1839),
.B(n_1740),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1840),
.B(n_1740),
.Y(n_1842)
);

AOI322xp5_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1841),
.A3(n_1723),
.B1(n_1713),
.B2(n_1739),
.C1(n_1737),
.C2(n_1724),
.Y(n_1843)
);

OAI221xp5_ASAP7_75t_R g1844 ( 
.A1(n_1843),
.A2(n_1727),
.B1(n_1737),
.B2(n_1724),
.C(n_1722),
.Y(n_1844)
);

AOI211xp5_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1727),
.B(n_1722),
.C(n_1341),
.Y(n_1845)
);


endmodule