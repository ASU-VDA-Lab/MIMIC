module fake_netlist_5_2198_n_1759 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1759);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1759;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_1070;
wire n_777;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_98),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_3),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_36),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_26),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_28),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_0),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_23),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_22),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_1),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_41),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_57),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_50),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_97),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_112),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_27),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_32),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_117),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_70),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_126),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_72),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_14),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_44),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_51),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_7),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_62),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_25),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_46),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_99),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_5),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_91),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_20),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_37),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_92),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_96),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_135),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_87),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_11),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_65),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_21),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_8),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_124),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_61),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_85),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_88),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_121),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_30),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_25),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_59),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_84),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_139),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_11),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_148),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_43),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_8),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_1),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_94),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_86),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_5),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_52),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_7),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_115),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_73),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_144),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_40),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_119),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_43),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_54),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_49),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_81),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_23),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_113),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_152),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_39),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_136),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_105),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_118),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_17),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_93),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_95),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_30),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_68),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_37),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_151),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_147),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_4),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_42),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_141),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_108),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_38),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_44),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_128),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_15),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_53),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_56),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_125),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_20),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_41),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_34),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_18),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_10),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_106),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_133),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_2),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_122),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_114),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_32),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_110),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_29),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_31),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_2),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_79),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_10),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_27),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_71),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_28),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_100),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_78),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_76),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_24),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_47),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_21),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_101),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_89),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_123),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_102),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_45),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_19),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_153),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_17),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_55),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_46),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_206),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_206),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_169),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_184),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_206),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_188),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_179),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_218),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_193),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_197),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_206),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_206),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_200),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_158),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_239),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_239),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_239),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_158),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_201),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_161),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_202),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_239),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_245),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_187),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_187),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_155),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_203),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_163),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_161),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_168),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_175),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_178),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_182),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_198),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_204),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_181),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_221),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_166),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_233),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_255),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_165),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_257),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_205),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_264),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_166),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_265),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_273),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_183),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_195),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_274),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_243),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_275),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_278),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_160),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_210),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_296),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_211),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_165),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_224),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_157),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_237),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_157),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_258),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_220),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_220),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_285),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_285),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_292),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_337),
.B(n_179),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_312),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_312),
.Y(n_387)
);

NOR2x1_ASAP7_75t_L g388 ( 
.A(n_308),
.B(n_227),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_309),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_319),
.B(n_227),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_322),
.B(n_219),
.Y(n_397)
);

BUFx8_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_328),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_351),
.B(n_359),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_310),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_359),
.B(n_280),
.Y(n_405)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_311),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_369),
.A2(n_217),
.B1(n_271),
.B2(n_283),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_324),
.B(n_280),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g410 ( 
.A1(n_325),
.A2(n_159),
.B(n_164),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_325),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_343),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_313),
.B(n_300),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_330),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_316),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_330),
.B(n_300),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_339),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_331),
.B(n_159),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_339),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_314),
.A2(n_189),
.B1(n_230),
.B2(n_267),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_333),
.B(n_156),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_348),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_317),
.Y(n_423)
);

AND2x2_ASAP7_75t_SL g424 ( 
.A(n_363),
.B(n_170),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_348),
.B(n_186),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_340),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_362),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_333),
.B(n_156),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_383),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_334),
.B(n_190),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_334),
.B(n_199),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_332),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_320),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_342),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_327),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_321),
.B(n_270),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_342),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_335),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_374),
.Y(n_446)
);

BUFx8_ASAP7_75t_L g447 ( 
.A(n_335),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_336),
.B(n_162),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_376),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_344),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_336),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_382),
.B(n_162),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_397),
.A2(n_315),
.B1(n_354),
.B2(n_345),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_384),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_L g457 ( 
.A1(n_385),
.A2(n_241),
.B1(n_207),
.B2(n_248),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_386),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_396),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_413),
.B(n_329),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_395),
.B(n_338),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_392),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_400),
.Y(n_468)
);

AO21x2_ASAP7_75t_L g469 ( 
.A1(n_421),
.A2(n_215),
.B(n_214),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_424),
.B(n_356),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_389),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_405),
.B(n_375),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

AO21x2_ASAP7_75t_L g480 ( 
.A1(n_421),
.A2(n_448),
.B(n_431),
.Y(n_480)
);

BUFx6f_ASAP7_75t_SL g481 ( 
.A(n_424),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_389),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_400),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_402),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_402),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_409),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_414),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_438),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_400),
.Y(n_495)
);

AND3x2_ASAP7_75t_L g496 ( 
.A(n_385),
.B(n_191),
.C(n_223),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

AND3x4_ASAP7_75t_L g498 ( 
.A(n_445),
.B(n_229),
.C(n_179),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_424),
.B(n_357),
.Y(n_499)
);

BUFx6f_ASAP7_75t_SL g500 ( 
.A(n_406),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_432),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_SL g502 ( 
.A(n_443),
.B(n_171),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_406),
.B(n_370),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_403),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_412),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_432),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_405),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_406),
.B(n_242),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_391),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_391),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_450),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_406),
.B(n_244),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_393),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_395),
.B(n_372),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_450),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_438),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_438),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_438),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_423),
.B(n_440),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_451),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_391),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_405),
.B(n_263),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_430),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_446),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_394),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_394),
.Y(n_535)
);

AOI21x1_ASAP7_75t_L g536 ( 
.A1(n_408),
.A2(n_286),
.B(n_282),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_431),
.B(n_167),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_394),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_394),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_436),
.B(n_375),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_429),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_396),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_429),
.Y(n_543)
);

BUFx8_ASAP7_75t_SL g544 ( 
.A(n_449),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_395),
.B(n_349),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_436),
.B(n_377),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_396),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_R g548 ( 
.A(n_401),
.B(n_167),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_436),
.B(n_346),
.C(n_344),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_397),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_429),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_429),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_395),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_397),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_407),
.B(n_171),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_397),
.B(n_365),
.Y(n_558)
);

INVxp33_ASAP7_75t_L g559 ( 
.A(n_393),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_442),
.B(n_398),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_425),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_429),
.Y(n_562)
);

INVxp33_ASAP7_75t_L g563 ( 
.A(n_399),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_429),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_452),
.B(n_295),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_442),
.B(n_377),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_410),
.Y(n_568)
);

CKINVDCx11_ASAP7_75t_R g569 ( 
.A(n_401),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_425),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_398),
.B(n_447),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_420),
.A2(n_172),
.B1(n_305),
.B2(n_304),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_448),
.B(n_379),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_399),
.B(n_382),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_428),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_451),
.Y(n_576)
);

NAND3xp33_ASAP7_75t_L g577 ( 
.A(n_435),
.B(n_360),
.C(n_346),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_426),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_416),
.B(n_238),
.Y(n_579)
);

NAND3xp33_ASAP7_75t_L g580 ( 
.A(n_435),
.B(n_360),
.C(n_347),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_435),
.B(n_379),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_426),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_426),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_425),
.Y(n_584)
);

AND3x1_ASAP7_75t_L g585 ( 
.A(n_428),
.B(n_381),
.C(n_380),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_433),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_416),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_416),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_410),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_452),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_425),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_433),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_445),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_425),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_433),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_437),
.Y(n_596)
);

BUFx4f_ASAP7_75t_L g597 ( 
.A(n_410),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_437),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_437),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_410),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_444),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_589),
.B(n_601),
.Y(n_603)
);

BUFx4_ASAP7_75t_L g604 ( 
.A(n_544),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_L g605 ( 
.A(n_473),
.B(n_407),
.C(n_420),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_590),
.B(n_447),
.Y(n_606)
);

INVx8_ASAP7_75t_L g607 ( 
.A(n_511),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_590),
.B(n_435),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_510),
.B(n_435),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_510),
.B(n_447),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_529),
.B(n_212),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_485),
.B(n_447),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_480),
.B(n_416),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_458),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_485),
.B(n_398),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_554),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_554),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_555),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_480),
.B(n_416),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_550),
.B(n_398),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_480),
.B(n_408),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_568),
.A2(n_410),
.B1(n_306),
.B2(n_303),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_588),
.B(n_388),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_588),
.B(n_388),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_501),
.B(n_434),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_550),
.B(n_173),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_555),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_495),
.B(n_266),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_501),
.B(n_434),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_599),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_599),
.B(n_418),
.Y(n_632)
);

OAI221xp5_ASAP7_75t_L g633 ( 
.A1(n_572),
.A2(n_441),
.B1(n_439),
.B2(n_289),
.C(n_276),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_529),
.B(n_216),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_537),
.A2(n_441),
.B(n_439),
.C(n_444),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_459),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_464),
.B(n_418),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_468),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_468),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_593),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_556),
.B(n_444),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_459),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_556),
.B(n_573),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_561),
.B(n_299),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_503),
.B(n_417),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_561),
.B(n_417),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_455),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_454),
.B(n_380),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_570),
.B(n_584),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_527),
.B(n_173),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_455),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_460),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_519),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_570),
.B(n_419),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_463),
.Y(n_655)
);

NOR2xp67_ASAP7_75t_SL g656 ( 
.A(n_571),
.B(n_174),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_519),
.Y(n_657)
);

NOR2xp67_ASAP7_75t_SL g658 ( 
.A(n_589),
.B(n_174),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_584),
.B(n_419),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_594),
.B(n_422),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_591),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_591),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_575),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_567),
.B(n_176),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_594),
.B(n_422),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_463),
.B(n_427),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_509),
.B(n_381),
.Y(n_667)
);

INVx3_ASAP7_75t_R g668 ( 
.A(n_574),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_465),
.B(n_176),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_466),
.B(n_427),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_504),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_466),
.B(n_222),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_591),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_470),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_470),
.B(n_226),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_576),
.B(n_177),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_520),
.B(n_177),
.Y(n_677)
);

BUFx5_ASAP7_75t_L g678 ( 
.A(n_515),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_460),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_558),
.B(n_180),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_509),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_574),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_559),
.B(n_229),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_563),
.B(n_347),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_560),
.B(n_350),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_587),
.B(n_231),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_565),
.A2(n_172),
.B1(n_260),
.B2(n_261),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_462),
.Y(n_688)
);

BUFx6f_ASAP7_75t_SL g689 ( 
.A(n_525),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_476),
.B(n_232),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_589),
.B(n_350),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_476),
.B(n_234),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_486),
.B(n_236),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_L g694 ( 
.A(n_529),
.B(n_240),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_591),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_581),
.B(n_352),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_568),
.A2(n_305),
.B1(n_260),
.B2(n_261),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_499),
.B(n_180),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_591),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_579),
.B(n_213),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_486),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_566),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_478),
.B(n_352),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_565),
.A2(n_268),
.B1(n_246),
.B2(n_247),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_568),
.A2(n_272),
.B1(n_301),
.B2(n_302),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_566),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_479),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_568),
.A2(n_272),
.B1(n_301),
.B2(n_302),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_488),
.B(n_492),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_585),
.B(n_213),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_488),
.B(n_249),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_492),
.B(n_250),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_585),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_493),
.B(n_251),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_462),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_493),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_471),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_471),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_478),
.B(n_253),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_565),
.B(n_253),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_565),
.A2(n_279),
.B1(n_291),
.B2(n_277),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_505),
.B(n_293),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_457),
.B(n_254),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_505),
.B(n_254),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_565),
.B(n_256),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_472),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_525),
.B(n_256),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_479),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_515),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_517),
.B(n_518),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_SL g731 ( 
.A(n_498),
.B(n_304),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_517),
.B(n_259),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_469),
.A2(n_290),
.B1(n_229),
.B2(n_367),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_508),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_518),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_521),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_521),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_581),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_540),
.B(n_546),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_496),
.B(n_259),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_601),
.B(n_262),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_525),
.B(n_262),
.Y(n_742)
);

O2A1O1Ixp5_ASAP7_75t_L g743 ( 
.A1(n_597),
.A2(n_371),
.B(n_368),
.C(n_367),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_587),
.B(n_269),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_601),
.B(n_297),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_469),
.A2(n_290),
.B1(n_368),
.B2(n_366),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_534),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_545),
.B(n_297),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_511),
.B(n_298),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_508),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_511),
.A2(n_298),
.B1(n_270),
.B2(n_364),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_534),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_549),
.B(n_371),
.C(n_366),
.Y(n_753)
);

INVx8_ASAP7_75t_L g754 ( 
.A(n_511),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_597),
.A2(n_290),
.B1(n_355),
.B2(n_353),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_535),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_535),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_578),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_597),
.A2(n_361),
.B1(n_355),
.B2(n_353),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_540),
.B(n_546),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_578),
.B(n_361),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_472),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_582),
.B(n_294),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_582),
.B(n_287),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_583),
.B(n_512),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_583),
.B(n_281),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_512),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_548),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_475),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_513),
.B(n_225),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_643),
.B(n_511),
.Y(n_771)
);

NOR2x1p5_ASAP7_75t_L g772 ( 
.A(n_750),
.B(n_530),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_702),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_768),
.B(n_526),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_681),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_629),
.B(n_516),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_702),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_SL g778 ( 
.A(n_731),
.B(n_557),
.C(n_235),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_617),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_673),
.B(n_587),
.Y(n_780)
);

BUFx12f_ASAP7_75t_L g781 ( 
.A(n_734),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_618),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_738),
.A2(n_481),
.B1(n_500),
.B2(n_516),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_619),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_628),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_706),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_629),
.B(n_516),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_729),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_739),
.B(n_638),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_768),
.B(n_481),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_706),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_637),
.B(n_516),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_735),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_739),
.B(n_682),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_639),
.B(n_516),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_696),
.B(n_549),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_662),
.A2(n_587),
.B(n_467),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_671),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_713),
.B(n_481),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_760),
.A2(n_500),
.B1(n_502),
.B2(n_498),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_736),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_737),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_605),
.A2(n_500),
.B1(n_498),
.B2(n_580),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_696),
.B(n_577),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_653),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_747),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_640),
.B(n_577),
.Y(n_807)
);

INVx5_ASAP7_75t_L g808 ( 
.A(n_603),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_673),
.B(n_587),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_608),
.B(n_580),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_752),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_653),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_756),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_626),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_759),
.B(n_647),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_605),
.A2(n_557),
.B1(n_572),
.B2(n_602),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_757),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_673),
.B(n_587),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_630),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_651),
.B(n_530),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_655),
.B(n_531),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_689),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_707),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_759),
.B(n_602),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_674),
.B(n_513),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_697),
.A2(n_600),
.B1(n_598),
.B2(n_596),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_701),
.B(n_531),
.Y(n_827)
);

INVx5_ASAP7_75t_L g828 ( 
.A(n_603),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_716),
.B(n_514),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_673),
.B(n_525),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_603),
.B(n_645),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_657),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_662),
.A2(n_547),
.B(n_467),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_682),
.B(n_683),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_631),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_661),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_707),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_713),
.B(n_575),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_703),
.B(n_541),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_758),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_657),
.B(n_185),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_707),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_709),
.B(n_528),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_767),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_689),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_607),
.B(n_569),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_769),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_613),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_691),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_684),
.B(n_575),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_609),
.B(n_538),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_649),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_668),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_623),
.B(n_538),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_707),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_697),
.A2(n_600),
.B1(n_598),
.B2(n_596),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_728),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_623),
.B(n_650),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_663),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_641),
.Y(n_860)
);

AOI221xp5_ASAP7_75t_L g861 ( 
.A1(n_687),
.A2(n_196),
.B1(n_252),
.B2(n_228),
.C(n_208),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_615),
.Y(n_862)
);

AND2x6_ASAP7_75t_SL g863 ( 
.A(n_740),
.B(n_575),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_636),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_667),
.Y(n_865)
);

NAND2x1p5_ASAP7_75t_L g866 ( 
.A(n_661),
.B(n_539),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_705),
.A2(n_539),
.B(n_592),
.C(n_586),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_678),
.B(n_541),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_691),
.B(n_479),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_730),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_685),
.Y(n_871)
);

AND2x2_ASAP7_75t_SL g872 ( 
.A(n_755),
.B(n_522),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_642),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_720),
.A2(n_533),
.B1(n_524),
.B2(n_522),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_648),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_678),
.B(n_543),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_685),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_678),
.B(n_551),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_685),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_SL g880 ( 
.A1(n_633),
.A2(n_270),
.B1(n_194),
.B2(n_4),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_646),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_650),
.B(n_586),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_676),
.B(n_524),
.Y(n_883)
);

CKINVDCx11_ASAP7_75t_R g884 ( 
.A(n_604),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_676),
.B(n_533),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_741),
.B(n_592),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_763),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_770),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_678),
.B(n_551),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_764),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_745),
.B(n_595),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_652),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_654),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_728),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_678),
.B(n_552),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_719),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_695),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_666),
.B(n_453),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_670),
.B(n_453),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_659),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_727),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_679),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_695),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_699),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_723),
.B(n_453),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_622),
.B(n_461),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_742),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_688),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_699),
.B(n_461),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_614),
.B(n_552),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_705),
.A2(n_490),
.B1(n_475),
.B2(n_477),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_660),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_665),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_708),
.A2(n_491),
.B1(n_477),
.B2(n_482),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_761),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_620),
.B(n_553),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_766),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_746),
.B(n_461),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_715),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_717),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_755),
.B(n_553),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_765),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_624),
.B(n_562),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_680),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_728),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_728),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_746),
.B(n_474),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_720),
.A2(n_564),
.B1(n_562),
.B2(n_474),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_718),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_691),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_726),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_607),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_632),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_672),
.B(n_474),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_607),
.B(n_754),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_762),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_675),
.B(n_542),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_635),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_724),
.Y(n_939)
);

NOR3xp33_ASAP7_75t_SL g940 ( 
.A(n_687),
.B(n_0),
.C(n_3),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_616),
.B(n_564),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_732),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_SL g943 ( 
.A(n_708),
.B(n_489),
.C(n_507),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_625),
.A2(n_547),
.B(n_467),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_644),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_691),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_690),
.B(n_542),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_692),
.B(n_542),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_693),
.B(n_490),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_711),
.B(n_491),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_664),
.B(n_536),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_712),
.B(n_489),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_754),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_714),
.B(n_506),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_R g955 ( 
.A(n_754),
.B(n_536),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_743),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_710),
.B(n_547),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_611),
.A2(n_547),
.B(n_467),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_691),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_958),
.A2(n_906),
.B(n_828),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_852),
.B(n_725),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_933),
.B(n_725),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_858),
.A2(n_749),
.B1(n_751),
.B2(n_722),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_784),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_945),
.B(n_621),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_932),
.B(n_612),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_854),
.A2(n_743),
.B(n_744),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_939),
.B(n_749),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_808),
.A2(n_694),
.B(n_634),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_798),
.B(n_748),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_784),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_823),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_933),
.B(n_733),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_811),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_823),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_776),
.A2(n_733),
.B1(n_704),
.B2(n_721),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_932),
.B(n_606),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_870),
.B(n_881),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_823),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_787),
.A2(n_740),
.B(n_698),
.C(n_656),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_834),
.B(n_814),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_774),
.B(n_669),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_774),
.B(n_677),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_875),
.B(n_610),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_850),
.B(n_753),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_893),
.B(n_700),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_811),
.Y(n_987)
);

AOI33xp33_ASAP7_75t_L g988 ( 
.A1(n_880),
.A2(n_753),
.A3(n_497),
.B1(n_507),
.B2(n_506),
.B3(n_487),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_808),
.A2(n_686),
.B(n_744),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_794),
.B(n_627),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_828),
.A2(n_831),
.B(n_869),
.Y(n_991)
);

AOI22x1_ASAP7_75t_L g992 ( 
.A1(n_938),
.A2(n_487),
.B1(n_482),
.B2(n_483),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_779),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_900),
.B(n_912),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_815),
.A2(n_658),
.B1(n_532),
.B2(n_523),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_781),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_913),
.B(n_497),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_860),
.B(n_484),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_SL g999 ( 
.A1(n_880),
.A2(n_6),
.B1(n_9),
.B2(n_12),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_782),
.Y(n_1000)
);

O2A1O1Ixp5_ASAP7_75t_L g1001 ( 
.A1(n_792),
.A2(n_484),
.B(n_483),
.C(n_494),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_819),
.B(n_532),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_882),
.B(n_532),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_922),
.B(n_532),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_785),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_771),
.A2(n_523),
.B1(n_494),
.B2(n_479),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_816),
.A2(n_523),
.B(n_494),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_849),
.A2(n_523),
.B1(n_494),
.B2(n_456),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_803),
.A2(n_896),
.B(n_804),
.C(n_796),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_817),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_849),
.A2(n_494),
.B1(n_456),
.B2(n_58),
.Y(n_1011)
);

NAND2xp33_ASAP7_75t_L g1012 ( 
.A(n_959),
.B(n_456),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_934),
.A2(n_456),
.B(n_48),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_789),
.B(n_456),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_833),
.A2(n_456),
.B(n_60),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_L g1016 ( 
.A(n_887),
.B(n_146),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_868),
.A2(n_145),
.B(n_143),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_817),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_823),
.Y(n_1019)
);

AO32x2_ASAP7_75t_L g1020 ( 
.A1(n_888),
.A2(n_9),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_896),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_835),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_915),
.B(n_16),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_775),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_865),
.B(n_18),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_890),
.B(n_19),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_837),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_921),
.A2(n_66),
.B(n_134),
.C(n_116),
.Y(n_1028)
);

OAI22x1_ASAP7_75t_L g1029 ( 
.A1(n_799),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_789),
.B(n_67),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_917),
.B(n_29),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_796),
.B(n_74),
.Y(n_1032)
);

INVx5_ASAP7_75t_L g1033 ( 
.A(n_837),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_942),
.B(n_31),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_788),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_837),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_937),
.A2(n_75),
.B(n_107),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_800),
.B(n_63),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_832),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_841),
.B(n_33),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_L g1041 ( 
.A(n_859),
.B(n_82),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_805),
.Y(n_1042)
);

CKINVDCx8_ASAP7_75t_R g1043 ( 
.A(n_863),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_SL g1044 ( 
.A(n_901),
.B(n_33),
.C(n_34),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_793),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_837),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_842),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_812),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_806),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_842),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_813),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_822),
.B(n_83),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_947),
.A2(n_90),
.B(n_104),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_872),
.A2(n_103),
.B1(n_142),
.B2(n_42),
.Y(n_1054)
);

INVx5_ASAP7_75t_L g1055 ( 
.A(n_842),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_839),
.B(n_45),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_839),
.B(n_35),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_842),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_825),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_838),
.B(n_35),
.Y(n_1060)
);

CKINVDCx16_ASAP7_75t_R g1061 ( 
.A(n_846),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_853),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_847),
.Y(n_1063)
);

OR2x6_ASAP7_75t_SL g1064 ( 
.A(n_845),
.B(n_907),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_838),
.B(n_790),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_804),
.A2(n_816),
.B1(n_807),
.B2(n_799),
.Y(n_1066)
);

OAI21xp33_ASAP7_75t_SL g1067 ( 
.A1(n_824),
.A2(n_872),
.B(n_810),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_857),
.Y(n_1068)
);

OA22x2_ASAP7_75t_L g1069 ( 
.A1(n_924),
.A2(n_820),
.B1(n_827),
.B2(n_821),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_829),
.Y(n_1070)
);

BUFx2_ASAP7_75t_SL g1071 ( 
.A(n_853),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_857),
.Y(n_1072)
);

AND3x1_ASAP7_75t_SL g1073 ( 
.A(n_772),
.B(n_861),
.C(n_940),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_857),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_857),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_783),
.A2(n_959),
.B1(n_927),
.B2(n_918),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_921),
.A2(n_867),
.B(n_916),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_948),
.A2(n_944),
.B(n_886),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_807),
.A2(n_790),
.B1(n_795),
.B2(n_802),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_801),
.Y(n_1080)
);

OA22x2_ASAP7_75t_L g1081 ( 
.A1(n_820),
.A2(n_827),
.B1(n_821),
.B2(n_877),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_847),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_840),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_871),
.B(n_879),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_891),
.A2(n_851),
.B(n_916),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_844),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_897),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_848),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_897),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_884),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_910),
.A2(n_954),
.B(n_952),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_SL g1092 ( 
.A(n_935),
.B(n_953),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_940),
.A2(n_885),
.B(n_883),
.C(n_830),
.Y(n_1093)
);

BUFx12f_ASAP7_75t_L g1094 ( 
.A(n_884),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_830),
.A2(n_867),
.B(n_923),
.C(n_950),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_846),
.B(n_859),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_923),
.A2(n_949),
.B(n_943),
.C(n_843),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_904),
.B(n_795),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_778),
.B(n_953),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_904),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_836),
.B(n_903),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_848),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_957),
.B(n_941),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_778),
.B(n_941),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_894),
.B(n_903),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_773),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_874),
.A2(n_905),
.B1(n_957),
.B2(n_930),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_978),
.B(n_910),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_1039),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1067),
.A2(n_905),
.B(n_951),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_972),
.Y(n_1111)
);

AO21x2_ASAP7_75t_L g1112 ( 
.A1(n_1077),
.A2(n_956),
.B(n_955),
.Y(n_1112)
);

AO21x1_ASAP7_75t_L g1113 ( 
.A1(n_963),
.A2(n_898),
.B(n_899),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1067),
.A2(n_928),
.B(n_911),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_974),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_1107),
.A2(n_909),
.A3(n_946),
.B(n_786),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_994),
.B(n_836),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_982),
.A2(n_930),
.B(n_902),
.C(n_864),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_961),
.B(n_894),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_SL g1120 ( 
.A1(n_1079),
.A2(n_786),
.B(n_855),
.Y(n_1120)
);

AO31x2_ASAP7_75t_L g1121 ( 
.A1(n_1076),
.A2(n_936),
.A3(n_931),
.B(n_908),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1078),
.A2(n_889),
.B(n_876),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1001),
.A2(n_826),
.B(n_856),
.Y(n_1123)
);

AO21x2_ASAP7_75t_L g1124 ( 
.A1(n_967),
.A2(n_1091),
.B(n_1085),
.Y(n_1124)
);

AOI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_976),
.A2(n_911),
.B(n_914),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_SL g1126 ( 
.A(n_996),
.B(n_894),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1059),
.B(n_908),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_993),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_1024),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_969),
.A2(n_878),
.B(n_889),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_983),
.A2(n_846),
.B1(n_935),
.B2(n_892),
.Y(n_1131)
);

NOR4xp25_ASAP7_75t_L g1132 ( 
.A(n_1021),
.B(n_826),
.C(n_856),
.D(n_914),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1070),
.B(n_931),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1065),
.B(n_936),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_981),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_SL g1136 ( 
.A1(n_1079),
.A2(n_855),
.B(n_797),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_972),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1060),
.A2(n_862),
.B(n_873),
.C(n_920),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1000),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_962),
.B(n_919),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1005),
.Y(n_1141)
);

NOR2xp67_ASAP7_75t_L g1142 ( 
.A(n_1048),
.B(n_929),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1012),
.A2(n_895),
.B(n_894),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_992),
.A2(n_866),
.B(n_780),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_L g1145 ( 
.A(n_1046),
.B(n_1041),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_995),
.A2(n_777),
.A3(n_791),
.B(n_955),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1022),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_985),
.B(n_935),
.Y(n_1148)
);

OAI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_986),
.A2(n_780),
.B(n_809),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_989),
.A2(n_809),
.B(n_818),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1035),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_987),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1063),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1082),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_991),
.A2(n_818),
.B(n_926),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_SL g1156 ( 
.A1(n_980),
.A2(n_925),
.B(n_926),
.C(n_1038),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1042),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1006),
.A2(n_1103),
.A3(n_1054),
.B(n_1009),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1097),
.A2(n_1007),
.B(n_1003),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1066),
.B(n_964),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1066),
.A2(n_999),
.B1(n_973),
.B2(n_1007),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1093),
.A2(n_1011),
.B(n_1032),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1013),
.A2(n_1029),
.A3(n_1101),
.B(n_1004),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1017),
.A2(n_1028),
.B(n_998),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_972),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_990),
.B(n_968),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1008),
.A2(n_997),
.B(n_1105),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1062),
.B(n_1084),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_988),
.B(n_1023),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_971),
.A2(n_1018),
.A3(n_1010),
.B(n_1053),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1088),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_966),
.B(n_977),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1069),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_999),
.A2(n_1051),
.B1(n_1049),
.B2(n_1045),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1098),
.B(n_1080),
.Y(n_1175)
);

OAI21xp33_ASAP7_75t_SL g1176 ( 
.A1(n_965),
.A2(n_984),
.B(n_1026),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1081),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_965),
.A2(n_1104),
.B(n_1056),
.C(n_1057),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1037),
.A2(n_1102),
.B(n_1014),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1083),
.Y(n_1180)
);

NOR2x1_ASAP7_75t_SL g1181 ( 
.A(n_1033),
.B(n_1055),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1031),
.A2(n_1002),
.B(n_1016),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_966),
.B(n_977),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1096),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1073),
.A2(n_1099),
.B1(n_1030),
.B2(n_1092),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_SL g1187 ( 
.A(n_1092),
.B(n_1043),
.Y(n_1187)
);

AO32x2_ASAP7_75t_L g1188 ( 
.A1(n_1020),
.A2(n_1046),
.A3(n_1044),
.B1(n_1040),
.B2(n_1034),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1016),
.A2(n_1106),
.B(n_1100),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1089),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1025),
.B(n_1071),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_975),
.A2(n_1068),
.B(n_979),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1058),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1068),
.B(n_1074),
.Y(n_1194)
);

AOI22x1_ASAP7_75t_L g1195 ( 
.A1(n_1074),
.A2(n_1047),
.B1(n_1019),
.B2(n_1075),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1019),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1033),
.A2(n_1055),
.B(n_1019),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_970),
.B(n_1055),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1033),
.A2(n_1050),
.B(n_1027),
.C(n_1036),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1027),
.B(n_1075),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1027),
.A2(n_1036),
.B1(n_1047),
.B2(n_1050),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1036),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_L g1203 ( 
.A(n_1061),
.B(n_1090),
.C(n_1047),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1050),
.B(n_1072),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1072),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1052),
.B(n_1064),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1020),
.A2(n_1094),
.B(n_1015),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1020),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_982),
.A2(n_983),
.B(n_1060),
.C(n_858),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_978),
.A2(n_858),
.B1(n_994),
.B2(n_759),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1015),
.A2(n_960),
.B(n_969),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1039),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_SL g1214 ( 
.A1(n_982),
.A2(n_605),
.B(n_880),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_978),
.B(n_994),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_982),
.A2(n_983),
.B(n_1060),
.C(n_858),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1039),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_SL g1218 ( 
.A1(n_1079),
.A2(n_1066),
.B(n_1077),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_963),
.A2(n_976),
.B(n_982),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_981),
.B(n_834),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1039),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_978),
.B(n_994),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_993),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_960),
.A2(n_1078),
.B(n_969),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1039),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1033),
.B(n_1055),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1067),
.A2(n_1077),
.B(n_1095),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1015),
.A2(n_960),
.B(n_969),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_978),
.B(n_994),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_978),
.B(n_994),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_978),
.B(n_994),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_981),
.B(n_834),
.Y(n_1232)
);

O2A1O1Ixp5_ASAP7_75t_L g1233 ( 
.A1(n_1060),
.A2(n_1065),
.B(n_983),
.C(n_982),
.Y(n_1233)
);

NOR2x1_ASAP7_75t_SL g1234 ( 
.A(n_1033),
.B(n_1055),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1107),
.A2(n_1076),
.A3(n_995),
.B(n_1078),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_960),
.A2(n_1078),
.B(n_969),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_982),
.A2(n_983),
.B(n_1060),
.C(n_858),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1039),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_982),
.A2(n_983),
.B(n_1060),
.C(n_858),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1039),
.Y(n_1240)
);

OR2x6_ASAP7_75t_L g1241 ( 
.A(n_1081),
.B(n_935),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_978),
.B(n_852),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1015),
.A2(n_960),
.B(n_969),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_978),
.B(n_852),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_981),
.B(n_834),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_SL g1246 ( 
.A1(n_982),
.A2(n_605),
.B(n_880),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_974),
.Y(n_1247)
);

AOI21x1_ASAP7_75t_L g1248 ( 
.A1(n_960),
.A2(n_1107),
.B(n_1085),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1067),
.A2(n_1077),
.B(n_1095),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1039),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_961),
.B(n_814),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1214),
.B(n_1246),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1226),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1128),
.Y(n_1254)
);

OAI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1214),
.A2(n_1246),
.B1(n_1174),
.B2(n_1229),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1112),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1172),
.B(n_1241),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_1109),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1111),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1111),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1112),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1139),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1171),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1135),
.B(n_1251),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1141),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1147),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1153),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1217),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1213),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1215),
.B(n_1222),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1172),
.B(n_1241),
.Y(n_1271)
);

AOI22x1_ASAP7_75t_L g1272 ( 
.A1(n_1189),
.A2(n_1173),
.B1(n_1159),
.B2(n_1136),
.Y(n_1272)
);

OAI21xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1219),
.A2(n_1230),
.B(n_1231),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1226),
.Y(n_1274)
);

OR2x6_ASAP7_75t_L g1275 ( 
.A(n_1241),
.B(n_1162),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1210),
.A2(n_1216),
.B(n_1237),
.C(n_1239),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1154),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1213),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1115),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1220),
.B(n_1232),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1135),
.B(n_1166),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1184),
.B(n_1177),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1144),
.A2(n_1130),
.B(n_1122),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1152),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_SL g1285 ( 
.A1(n_1189),
.A2(n_1120),
.B(n_1169),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1221),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1247),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1248),
.A2(n_1164),
.B(n_1179),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1242),
.B(n_1244),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1155),
.A2(n_1150),
.B(n_1167),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1121),
.Y(n_1291)
);

OR2x6_ASAP7_75t_L g1292 ( 
.A(n_1218),
.B(n_1148),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1151),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1225),
.Y(n_1294)
);

NAND2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1126),
.B(n_1145),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1143),
.A2(n_1249),
.B(n_1227),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1192),
.B(n_1186),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1180),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1174),
.A2(n_1161),
.B1(n_1125),
.B2(n_1249),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1227),
.A2(n_1114),
.B(n_1110),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1233),
.A2(n_1178),
.B(n_1176),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1111),
.Y(n_1302)
);

NOR3xp33_ASAP7_75t_L g1303 ( 
.A(n_1242),
.B(n_1244),
.C(n_1161),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1245),
.B(n_1140),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1191),
.B(n_1190),
.Y(n_1305)
);

AOI221xp5_ASAP7_75t_L g1306 ( 
.A1(n_1132),
.A2(n_1211),
.B1(n_1168),
.B2(n_1160),
.C(n_1182),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1192),
.A2(n_1208),
.B(n_1113),
.Y(n_1307)
);

AOI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1119),
.A2(n_1160),
.B(n_1211),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1137),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1129),
.B(n_1240),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1123),
.A2(n_1108),
.B(n_1195),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1238),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1223),
.Y(n_1313)
);

OAI211xp5_ASAP7_75t_L g1314 ( 
.A1(n_1131),
.A2(n_1182),
.B(n_1132),
.C(n_1142),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_SL g1315 ( 
.A1(n_1134),
.A2(n_1117),
.B(n_1181),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_SL g1316 ( 
.A1(n_1199),
.A2(n_1118),
.B(n_1134),
.C(n_1138),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1124),
.A2(n_1156),
.B(n_1123),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1201),
.A2(n_1117),
.B(n_1133),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1175),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1201),
.A2(n_1127),
.B(n_1133),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1127),
.B(n_1185),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1149),
.A2(n_1194),
.B(n_1193),
.Y(n_1322)
);

BUFx4f_ASAP7_75t_SL g1323 ( 
.A(n_1250),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1121),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1137),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1170),
.Y(n_1326)
);

O2A1O1Ixp5_ASAP7_75t_L g1327 ( 
.A1(n_1209),
.A2(n_1194),
.B(n_1198),
.C(n_1197),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1196),
.B(n_1205),
.Y(n_1328)
);

INVxp67_ASAP7_75t_SL g1329 ( 
.A(n_1234),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1137),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1204),
.A2(n_1206),
.B(n_1200),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1187),
.A2(n_1207),
.B(n_1203),
.C(n_1183),
.Y(n_1332)
);

NAND2xp33_ASAP7_75t_L g1333 ( 
.A(n_1165),
.B(n_1209),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1235),
.A2(n_1146),
.B(n_1116),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1202),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1170),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1165),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1183),
.A2(n_1235),
.B(n_1170),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1188),
.A2(n_1165),
.B1(n_1158),
.B2(n_1163),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1163),
.B(n_1158),
.Y(n_1340)
);

AO21x2_ASAP7_75t_L g1341 ( 
.A1(n_1146),
.A2(n_1158),
.B(n_1163),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1215),
.B(n_1222),
.Y(n_1342)
);

AOI222xp33_ASAP7_75t_L g1343 ( 
.A1(n_1214),
.A2(n_999),
.B1(n_1246),
.B2(n_407),
.C1(n_557),
.C2(n_1174),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1215),
.B(n_1222),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1214),
.A2(n_1246),
.B1(n_1174),
.B2(n_1066),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1212),
.A2(n_1243),
.B(n_1228),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1227),
.A2(n_1249),
.B(n_1219),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1171),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1212),
.A2(n_1243),
.B(n_1228),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1113),
.A2(n_1159),
.A3(n_1236),
.B(n_1224),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1219),
.A2(n_999),
.B1(n_605),
.B2(n_880),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1126),
.B(n_1033),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1224),
.A2(n_1236),
.B(n_1219),
.Y(n_1353)
);

OA21x2_ASAP7_75t_L g1354 ( 
.A1(n_1227),
.A2(n_1249),
.B(n_1219),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1171),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1174),
.A2(n_481),
.B1(n_385),
.B2(n_999),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1128),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1212),
.A2(n_1243),
.B(n_1228),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1113),
.A2(n_1159),
.A3(n_1236),
.B(n_1224),
.Y(n_1359)
);

CKINVDCx11_ASAP7_75t_R g1360 ( 
.A(n_1213),
.Y(n_1360)
);

AOI22x1_ASAP7_75t_L g1361 ( 
.A1(n_1189),
.A2(n_1029),
.B1(n_590),
.B2(n_939),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1171),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1212),
.A2(n_1243),
.B(n_1228),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1219),
.A2(n_999),
.B1(n_605),
.B2(n_880),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1210),
.A2(n_1237),
.B1(n_1239),
.B2(n_1216),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1227),
.A2(n_1249),
.B(n_1219),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1157),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1109),
.Y(n_1368)
);

OAI222xp33_ASAP7_75t_L g1369 ( 
.A1(n_1174),
.A2(n_880),
.B1(n_557),
.B2(n_1161),
.C1(n_1066),
.C2(n_633),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1219),
.A2(n_999),
.B1(n_605),
.B2(n_880),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1210),
.A2(n_1237),
.B1(n_1239),
.B2(n_1216),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1233),
.A2(n_1216),
.B(n_1210),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1212),
.A2(n_1243),
.B(n_1228),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1112),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1112),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1356),
.A2(n_1364),
.B1(n_1370),
.B2(n_1351),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1351),
.A2(n_1364),
.B1(n_1370),
.B2(n_1252),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1252),
.A2(n_1299),
.B1(n_1342),
.B2(n_1344),
.Y(n_1378)
);

CKINVDCx6p67_ASAP7_75t_R g1379 ( 
.A(n_1269),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1321),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1264),
.B(n_1304),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1299),
.A2(n_1270),
.B1(n_1345),
.B2(n_1255),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1280),
.B(n_1305),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1254),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1262),
.Y(n_1385)
);

OA22x2_ASAP7_75t_L g1386 ( 
.A1(n_1314),
.A2(n_1372),
.B1(n_1282),
.B2(n_1285),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1317),
.A2(n_1353),
.B(n_1301),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1369),
.A2(n_1343),
.B(n_1365),
.C(n_1371),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1281),
.B(n_1292),
.Y(n_1389)
);

AND2x2_ASAP7_75t_SL g1390 ( 
.A(n_1347),
.B(n_1354),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1291),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1345),
.A2(n_1255),
.B1(n_1289),
.B2(n_1361),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1338),
.A2(n_1288),
.B(n_1307),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1276),
.A2(n_1273),
.B(n_1332),
.C(n_1303),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1319),
.B(n_1306),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1265),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1269),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1300),
.B(n_1339),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1278),
.B(n_1310),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1257),
.B(n_1271),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1331),
.Y(n_1401)
);

O2A1O1Ixp5_ASAP7_75t_L g1402 ( 
.A1(n_1308),
.A2(n_1327),
.B(n_1340),
.C(n_1297),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1316),
.A2(n_1315),
.B(n_1292),
.C(n_1275),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1266),
.B(n_1293),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1296),
.A2(n_1283),
.B(n_1290),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1275),
.A2(n_1323),
.B1(n_1286),
.B2(n_1258),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1296),
.A2(n_1290),
.B(n_1300),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1331),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1258),
.A2(n_1286),
.B1(n_1323),
.B2(n_1268),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1298),
.Y(n_1410)
);

O2A1O1Ixp5_ASAP7_75t_L g1411 ( 
.A1(n_1329),
.A2(n_1336),
.B(n_1326),
.C(n_1324),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1257),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1313),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1310),
.B(n_1267),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1349),
.A2(n_1358),
.B(n_1373),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1267),
.B(n_1277),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1333),
.A2(n_1339),
.B(n_1320),
.C(n_1318),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1294),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1268),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1277),
.B(n_1287),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1335),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1357),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1279),
.B(n_1284),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1312),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1368),
.A2(n_1367),
.B1(n_1272),
.B2(n_1295),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1352),
.A2(n_1366),
.B(n_1354),
.Y(n_1426)
);

INVxp33_ASAP7_75t_L g1427 ( 
.A(n_1360),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1263),
.B(n_1348),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1348),
.Y(n_1429)
);

O2A1O1Ixp5_ASAP7_75t_L g1430 ( 
.A1(n_1274),
.A2(n_1253),
.B(n_1355),
.C(n_1362),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1328),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1360),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1318),
.B(n_1322),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1295),
.A2(n_1328),
.B(n_1256),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1341),
.B(n_1256),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1261),
.B(n_1375),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1333),
.A2(n_1374),
.B(n_1311),
.C(n_1316),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1309),
.A2(n_1330),
.B1(n_1260),
.B2(n_1259),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1334),
.B(n_1359),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1334),
.B(n_1359),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1334),
.B(n_1359),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1309),
.B(n_1330),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1350),
.B(n_1359),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1302),
.A2(n_1325),
.B1(n_1337),
.B2(n_1350),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1337),
.B(n_1346),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1337),
.B(n_1363),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1317),
.A2(n_1353),
.B(n_1301),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1369),
.A2(n_1214),
.B(n_1246),
.C(n_1216),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1269),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1270),
.A2(n_1344),
.B(n_1342),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1280),
.B(n_1305),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1252),
.B(n_1300),
.Y(n_1452)
);

INVx8_ASAP7_75t_L g1453 ( 
.A(n_1258),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1252),
.A2(n_1214),
.B(n_1246),
.C(n_1233),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1395),
.B(n_1378),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1452),
.B(n_1398),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1391),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1452),
.B(n_1398),
.Y(n_1458)
);

INVxp67_ASAP7_75t_SL g1459 ( 
.A(n_1401),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1437),
.A2(n_1417),
.B(n_1426),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1390),
.B(n_1439),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1411),
.A2(n_1402),
.B(n_1417),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1389),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1407),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1415),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1408),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1384),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1432),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1436),
.B(n_1435),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1380),
.B(n_1450),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1385),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1396),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1435),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1410),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1413),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1415),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1422),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1388),
.A2(n_1394),
.B(n_1392),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1415),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1450),
.B(n_1454),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1429),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1443),
.B(n_1387),
.Y(n_1483)
);

AOI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1382),
.A2(n_1444),
.B(n_1425),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1404),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1445),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1381),
.B(n_1399),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1419),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1433),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1387),
.B(n_1447),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1428),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1454),
.B(n_1377),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1447),
.B(n_1428),
.Y(n_1493)
);

AOI21xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1376),
.A2(n_1448),
.B(n_1406),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1428),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1421),
.B(n_1414),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1434),
.A2(n_1403),
.B(n_1446),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1416),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1420),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1405),
.B(n_1431),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1423),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1467),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1471),
.Y(n_1503)
);

CKINVDCx14_ASAP7_75t_R g1504 ( 
.A(n_1469),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1500),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1492),
.A2(n_1479),
.B1(n_1455),
.B2(n_1494),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1481),
.A2(n_1434),
.B(n_1430),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1457),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1497),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1466),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1497),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1483),
.B(n_1405),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1500),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1489),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1493),
.B(n_1400),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1465),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1489),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1463),
.B(n_1393),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1496),
.B(n_1386),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1474),
.B(n_1470),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1479),
.A2(n_1386),
.B1(n_1451),
.B2(n_1383),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1468),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1463),
.B(n_1393),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1463),
.B(n_1393),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1481),
.A2(n_1418),
.B(n_1427),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1468),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1488),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1506),
.B(n_1494),
.C(n_1455),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1506),
.A2(n_1492),
.B1(n_1460),
.B2(n_1471),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1522),
.Y(n_1530)
);

OAI221xp5_ASAP7_75t_L g1531 ( 
.A1(n_1525),
.A2(n_1484),
.B1(n_1487),
.B2(n_1397),
.C(n_1409),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_L g1532 ( 
.A(n_1525),
.B(n_1484),
.C(n_1438),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1514),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1507),
.B(n_1488),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1505),
.Y(n_1535)
);

AOI222xp33_ASAP7_75t_L g1536 ( 
.A1(n_1521),
.A2(n_1427),
.B1(n_1453),
.B2(n_1449),
.C1(n_1432),
.C2(n_1424),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1522),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1519),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1521),
.A2(n_1464),
.B1(n_1485),
.B2(n_1495),
.C(n_1491),
.Y(n_1539)
);

OAI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1519),
.A2(n_1464),
.B1(n_1412),
.B2(n_1379),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1503),
.A2(n_1485),
.B1(n_1491),
.B2(n_1495),
.C(n_1499),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1503),
.A2(n_1501),
.B1(n_1499),
.B2(n_1498),
.C(n_1486),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1514),
.B(n_1474),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1504),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1526),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1510),
.A2(n_1477),
.B(n_1480),
.Y(n_1546)
);

AND2x4_ASAP7_75t_SL g1547 ( 
.A(n_1515),
.B(n_1379),
.Y(n_1547)
);

BUFx5_ASAP7_75t_L g1548 ( 
.A(n_1508),
.Y(n_1548)
);

AOI221xp5_ASAP7_75t_L g1549 ( 
.A1(n_1507),
.A2(n_1501),
.B1(n_1486),
.B2(n_1472),
.C(n_1478),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1526),
.Y(n_1550)
);

NOR2x1_ASAP7_75t_SL g1551 ( 
.A(n_1509),
.B(n_1497),
.Y(n_1551)
);

INVxp67_ASAP7_75t_SL g1552 ( 
.A(n_1502),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1527),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_L g1554 ( 
.A(n_1509),
.B(n_1497),
.Y(n_1554)
);

OAI21xp33_ASAP7_75t_L g1555 ( 
.A1(n_1509),
.A2(n_1458),
.B(n_1456),
.Y(n_1555)
);

AOI33xp33_ASAP7_75t_L g1556 ( 
.A1(n_1505),
.A2(n_1490),
.A3(n_1473),
.B1(n_1472),
.B2(n_1475),
.B3(n_1476),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1502),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_SL g1558 ( 
.A1(n_1511),
.A2(n_1460),
.B1(n_1453),
.B2(n_1462),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1517),
.B(n_1513),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1517),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1515),
.B(n_1461),
.Y(n_1561)
);

OAI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1511),
.A2(n_1462),
.B1(n_1459),
.B2(n_1442),
.C(n_1482),
.Y(n_1562)
);

BUFx8_ASAP7_75t_L g1563 ( 
.A(n_1504),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1546),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1534),
.Y(n_1565)
);

INVx4_ASAP7_75t_SL g1566 ( 
.A(n_1534),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1554),
.B(n_1516),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1530),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1529),
.A2(n_1460),
.B(n_1534),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1546),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1538),
.B(n_1520),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1537),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1553),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1533),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1563),
.Y(n_1575)
);

INVx4_ASAP7_75t_L g1576 ( 
.A(n_1547),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1513),
.Y(n_1577)
);

INVx5_ASAP7_75t_L g1578 ( 
.A(n_1535),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1560),
.Y(n_1579)
);

BUFx8_ASAP7_75t_L g1580 ( 
.A(n_1563),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1549),
.B(n_1556),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1548),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1545),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1559),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1551),
.B(n_1561),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1559),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1550),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1528),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1557),
.Y(n_1589)
);

INVx4_ASAP7_75t_SL g1590 ( 
.A(n_1544),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_SL g1591 ( 
.A(n_1531),
.B(n_1449),
.C(n_1527),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1543),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1565),
.B(n_1558),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1570),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1585),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_R g1596 ( 
.A(n_1580),
.B(n_1453),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1581),
.B(n_1552),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1592),
.B(n_1520),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1570),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1568),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1570),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1585),
.B(n_1567),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1577),
.B(n_1513),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1568),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1570),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1581),
.B(n_1541),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1566),
.B(n_1518),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1584),
.B(n_1523),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1572),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1564),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1564),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1577),
.B(n_1456),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1572),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1566),
.B(n_1523),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1566),
.B(n_1511),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1523),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1571),
.B(n_1458),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1583),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1566),
.B(n_1524),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1578),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_R g1621 ( 
.A(n_1580),
.B(n_1453),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1588),
.B(n_1512),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1583),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1564),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1587),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1612),
.B(n_1622),
.Y(n_1626)
);

OAI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1606),
.A2(n_1588),
.B(n_1569),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1606),
.B(n_1590),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1590),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1597),
.B(n_1590),
.Y(n_1631)
);

NAND2x1p5_ASAP7_75t_L g1632 ( 
.A(n_1615),
.B(n_1576),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1612),
.B(n_1590),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1595),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1594),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1622),
.B(n_1574),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1603),
.A2(n_1591),
.B1(n_1531),
.B2(n_1569),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1595),
.B(n_1590),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1593),
.B(n_1574),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1595),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1594),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1600),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1593),
.B(n_1586),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1593),
.B(n_1586),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1571),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1617),
.B(n_1579),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1602),
.B(n_1586),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1594),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1594),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1615),
.A2(n_1591),
.B(n_1575),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1617),
.B(n_1589),
.Y(n_1651)
);

NOR2x1p5_ASAP7_75t_SL g1652 ( 
.A(n_1599),
.B(n_1582),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1604),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1620),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1604),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1609),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1609),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1598),
.B(n_1589),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1613),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1613),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1627),
.B(n_1586),
.Y(n_1661)
);

AOI222xp33_ASAP7_75t_L g1662 ( 
.A1(n_1637),
.A2(n_1539),
.B1(n_1580),
.B2(n_1562),
.C1(n_1555),
.C2(n_1575),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1660),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1638),
.B(n_1575),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1634),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1636),
.B(n_1618),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1629),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1638),
.B(n_1643),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1636),
.B(n_1618),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1639),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1643),
.B(n_1602),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1642),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1628),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1634),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1630),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1631),
.B(n_1640),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1640),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1646),
.B(n_1623),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1644),
.B(n_1602),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1654),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_SL g1681 ( 
.A(n_1644),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_SL g1682 ( 
.A(n_1650),
.B(n_1580),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1647),
.B(n_1607),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1653),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1645),
.B(n_1623),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1675),
.B(n_1673),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1665),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1677),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1681),
.A2(n_1633),
.B1(n_1632),
.B2(n_1645),
.Y(n_1689)
);

OAI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1682),
.A2(n_1632),
.B1(n_1626),
.B2(n_1657),
.C(n_1656),
.Y(n_1690)
);

AOI322xp5_ASAP7_75t_L g1691 ( 
.A1(n_1670),
.A2(n_1614),
.A3(n_1616),
.B1(n_1619),
.B2(n_1607),
.C1(n_1647),
.C2(n_1608),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1668),
.B(n_1655),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1664),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1685),
.Y(n_1694)
);

OAI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1662),
.A2(n_1626),
.B1(n_1654),
.B2(n_1532),
.C(n_1659),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1685),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1668),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1675),
.A2(n_1573),
.B1(n_1576),
.B2(n_1621),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1671),
.B(n_1651),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1667),
.Y(n_1700)
);

OAI21xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1661),
.A2(n_1620),
.B(n_1658),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1671),
.B(n_1651),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1676),
.A2(n_1536),
.B(n_1679),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1663),
.B(n_1573),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1697),
.B(n_1679),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1694),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1693),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1696),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1698),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1687),
.B(n_1674),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_SL g1711 ( 
.A(n_1686),
.B(n_1680),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1688),
.B(n_1674),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1699),
.B(n_1678),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1700),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1695),
.A2(n_1680),
.B(n_1669),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1709),
.A2(n_1690),
.B1(n_1686),
.B2(n_1702),
.Y(n_1716)
);

NAND2xp33_ASAP7_75t_L g1717 ( 
.A(n_1709),
.B(n_1596),
.Y(n_1717)
);

AOI311xp33_ASAP7_75t_L g1718 ( 
.A1(n_1715),
.A2(n_1689),
.A3(n_1701),
.B(n_1704),
.C(n_1692),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1711),
.B(n_1704),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1711),
.B(n_1703),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1707),
.Y(n_1721)
);

OAI321xp33_ASAP7_75t_L g1722 ( 
.A1(n_1705),
.A2(n_1683),
.A3(n_1672),
.B1(n_1667),
.B2(n_1684),
.C(n_1666),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1713),
.A2(n_1691),
.B1(n_1678),
.B2(n_1669),
.C(n_1666),
.Y(n_1723)
);

OAI221xp5_ASAP7_75t_SL g1724 ( 
.A1(n_1710),
.A2(n_1683),
.B1(n_1684),
.B2(n_1672),
.C(n_1635),
.Y(n_1724)
);

NAND4xp25_ASAP7_75t_L g1725 ( 
.A(n_1712),
.B(n_1536),
.C(n_1649),
.D(n_1648),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1721),
.Y(n_1726)
);

O2A1O1Ixp5_ASAP7_75t_L g1727 ( 
.A1(n_1720),
.A2(n_1708),
.B(n_1706),
.C(n_1714),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1719),
.Y(n_1728)
);

OAI21xp33_ASAP7_75t_L g1729 ( 
.A1(n_1717),
.A2(n_1652),
.B(n_1635),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1716),
.A2(n_1615),
.B1(n_1573),
.B2(n_1607),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1722),
.A2(n_1649),
.B1(n_1648),
.B2(n_1641),
.C(n_1624),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1728),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1726),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1730),
.B(n_1723),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1727),
.B(n_1718),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1729),
.A2(n_1724),
.B(n_1725),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1731),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1735),
.A2(n_1615),
.B1(n_1641),
.B2(n_1573),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1732),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1733),
.Y(n_1740)
);

OAI21xp33_ASAP7_75t_L g1741 ( 
.A1(n_1734),
.A2(n_1605),
.B(n_1599),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1735),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_L g1743 ( 
.A(n_1738),
.B(n_1737),
.C(n_1736),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1742),
.B(n_1740),
.Y(n_1744)
);

NAND4xp25_ASAP7_75t_L g1745 ( 
.A(n_1741),
.B(n_1599),
.C(n_1605),
.D(n_1601),
.Y(n_1745)
);

XNOR2xp5_ASAP7_75t_L g1746 ( 
.A(n_1743),
.B(n_1739),
.Y(n_1746)
);

OA22x2_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1744),
.B1(n_1601),
.B2(n_1605),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1747),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1747),
.A2(n_1745),
.B(n_1601),
.Y(n_1749)
);

AOI211xp5_ASAP7_75t_L g1750 ( 
.A1(n_1748),
.A2(n_1610),
.B(n_1611),
.C(n_1624),
.Y(n_1750)
);

XNOR2x1_ASAP7_75t_L g1751 ( 
.A(n_1749),
.B(n_1573),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_SL g1752 ( 
.A1(n_1751),
.A2(n_1620),
.B1(n_1573),
.B2(n_1624),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1750),
.Y(n_1753)
);

OAI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1753),
.A2(n_1610),
.B(n_1611),
.C(n_1658),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1754),
.A2(n_1752),
.B1(n_1611),
.B2(n_1610),
.Y(n_1755)
);

XNOR2xp5_ASAP7_75t_L g1756 ( 
.A(n_1755),
.B(n_1540),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1625),
.B(n_1616),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1757),
.A2(n_1614),
.B1(n_1616),
.B2(n_1619),
.Y(n_1758)
);

AOI211xp5_ASAP7_75t_L g1759 ( 
.A1(n_1758),
.A2(n_1625),
.B(n_1614),
.C(n_1619),
.Y(n_1759)
);


endmodule