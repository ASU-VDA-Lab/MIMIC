module fake_jpeg_32173_n_526 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_1),
.B(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_51),
.Y(n_137)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_52),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_16),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_56),
.Y(n_101)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_68),
.Y(n_115)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_22),
.B(n_15),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_75),
.B(n_76),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_14),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_34),
.B(n_0),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_78),
.A2(n_49),
.B1(n_21),
.B2(n_27),
.Y(n_154)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_80),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_83),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_13),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_92),
.B(n_95),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_28),
.B(n_0),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_28),
.B(n_1),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_48),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_100),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_110),
.B(n_116),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_24),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_117),
.B(n_162),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_54),
.B(n_24),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_124),
.B(n_133),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_94),
.A2(n_34),
.B1(n_25),
.B2(n_47),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_126),
.A2(n_89),
.B1(n_99),
.B2(n_88),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_60),
.A2(n_39),
.B1(n_41),
.B2(n_46),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_128),
.A2(n_46),
.B1(n_47),
.B2(n_35),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_85),
.B(n_39),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_59),
.B(n_41),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_50),
.B(n_24),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_136),
.B(n_145),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_87),
.B(n_38),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_51),
.B(n_24),
.Y(n_145)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_52),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_64),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_152),
.B(n_161),
.Y(n_188)
);

OR2x4_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_49),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_64),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_77),
.B(n_18),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_165),
.B(n_175),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_25),
.B1(n_80),
.B2(n_120),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_166),
.A2(n_186),
.B1(n_192),
.B2(n_214),
.Y(n_267)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_167),
.Y(n_270)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_168),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_101),
.A2(n_79),
.B1(n_93),
.B2(n_91),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_169),
.A2(n_220),
.B1(n_113),
.B2(n_102),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_78),
.C(n_90),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_171),
.B(n_197),
.C(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_119),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_172),
.B(n_178),
.Y(n_240)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_173),
.Y(n_258)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_108),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_176),
.Y(n_264)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_137),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_181),
.A2(n_218),
.B1(n_127),
.B2(n_159),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_21),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_191),
.Y(n_227)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_120),
.A2(n_25),
.B1(n_80),
.B2(n_46),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_108),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_187),
.B(n_199),
.Y(n_259)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_189),
.Y(n_269)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_190),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_115),
.B(n_18),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_109),
.A2(n_74),
.B1(n_73),
.B2(n_70),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_20),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_194),
.B(n_204),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_1),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_49),
.B(n_38),
.C(n_32),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_32),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_113),
.Y(n_231)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_203),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_20),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_104),
.B(n_30),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_211),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_207),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_104),
.B(n_121),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_132),
.Y(n_212)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_126),
.A2(n_47),
.B1(n_35),
.B2(n_27),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_102),
.A2(n_47),
.B1(n_35),
.B2(n_27),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_221),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_107),
.B(n_27),
.C(n_30),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_224),
.A2(n_105),
.B1(n_118),
.B2(n_142),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_225),
.B(n_231),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_229),
.A2(n_251),
.B1(n_173),
.B2(n_189),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_159),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_107),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_246),
.C(n_247),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_104),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_171),
.B(n_155),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_178),
.A2(n_214),
.B1(n_197),
.B2(n_199),
.Y(n_251)
);

OR2x6_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_200),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_252),
.B(n_27),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_206),
.B1(n_129),
.B2(n_146),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_127),
.C(n_160),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_209),
.C(n_196),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_170),
.B(n_157),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_174),
.B(n_157),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_272),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_164),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_164),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_179),
.A2(n_135),
.B(n_3),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_274),
.B(n_167),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_177),
.B(n_146),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_172),
.A2(n_135),
.B(n_3),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_275),
.Y(n_337)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_277),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_278),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_247),
.B(n_182),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_300),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_176),
.B1(n_185),
.B2(n_142),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_287),
.B1(n_313),
.B2(n_235),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_221),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_283),
.B(n_293),
.Y(n_329)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_240),
.A2(n_166),
.B(n_186),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_295),
.B(n_298),
.Y(n_333)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_180),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_316),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_236),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_291),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_292),
.B(n_296),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_227),
.B(n_168),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_253),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_258),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_297),
.B(n_306),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_190),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_299),
.A2(n_274),
.B(n_242),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_240),
.A2(n_184),
.B(n_201),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_129),
.B1(n_148),
.B2(n_118),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_301),
.A2(n_314),
.B1(n_229),
.B2(n_239),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_234),
.B(n_198),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_307),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_269),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_303),
.Y(n_350)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_304),
.Y(n_335)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_236),
.Y(n_305)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_305),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_246),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_238),
.B(n_193),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_309),
.A2(n_255),
.B1(n_248),
.B2(n_242),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_231),
.B(n_215),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_310),
.B(n_311),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_258),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_315),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_239),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_252),
.A2(n_148),
.B1(n_222),
.B2(n_210),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_237),
.B(n_206),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_252),
.A2(n_196),
.B(n_30),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_316),
.B(n_318),
.Y(n_358)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_252),
.B(n_30),
.CI(n_4),
.CON(n_318),
.SN(n_318)
);

INVx11_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_226),
.Y(n_320)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_322),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_323),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_251),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_360),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_309),
.A2(n_237),
.B1(n_256),
.B2(n_268),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_331),
.A2(n_344),
.B1(n_349),
.B2(n_134),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_341),
.A2(n_298),
.B(n_279),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_294),
.A2(n_264),
.B1(n_245),
.B2(n_232),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_345),
.A2(n_348),
.B1(n_352),
.B2(n_284),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_260),
.B(n_265),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_319),
.B(n_134),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_245),
.B1(n_232),
.B2(n_208),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_276),
.A2(n_224),
.B1(n_271),
.B2(n_241),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_295),
.A2(n_230),
.B1(n_243),
.B2(n_257),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_313),
.A2(n_269),
.B1(n_271),
.B2(n_233),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_278),
.Y(n_374)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_280),
.Y(n_357)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_292),
.B(n_244),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_359),
.B(n_300),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_280),
.B(n_244),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_355),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_361),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_362),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_363),
.A2(n_366),
.B1(n_378),
.B2(n_337),
.Y(n_404)
);

NOR2x1_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_295),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_390),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_279),
.B1(n_285),
.B2(n_290),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_370),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_331),
.A2(n_298),
.B1(n_318),
.B2(n_305),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_333),
.B(n_347),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_374),
.Y(n_396)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_281),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_376),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g376 ( 
.A(n_332),
.B(n_315),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_339),
.A2(n_286),
.B1(n_302),
.B2(n_307),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_346),
.B(n_318),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_379),
.B(n_392),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_360),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_380),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_340),
.B(n_288),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_382),
.C(n_385),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_288),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_341),
.A2(n_312),
.B(n_277),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_394),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_329),
.B(n_278),
.Y(n_384)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_326),
.B(n_291),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_326),
.B(n_330),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_389),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_308),
.Y(n_387)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_325),
.B(n_304),
.Y(n_388)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_325),
.B(n_303),
.C(n_278),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_30),
.Y(n_391)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_2),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_5),
.Y(n_393)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_393),
.Y(n_421)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_400),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_388),
.B1(n_376),
.B2(n_393),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_361),
.B(n_328),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_405),
.B(n_422),
.Y(n_448)
);

AOI22x1_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_358),
.B1(n_323),
.B2(n_334),
.Y(n_409)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_409),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_349),
.Y(n_411)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_411),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_371),
.A2(n_324),
.B1(n_336),
.B2(n_351),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_412),
.A2(n_414),
.B1(n_420),
.B2(n_394),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_366),
.A2(n_324),
.B1(n_336),
.B2(n_351),
.Y(n_414)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_377),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_424),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_363),
.A2(n_354),
.B1(n_350),
.B2(n_334),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_379),
.B(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_368),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_426),
.A2(n_427),
.B1(n_441),
.B2(n_421),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_404),
.A2(n_370),
.B1(n_380),
.B2(n_373),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_389),
.Y(n_428)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_415),
.A2(n_364),
.B1(n_383),
.B2(n_367),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_430),
.A2(n_446),
.B1(n_447),
.B2(n_414),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_378),
.Y(n_431)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_431),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_398),
.A2(n_390),
.B(n_369),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_432),
.A2(n_444),
.B(n_327),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_381),
.C(n_382),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_442),
.C(n_443),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_368),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_436),
.B(n_397),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_439),
.Y(n_470)
);

AO21x1_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_375),
.B(n_364),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_402),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_440),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_385),
.C(n_386),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_345),
.C(n_348),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_398),
.A2(n_343),
.B(n_342),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_407),
.B(n_338),
.Y(n_445)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_342),
.B1(n_338),
.B2(n_335),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_403),
.A2(n_335),
.B1(n_327),
.B2(n_343),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_448),
.B(n_406),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_452),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_451),
.B(n_456),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_437),
.B(n_413),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_454),
.A2(n_466),
.B1(n_425),
.B2(n_433),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_401),
.C(n_409),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_458),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_423),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_425),
.A2(n_430),
.B1(n_420),
.B2(n_433),
.Y(n_457)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_457),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_409),
.C(n_416),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_444),
.A2(n_411),
.B(n_421),
.Y(n_462)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_462),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_463),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_416),
.C(n_419),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_465),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_427),
.B(n_424),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_426),
.A2(n_419),
.B1(n_418),
.B2(n_417),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_446),
.B(n_412),
.C(n_400),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_8),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_438),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_459),
.Y(n_471)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_471),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_478),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_470),
.A2(n_461),
.B(n_439),
.Y(n_473)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_473),
.Y(n_490)
);

A2O1A1O1Ixp25_ASAP7_75t_L g478 ( 
.A1(n_470),
.A2(n_439),
.B(n_449),
.C(n_445),
.D(n_432),
.Y(n_478)
);

AOI321xp33_ASAP7_75t_L g479 ( 
.A1(n_469),
.A2(n_449),
.A3(n_438),
.B1(n_429),
.B2(n_435),
.C(n_9),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_468),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_480),
.B(n_464),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_451),
.A2(n_429),
.B1(n_435),
.B2(n_7),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_481),
.A2(n_482),
.B1(n_8),
.B2(n_9),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_460),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_460),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_499),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_485),
.B(n_467),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_491),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_486),
.B(n_454),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_493),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_456),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_453),
.C(n_455),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_497),
.C(n_474),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_466),
.Y(n_495)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_495),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_496),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_453),
.C(n_458),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_506),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_483),
.C(n_480),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_493),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_490),
.A2(n_477),
.B1(n_481),
.B2(n_479),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_498),
.A2(n_478),
.B(n_482),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_508),
.B(n_8),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_494),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_509),
.B(n_510),
.Y(n_517)
);

O2A1O1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_504),
.A2(n_487),
.B(n_498),
.C(n_488),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_511),
.A2(n_505),
.B(n_501),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_514),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_8),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_512),
.A2(n_500),
.B(n_502),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_515),
.A2(n_516),
.B(n_517),
.Y(n_519)
);

AOI322xp5_ASAP7_75t_L g521 ( 
.A1(n_519),
.A2(n_520),
.A3(n_508),
.B1(n_513),
.B2(n_507),
.C1(n_12),
.C2(n_11),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g520 ( 
.A(n_518),
.Y(n_520)
);

AOI21xp33_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_9),
.B(n_10),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_522),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_9),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_10),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_SL g526 ( 
.A1(n_525),
.A2(n_10),
.B(n_11),
.C(n_516),
.Y(n_526)
);


endmodule