module fake_jpeg_3305_n_173 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_0),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_50),
.B1(n_53),
.B2(n_45),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_61),
.B1(n_66),
.B2(n_58),
.Y(n_87)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_50),
.B1(n_53),
.B2(n_42),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_76),
.B1(n_43),
.B2(n_48),
.Y(n_86)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_96),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_61),
.B1(n_66),
.B2(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_57),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_57),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_45),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_69),
.B1(n_78),
.B2(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_104),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_69),
.C(n_62),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_24),
.C(n_40),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_55),
.B(n_44),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_102),
.B(n_5),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_55),
.B(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_55),
.B(n_44),
.C(n_20),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_114),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_111),
.B(n_4),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_19),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_7),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_118),
.C(n_123),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_133),
.B(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_6),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_98),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_134),
.C(n_111),
.Y(n_145)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_126),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_23),
.C(n_39),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_11),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_11),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_108),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_28),
.C(n_38),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_141),
.B(n_150),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_117),
.B(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_149),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_103),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_147),
.C(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_134),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_105),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_31),
.B(n_15),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_144),
.C(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_128),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_140),
.C(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_161),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_147),
.B(n_156),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_160),
.A2(n_154),
.B(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_166),
.B1(n_165),
.B2(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_146),
.B1(n_159),
.B2(n_21),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

AOI321xp33_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_146),
.A3(n_17),
.B1(n_27),
.B2(n_29),
.C(n_33),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_35),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_37),
.Y(n_173)
);


endmodule