module fake_jpeg_17901_n_97 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_0),
.C(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_2),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_2),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_3),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_3),
.B1(n_42),
.B2(n_41),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_39),
.B1(n_46),
.B2(n_47),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_66),
.B1(n_62),
.B2(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_46),
.B1(n_50),
.B2(n_43),
.Y(n_66)
);

OR2x4_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_7),
.Y(n_72)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_38),
.B1(n_37),
.B2(n_10),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_12),
.C(n_14),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_77),
.B1(n_64),
.B2(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_77),
.B1(n_81),
.B2(n_75),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_87),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_81),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_15),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_16),
.Y(n_92)
);

NAND4xp25_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_17),
.C(n_20),
.D(n_21),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_35),
.C(n_27),
.Y(n_94)
);

NOR4xp25_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_34),
.C(n_29),
.D(n_30),
.Y(n_95)
);

BUFx24_ASAP7_75t_SL g96 ( 
.A(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_22),
.Y(n_97)
);


endmodule