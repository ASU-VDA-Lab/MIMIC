module fake_aes_7648_n_1351 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1351);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1351;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_584;
wire n_1130;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1204;
wire n_1094;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_291), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_66), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_156), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_60), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_48), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_25), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_27), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_243), .Y(n_330) );
CKINVDCx16_ASAP7_75t_R g331 ( .A(n_26), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_6), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_75), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_219), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_74), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_186), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_22), .Y(n_337) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_125), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_299), .Y(n_339) );
CKINVDCx14_ASAP7_75t_R g340 ( .A(n_198), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_207), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_300), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_284), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_173), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_31), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_311), .Y(n_346) );
NOR2xp67_ASAP7_75t_L g347 ( .A(n_8), .B(n_89), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_131), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_149), .Y(n_349) );
NOR2xp67_ASAP7_75t_L g350 ( .A(n_40), .B(n_101), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_240), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_164), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_39), .Y(n_353) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_66), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_7), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_241), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_119), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_200), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_242), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_146), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_227), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_189), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_1), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_86), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_184), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_151), .B(n_166), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_287), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_133), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_73), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_238), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_197), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_145), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_24), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_229), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_179), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_168), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_247), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_171), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_56), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_127), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_318), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_232), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_258), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_65), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_225), .Y(n_385) );
BUFx5_ASAP7_75t_L g386 ( .A(n_53), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_122), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_155), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_259), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_80), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_139), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_61), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_23), .Y(n_393) );
CKINVDCx14_ASAP7_75t_R g394 ( .A(n_251), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_50), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_129), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_159), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_215), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_165), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_303), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_233), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_38), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_152), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_157), .Y(n_404) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_298), .B(n_192), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_294), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_20), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_279), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_0), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_272), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_249), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_289), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_153), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_212), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_169), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_50), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_6), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_223), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_75), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_280), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_213), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_322), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_321), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_320), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_116), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_230), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_53), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_302), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_163), .B(n_221), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_193), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_5), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_180), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_208), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_111), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_305), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_236), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_27), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_135), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_52), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_121), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_70), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_136), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_86), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_29), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_13), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_72), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_315), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_263), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_307), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_148), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_57), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_202), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_56), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_126), .Y(n_454) );
BUFx10_ASAP7_75t_L g455 ( .A(n_134), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_83), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_138), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_260), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_256), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_94), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_288), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_286), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_26), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_178), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_39), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_226), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_290), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_269), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_255), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_204), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_128), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_4), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_87), .Y(n_473) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_150), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_73), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_105), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_201), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_94), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_116), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_292), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_244), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_222), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_235), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_167), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_181), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_211), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_41), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_147), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_187), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_114), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_218), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_252), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_210), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_266), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_63), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_234), .Y(n_496) );
BUFx3_ASAP7_75t_L g497 ( .A(n_158), .Y(n_497) );
NOR2xp67_ASAP7_75t_L g498 ( .A(n_140), .B(n_209), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_43), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_19), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_295), .Y(n_501) );
INVxp67_ASAP7_75t_SL g502 ( .A(n_309), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_422), .B(n_430), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_386), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_455), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_343), .B(n_0), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_386), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_469), .B(n_1), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_469), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_469), .B(n_2), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_386), .Y(n_511) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_336), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_451), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_329), .B(n_2), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_369), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_386), .Y(n_516) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_342), .A2(n_120), .B(n_118), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_386), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_349), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_380), .B(n_3), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_386), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_331), .A2(n_354), .B1(n_355), .B2(n_332), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_369), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_336), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_398), .B(n_3), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_336), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_344), .B(n_4), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_375), .B(n_5), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_336), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_500), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_455), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_386), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_349), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_500), .B(n_7), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_351), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_342), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_378), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_332), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_471), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_539) );
INVx6_ASAP7_75t_L g540 ( .A(n_455), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_337), .B(n_9), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_337), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_355), .Y(n_543) );
CKINVDCx11_ASAP7_75t_R g544 ( .A(n_327), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_351), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_401), .B(n_325), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_505), .B(n_338), .Y(n_547) );
INVx6_ASAP7_75t_L g548 ( .A(n_508), .Y(n_548) );
BUFx2_ASAP7_75t_L g549 ( .A(n_538), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_503), .B(n_406), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_508), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_508), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_504), .Y(n_553) );
BUFx3_ASAP7_75t_L g554 ( .A(n_508), .Y(n_554) );
OR2x6_ASAP7_75t_L g555 ( .A(n_539), .B(n_347), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_512), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_538), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_522), .A2(n_514), .B1(n_534), .B2(n_541), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_503), .B(n_373), .Y(n_559) );
BUFx10_ASAP7_75t_L g560 ( .A(n_540), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_543), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_504), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_513), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_512), .Y(n_564) );
BUFx4f_ASAP7_75t_L g565 ( .A(n_510), .Y(n_565) );
BUFx10_ASAP7_75t_L g566 ( .A(n_540), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_530), .B(n_378), .Y(n_567) );
INVx4_ASAP7_75t_L g568 ( .A(n_510), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_505), .B(n_339), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_507), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_512), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_512), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_533), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_515), .B(n_340), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_533), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_533), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_544), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_533), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_531), .B(n_373), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_533), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_515), .B(n_340), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_507), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_505), .B(n_377), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_510), .Y(n_584) );
INVx4_ASAP7_75t_L g585 ( .A(n_510), .Y(n_585) );
INVx3_ASAP7_75t_L g586 ( .A(n_541), .Y(n_586) );
BUFx10_ASAP7_75t_L g587 ( .A(n_540), .Y(n_587) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_539), .A2(n_472), .B1(n_479), .B2(n_327), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_513), .A2(n_437), .B1(n_444), .B2(n_379), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_514), .A2(n_471), .B1(n_456), .B2(n_463), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_565), .B(n_534), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_579), .B(n_531), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g593 ( .A1(n_588), .A2(n_479), .B1(n_487), .B2(n_472), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_568), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_563), .B(n_530), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_558), .B(n_531), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_563), .B(n_557), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_577), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g599 ( .A1(n_559), .A2(n_528), .B(n_527), .C(n_523), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_586), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_586), .A2(n_541), .B1(n_534), .B2(n_511), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_574), .B(n_531), .Y(n_602) );
AND2x6_ASAP7_75t_SL g603 ( .A(n_555), .B(n_546), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_568), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_574), .B(n_540), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_568), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_581), .B(n_540), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_581), .B(n_523), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_567), .B(n_527), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_557), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_567), .B(n_528), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_583), .B(n_520), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_550), .B(n_520), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_549), .B(n_534), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_558), .A2(n_541), .B1(n_506), .B2(n_525), .Y(n_615) );
AND2x6_ASAP7_75t_SL g616 ( .A(n_555), .B(n_525), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_555), .A2(n_456), .B1(n_463), .B2(n_446), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_586), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_569), .B(n_542), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_568), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_586), .Y(n_621) );
AND3x1_ASAP7_75t_L g622 ( .A(n_590), .B(n_328), .C(n_326), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_565), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_548), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_561), .B(n_446), .Y(n_625) );
BUFx3_ASAP7_75t_L g626 ( .A(n_561), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_585), .B(n_519), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_565), .B(n_511), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_585), .B(n_519), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_585), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_554), .B(n_339), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_554), .B(n_383), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_547), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_548), .B(n_542), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_548), .B(n_420), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g636 ( .A1(n_555), .A2(n_487), .B1(n_476), .B2(n_390), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_551), .B(n_516), .Y(n_637) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_548), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_551), .B(n_387), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_548), .A2(n_407), .B1(n_409), .B2(n_364), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_551), .B(n_387), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_590), .A2(n_427), .B1(n_335), .B2(n_345), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_551), .B(n_436), .Y(n_643) );
NOR2x1p5_ASAP7_75t_L g644 ( .A(n_589), .B(n_324), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_552), .B(n_436), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_552), .B(n_495), .C(n_490), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_552), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_584), .B(n_438), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_584), .B(n_438), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_584), .B(n_442), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_584), .B(n_442), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_553), .A2(n_353), .B1(n_363), .B2(n_333), .Y(n_652) );
INVx4_ASAP7_75t_L g653 ( .A(n_560), .Y(n_653) );
NAND3xp33_ASAP7_75t_SL g654 ( .A(n_553), .B(n_458), .C(n_454), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_566), .B(n_454), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_566), .Y(n_656) );
INVx4_ASAP7_75t_L g657 ( .A(n_566), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_566), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_562), .A2(n_518), .B1(n_532), .B2(n_521), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_562), .A2(n_521), .B1(n_532), .B2(n_536), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_570), .A2(n_499), .B1(n_392), .B2(n_395), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_587), .B(n_458), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_587), .B(n_459), .Y(n_663) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_587), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_570), .A2(n_536), .B1(n_537), .B2(n_509), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_582), .B(n_330), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_582), .B(n_461), .Y(n_667) );
INVx2_ASAP7_75t_SL g668 ( .A(n_573), .Y(n_668) );
INVx8_ASAP7_75t_L g669 ( .A(n_556), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_575), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_575), .A2(n_393), .B1(n_416), .B2(n_402), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_576), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_576), .B(n_509), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_576), .B(n_466), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_578), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_594), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_626), .B(n_509), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_637), .A2(n_517), .B(n_578), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_637), .A2(n_517), .B(n_578), .Y(n_679) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_664), .Y(n_680) );
NOR2x1p5_ASAP7_75t_SL g681 ( .A(n_647), .B(n_429), .Y(n_681) );
BUFx8_ASAP7_75t_L g682 ( .A(n_597), .Y(n_682) );
O2A1O1Ixp5_ASAP7_75t_L g683 ( .A1(n_591), .A2(n_474), .B(n_502), .C(n_367), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_591), .A2(n_517), .B(n_580), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_628), .A2(n_517), .B(n_580), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g686 ( .A(n_610), .B(n_350), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_609), .B(n_466), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_628), .A2(n_517), .B(n_580), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_625), .B(n_417), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_612), .A2(n_537), .B(n_431), .C(n_441), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_642), .A2(n_443), .B(n_445), .C(n_419), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_611), .B(n_613), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_612), .B(n_468), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_653), .B(n_468), .Y(n_694) );
NOR2xp33_ASAP7_75t_R g695 ( .A(n_598), .B(n_394), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_595), .B(n_453), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_601), .A2(n_394), .B1(n_483), .B2(n_481), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_633), .B(n_465), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_627), .A2(n_341), .B(n_334), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_601), .A2(n_483), .B1(n_484), .B2(n_481), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_636), .A2(n_475), .B1(n_478), .B2(n_473), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_604), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_606), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_608), .B(n_614), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_629), .A2(n_348), .B(n_346), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_644), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_593), .Y(n_707) );
BUFx3_ASAP7_75t_L g708 ( .A(n_638), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_615), .A2(n_488), .B1(n_501), .B2(n_484), .Y(n_709) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_596), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_592), .A2(n_356), .B(n_352), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_639), .A2(n_361), .B(n_358), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_622), .A2(n_646), .B1(n_619), .B2(n_618), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_599), .A2(n_390), .B(n_425), .C(n_384), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_653), .B(n_488), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_641), .A2(n_368), .B(n_362), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_620), .Y(n_717) );
NOR2xp67_ASAP7_75t_L g718 ( .A(n_617), .B(n_501), .Y(n_718) );
NAND2x1p5_ASAP7_75t_L g719 ( .A(n_657), .B(n_434), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_602), .B(n_460), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_640), .B(n_385), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_623), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_621), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_646), .A2(n_371), .B1(n_372), .B2(n_370), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_634), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_605), .B(n_460), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_607), .B(n_323), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_630), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_643), .A2(n_648), .B(n_645), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_667), .B(n_357), .Y(n_730) );
O2A1O1Ixp33_ASAP7_75t_L g731 ( .A1(n_636), .A2(n_374), .B(n_382), .C(n_376), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_623), .A2(n_439), .B1(n_545), .B2(n_535), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_657), .B(n_359), .Y(n_733) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_664), .Y(n_734) );
AO21x1_ASAP7_75t_L g735 ( .A1(n_666), .A2(n_391), .B(n_389), .Y(n_735) );
O2A1O1Ixp33_ASAP7_75t_L g736 ( .A1(n_652), .A2(n_397), .B(n_408), .C(n_403), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_649), .A2(n_411), .B(n_410), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_650), .A2(n_414), .B(n_412), .Y(n_738) );
OA22x2_ASAP7_75t_L g739 ( .A1(n_661), .A2(n_418), .B1(n_421), .B2(n_415), .Y(n_739) );
INVx5_ASAP7_75t_L g740 ( .A(n_623), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_664), .B(n_360), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_651), .A2(n_432), .B(n_423), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_619), .B(n_365), .Y(n_743) );
NOR2xp33_ASAP7_75t_SL g744 ( .A(n_664), .B(n_388), .Y(n_744) );
BUFx3_ASAP7_75t_L g745 ( .A(n_638), .Y(n_745) );
INVx4_ASAP7_75t_L g746 ( .A(n_623), .Y(n_746) );
NOR2xp67_ASAP7_75t_L g747 ( .A(n_654), .B(n_10), .Y(n_747) );
OAI22x1_ASAP7_75t_L g748 ( .A1(n_603), .A2(n_428), .B1(n_424), .B2(n_433), .Y(n_748) );
OAI21xp33_ASAP7_75t_L g749 ( .A1(n_665), .A2(n_440), .B(n_435), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_659), .A2(n_448), .B(n_447), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_631), .A2(n_450), .B(n_449), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g752 ( .A1(n_635), .A2(n_462), .B(n_464), .C(n_457), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_624), .B(n_467), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g754 ( .A1(n_635), .A2(n_477), .B(n_480), .C(n_470), .Y(n_754) );
NOR2xp67_ASAP7_75t_L g755 ( .A(n_671), .B(n_11), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g756 ( .A1(n_660), .A2(n_485), .B(n_486), .C(n_482), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_632), .A2(n_492), .B(n_491), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_666), .A2(n_494), .B1(n_493), .B2(n_399), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_638), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_655), .B(n_396), .Y(n_760) );
OAI22x1_ASAP7_75t_L g761 ( .A1(n_616), .A2(n_399), .B1(n_400), .B2(n_396), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_662), .B(n_400), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_660), .A2(n_665), .B1(n_659), .B2(n_663), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_674), .A2(n_413), .B(n_404), .Y(n_764) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_669), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_663), .B(n_496), .Y(n_766) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_656), .A2(n_439), .B1(n_496), .B2(n_381), .Y(n_767) );
BUFx6f_ASAP7_75t_L g768 ( .A(n_669), .Y(n_768) );
OR2x6_ASAP7_75t_SL g769 ( .A(n_673), .B(n_11), .Y(n_769) );
BUFx2_ASAP7_75t_L g770 ( .A(n_658), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_668), .B(n_12), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_672), .Y(n_772) );
AO21x1_ASAP7_75t_L g773 ( .A1(n_670), .A2(n_526), .B(n_524), .Y(n_773) );
INVx2_ASAP7_75t_SL g774 ( .A(n_669), .Y(n_774) );
A2O1A1Ixp33_ASAP7_75t_L g775 ( .A1(n_675), .A2(n_405), .B(n_498), .C(n_452), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_626), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_594), .Y(n_777) );
A2O1A1Ixp33_ASAP7_75t_L g778 ( .A1(n_612), .A2(n_426), .B(n_489), .C(n_452), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_609), .B(n_535), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g780 ( .A1(n_637), .A2(n_571), .B(n_564), .Y(n_780) );
NOR3xp33_ASAP7_75t_L g781 ( .A(n_593), .B(n_366), .C(n_426), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_596), .A2(n_545), .B1(n_535), .B2(n_497), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_612), .A2(n_497), .B(n_489), .C(n_524), .Y(n_783) );
NOR3xp33_ASAP7_75t_L g784 ( .A(n_593), .B(n_526), .C(n_524), .Y(n_784) );
O2A1O1Ixp33_ASAP7_75t_L g785 ( .A1(n_642), .A2(n_529), .B(n_526), .C(n_564), .Y(n_785) );
O2A1O1Ixp33_ASAP7_75t_L g786 ( .A1(n_642), .A2(n_529), .B(n_571), .C(n_14), .Y(n_786) );
NOR2xp67_ASAP7_75t_L g787 ( .A(n_626), .B(n_12), .Y(n_787) );
A2O1A1Ixp33_ASAP7_75t_L g788 ( .A1(n_612), .A2(n_572), .B(n_556), .C(n_15), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_600), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_609), .A2(n_15), .B1(n_13), .B2(n_14), .Y(n_790) );
A2O1A1Ixp33_ASAP7_75t_L g791 ( .A1(n_612), .A2(n_572), .B(n_556), .C(n_18), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_610), .B(n_16), .Y(n_792) );
AND2x4_ASAP7_75t_L g793 ( .A(n_626), .B(n_16), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_626), .B(n_572), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_609), .B(n_17), .Y(n_795) );
AO22x1_ASAP7_75t_L g796 ( .A1(n_626), .A2(n_19), .B1(n_17), .B2(n_18), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_626), .B(n_20), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_609), .B(n_21), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_609), .B(n_21), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_SL g800 ( .A1(n_592), .A2(n_572), .B(n_123), .C(n_124), .Y(n_800) );
BUFx6f_ASAP7_75t_L g801 ( .A(n_664), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_626), .B(n_22), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_646), .B(n_23), .C(n_24), .Y(n_803) );
NAND2xp5_ASAP7_75t_SL g804 ( .A(n_626), .B(n_25), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_610), .B(n_28), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_626), .B(n_28), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_692), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_677), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_684), .A2(n_30), .B(n_31), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_704), .B(n_32), .Y(n_810) );
AO31x2_ASAP7_75t_L g811 ( .A1(n_788), .A2(n_34), .A3(n_32), .B(n_33), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_729), .A2(n_34), .B(n_35), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_707), .A2(n_37), .B1(n_35), .B2(n_36), .Y(n_813) );
OAI21xp5_ASAP7_75t_L g814 ( .A1(n_685), .A2(n_36), .B(n_37), .Y(n_814) );
INVxp67_ASAP7_75t_L g815 ( .A(n_776), .Y(n_815) );
INVx1_ASAP7_75t_SL g816 ( .A(n_793), .Y(n_816) );
BUFx3_ASAP7_75t_L g817 ( .A(n_682), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_795), .Y(n_818) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_688), .A2(n_38), .B(n_40), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_763), .A2(n_43), .B1(n_41), .B2(n_42), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_713), .B(n_42), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_763), .A2(n_46), .B1(n_44), .B2(n_45), .Y(n_822) );
AO22x2_ASAP7_75t_L g823 ( .A1(n_793), .A2(n_46), .B1(n_44), .B2(n_45), .Y(n_823) );
AO31x2_ASAP7_75t_L g824 ( .A1(n_791), .A2(n_49), .A3(n_47), .B(n_48), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_798), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_682), .B(n_49), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_799), .A2(n_54), .B1(n_51), .B2(n_52), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_689), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_726), .Y(n_829) );
INVx2_ASAP7_75t_SL g830 ( .A(n_695), .Y(n_830) );
AO31x2_ASAP7_75t_L g831 ( .A1(n_773), .A2(n_55), .A3(n_51), .B(n_54), .Y(n_831) );
O2A1O1Ixp33_ASAP7_75t_SL g832 ( .A1(n_714), .A2(n_132), .B(n_137), .C(n_130), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_676), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_720), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_797), .Y(n_835) );
A2O1A1Ixp33_ASAP7_75t_L g836 ( .A1(n_681), .A2(n_58), .B(n_59), .C(n_60), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g837 ( .A1(n_678), .A2(n_142), .B(n_141), .Y(n_837) );
AND2x2_ASAP7_75t_L g838 ( .A(n_769), .B(n_59), .Y(n_838) );
O2A1O1Ixp33_ASAP7_75t_L g839 ( .A1(n_690), .A2(n_61), .B(n_62), .C(n_63), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_706), .B(n_64), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_802), .Y(n_841) );
O2A1O1Ixp33_ASAP7_75t_L g842 ( .A1(n_752), .A2(n_64), .B(n_65), .C(n_67), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_679), .A2(n_144), .B(n_143), .Y(n_843) );
BUFx3_ASAP7_75t_L g844 ( .A(n_765), .Y(n_844) );
OAI21xp5_ASAP7_75t_L g845 ( .A1(n_756), .A2(n_67), .B(n_68), .Y(n_845) );
OAI21x1_ASAP7_75t_SL g846 ( .A1(n_750), .A2(n_68), .B(n_69), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_710), .B(n_69), .Y(n_847) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_680), .Y(n_848) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_765), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_761), .Y(n_850) );
OAI21xp5_ASAP7_75t_L g851 ( .A1(n_786), .A2(n_71), .B(n_72), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_753), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_784), .A2(n_71), .B1(n_74), .B2(n_76), .Y(n_853) );
AO31x2_ASAP7_75t_L g854 ( .A1(n_778), .A2(n_76), .A3(n_77), .B(n_78), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_779), .Y(n_855) );
INVx3_ASAP7_75t_L g856 ( .A(n_765), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g857 ( .A1(n_780), .A2(n_160), .B(n_154), .Y(n_857) );
OA21x2_ASAP7_75t_L g858 ( .A1(n_783), .A2(n_162), .B(n_161), .Y(n_858) );
AOI221x1_ASAP7_75t_L g859 ( .A1(n_775), .A2(n_77), .B1(n_78), .B2(n_79), .C(n_80), .Y(n_859) );
NOR4xp25_ASAP7_75t_L g860 ( .A(n_731), .B(n_79), .C(n_81), .D(n_82), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g861 ( .A1(n_766), .A2(n_172), .B(n_170), .Y(n_861) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_768), .B(n_81), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_713), .B(n_82), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_760), .A2(n_175), .B(n_174), .Y(n_864) );
A2O1A1Ixp33_ASAP7_75t_L g865 ( .A1(n_712), .A2(n_737), .B(n_738), .C(n_716), .Y(n_865) );
AO32x2_ASAP7_75t_L g866 ( .A1(n_767), .A2(n_83), .A3(n_84), .B1(n_85), .B2(n_87), .Y(n_866) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_762), .A2(n_177), .B(n_176), .Y(n_867) );
NAND2xp5_ASAP7_75t_SL g868 ( .A(n_768), .B(n_84), .Y(n_868) );
OAI21xp5_ASAP7_75t_L g869 ( .A1(n_683), .A2(n_183), .B(n_182), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_687), .B(n_85), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g871 ( .A1(n_742), .A2(n_239), .B(n_317), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_723), .Y(n_872) );
AND2x4_ASAP7_75t_L g873 ( .A(n_740), .B(n_88), .Y(n_873) );
BUFx10_ASAP7_75t_L g874 ( .A(n_768), .Y(n_874) );
OAI22x1_ASAP7_75t_L g875 ( .A1(n_724), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_875) );
OAI21xp5_ASAP7_75t_L g876 ( .A1(n_711), .A2(n_90), .B(n_91), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_696), .B(n_92), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_702), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_693), .B(n_92), .Y(n_879) );
NAND2xp5_ASAP7_75t_SL g880 ( .A(n_744), .B(n_93), .Y(n_880) );
A2O1A1Ixp33_ASAP7_75t_L g881 ( .A1(n_751), .A2(n_93), .B(n_95), .C(n_96), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_725), .B(n_95), .Y(n_882) );
AO21x2_ASAP7_75t_L g883 ( .A1(n_800), .A2(n_246), .B(n_316), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g884 ( .A1(n_730), .A2(n_245), .B(n_314), .Y(n_884) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_680), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_701), .B(n_96), .Y(n_886) );
NOR2xp67_ASAP7_75t_L g887 ( .A(n_740), .B(n_185), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_757), .A2(n_237), .B(n_313), .Y(n_888) );
BUFx12f_ASAP7_75t_L g889 ( .A(n_686), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_718), .B(n_97), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_740), .B(n_98), .Y(n_891) );
BUFx6f_ASAP7_75t_L g892 ( .A(n_680), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_709), .B(n_99), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_724), .B(n_99), .Y(n_894) );
O2A1O1Ixp5_ASAP7_75t_SL g895 ( .A1(n_804), .A2(n_231), .B(n_312), .C(n_310), .Y(n_895) );
OAI22x1_ASAP7_75t_L g896 ( .A1(n_792), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_703), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_772), .A2(n_228), .B(n_308), .Y(n_898) );
OR2x2_ASAP7_75t_L g899 ( .A(n_700), .B(n_100), .Y(n_899) );
OAI21xp5_ASAP7_75t_L g900 ( .A1(n_789), .A2(n_102), .B(n_103), .Y(n_900) );
O2A1O1Ixp33_ASAP7_75t_SL g901 ( .A1(n_794), .A2(n_248), .B(n_306), .C(n_304), .Y(n_901) );
AO31x2_ASAP7_75t_L g902 ( .A1(n_735), .A2(n_103), .A3(n_104), .B(n_105), .Y(n_902) );
INVx2_ASAP7_75t_SL g903 ( .A(n_719), .Y(n_903) );
AND2x4_ASAP7_75t_L g904 ( .A(n_770), .B(n_106), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_739), .B(n_106), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g906 ( .A1(n_755), .A2(n_107), .B1(n_108), .B2(n_109), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g907 ( .A1(n_727), .A2(n_253), .B(n_301), .Y(n_907) );
OA21x2_ASAP7_75t_L g908 ( .A1(n_764), .A2(n_250), .B(n_297), .Y(n_908) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_734), .Y(n_909) );
BUFx2_ASAP7_75t_L g910 ( .A(n_774), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_691), .B(n_107), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_698), .B(n_108), .Y(n_912) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_767), .Y(n_913) );
BUFx2_ASAP7_75t_L g914 ( .A(n_746), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_721), .B(n_109), .Y(n_915) );
AOI21xp5_ASAP7_75t_L g916 ( .A1(n_743), .A2(n_254), .B(n_296), .Y(n_916) );
INVx1_ASAP7_75t_SL g917 ( .A(n_734), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_790), .Y(n_918) );
INVx2_ASAP7_75t_SL g919 ( .A(n_806), .Y(n_919) );
NAND2xp5_ASAP7_75t_SL g920 ( .A(n_801), .B(n_110), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_699), .A2(n_224), .B(n_293), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_705), .A2(n_220), .B(n_285), .Y(n_922) );
O2A1O1Ixp33_ASAP7_75t_L g923 ( .A1(n_736), .A2(n_110), .B(n_111), .C(n_112), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_697), .B(n_112), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_717), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_749), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_926) );
OAI21xp5_ASAP7_75t_L g927 ( .A1(n_785), .A2(n_115), .B(n_117), .Y(n_927) );
AOI211x1_ASAP7_75t_L g928 ( .A1(n_796), .A2(n_117), .B(n_188), .C(n_190), .Y(n_928) );
BUFx3_ASAP7_75t_L g929 ( .A(n_708), .Y(n_929) );
BUFx6f_ASAP7_75t_L g930 ( .A(n_801), .Y(n_930) );
NAND3xp33_ASAP7_75t_SL g931 ( .A(n_781), .B(n_191), .C(n_194), .Y(n_931) );
BUFx3_ASAP7_75t_L g932 ( .A(n_745), .Y(n_932) );
A2O1A1Ixp33_ASAP7_75t_L g933 ( .A1(n_749), .A2(n_195), .B(n_196), .C(n_199), .Y(n_933) );
INVx2_ASAP7_75t_SL g934 ( .A(n_748), .Y(n_934) );
A2O1A1Ixp33_ASAP7_75t_L g935 ( .A1(n_787), .A2(n_203), .B(n_205), .C(n_206), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_805), .A2(n_214), .B1(n_216), .B2(n_217), .Y(n_936) );
OAI21xp5_ASAP7_75t_L g937 ( .A1(n_758), .A2(n_782), .B(n_728), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_758), .B(n_257), .Y(n_938) );
OA21x2_ASAP7_75t_L g939 ( .A1(n_782), .A2(n_261), .B(n_262), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_801), .A2(n_771), .B1(n_777), .B2(n_803), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_747), .Y(n_941) );
OAI21xp5_ASAP7_75t_L g942 ( .A1(n_759), .A2(n_264), .B(n_265), .Y(n_942) );
OA21x2_ASAP7_75t_L g943 ( .A1(n_732), .A2(n_267), .B(n_268), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_722), .A2(n_270), .B1(n_271), .B2(n_273), .Y(n_944) );
AND2x4_ASAP7_75t_L g945 ( .A(n_733), .B(n_319), .Y(n_945) );
OAI21x1_ASAP7_75t_L g946 ( .A1(n_741), .A2(n_274), .B(n_275), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_694), .Y(n_947) );
BUFx2_ASAP7_75t_L g948 ( .A(n_715), .Y(n_948) );
A2O1A1Ixp33_ASAP7_75t_L g949 ( .A1(n_729), .A2(n_276), .B(n_277), .C(n_278), .Y(n_949) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_729), .A2(n_281), .B(n_282), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_692), .B(n_283), .Y(n_951) );
AOI21xp5_ASAP7_75t_L g952 ( .A1(n_729), .A2(n_565), .B(n_684), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_692), .B(n_626), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_676), .Y(n_954) );
INVx2_ASAP7_75t_L g955 ( .A(n_676), .Y(n_955) );
INVxp67_ASAP7_75t_L g956 ( .A(n_692), .Y(n_956) );
INVx2_ASAP7_75t_SL g957 ( .A(n_682), .Y(n_957) );
OAI22x1_ASAP7_75t_L g958 ( .A1(n_793), .A2(n_590), .B1(n_610), .B2(n_577), .Y(n_958) );
O2A1O1Ixp33_ASAP7_75t_L g959 ( .A1(n_714), .A2(n_690), .B(n_754), .C(n_752), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_956), .Y(n_960) );
NAND2x1p5_ASAP7_75t_L g961 ( .A(n_817), .B(n_957), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_807), .B(n_953), .Y(n_962) );
BUFx2_ASAP7_75t_L g963 ( .A(n_844), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_872), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_833), .Y(n_965) );
BUFx12f_ASAP7_75t_L g966 ( .A(n_889), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_828), .Y(n_967) );
AOI21xp5_ASAP7_75t_L g968 ( .A1(n_865), .A2(n_951), .B(n_825), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_834), .B(n_829), .Y(n_969) );
BUFx2_ASAP7_75t_R g970 ( .A(n_850), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_905), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_823), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_823), .Y(n_973) );
INVx2_ASAP7_75t_L g974 ( .A(n_878), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_918), .B(n_818), .Y(n_975) );
OA21x2_ASAP7_75t_L g976 ( .A1(n_814), .A2(n_819), .B(n_809), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_877), .B(n_838), .Y(n_977) );
OA21x2_ASAP7_75t_L g978 ( .A1(n_814), .A2(n_819), .B(n_809), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_810), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_882), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g981 ( .A1(n_940), .A2(n_843), .B(n_837), .Y(n_981) );
AO21x2_ASAP7_75t_L g982 ( .A1(n_812), .A2(n_927), .B(n_869), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_904), .Y(n_983) );
AND2x4_ASAP7_75t_L g984 ( .A(n_903), .B(n_808), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_816), .B(n_815), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_886), .Y(n_986) );
AND2x4_ASAP7_75t_L g987 ( .A(n_941), .B(n_852), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_875), .Y(n_988) );
BUFx3_ASAP7_75t_L g989 ( .A(n_874), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_913), .B(n_958), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_835), .B(n_841), .Y(n_991) );
OAI21xp5_ASAP7_75t_L g992 ( .A1(n_959), .A2(n_812), .B(n_855), .Y(n_992) );
CKINVDCx5p33_ASAP7_75t_R g993 ( .A(n_826), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_870), .B(n_821), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_911), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_900), .Y(n_996) );
AO31x2_ASAP7_75t_L g997 ( .A1(n_836), .A2(n_949), .A3(n_859), .B(n_933), .Y(n_997) );
INVx2_ASAP7_75t_SL g998 ( .A(n_910), .Y(n_998) );
BUFx8_ASAP7_75t_L g999 ( .A(n_830), .Y(n_999) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_873), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_906), .A2(n_899), .B1(n_863), .B2(n_893), .Y(n_1001) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_848), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_900), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_906), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_879), .B(n_897), .Y(n_1005) );
OAI21x1_ASAP7_75t_SL g1006 ( .A1(n_846), .A2(n_927), .B(n_845), .Y(n_1006) );
A2O1A1Ixp33_ASAP7_75t_L g1007 ( .A1(n_924), .A2(n_851), .B(n_839), .C(n_923), .Y(n_1007) );
INVx3_ASAP7_75t_L g1008 ( .A(n_856), .Y(n_1008) );
INVx4_ASAP7_75t_L g1009 ( .A(n_873), .Y(n_1009) );
OAI21xp5_ASAP7_75t_L g1010 ( .A1(n_851), .A2(n_937), .B(n_895), .Y(n_1010) );
CKINVDCx11_ASAP7_75t_R g1011 ( .A(n_891), .Y(n_1011) );
CKINVDCx16_ASAP7_75t_R g1012 ( .A(n_891), .Y(n_1012) );
AOI21xp5_ASAP7_75t_L g1013 ( .A1(n_950), .A2(n_832), .B(n_937), .Y(n_1013) );
INVx1_ASAP7_75t_SL g1014 ( .A(n_914), .Y(n_1014) );
NOR2xp33_ASAP7_75t_L g1015 ( .A(n_948), .B(n_915), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_925), .B(n_954), .Y(n_1016) );
CKINVDCx5p33_ASAP7_75t_R g1017 ( .A(n_934), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_955), .B(n_894), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_847), .A2(n_919), .B1(n_945), .B2(n_840), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_827), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_947), .B(n_912), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_890), .B(n_849), .Y(n_1022) );
AO21x2_ASAP7_75t_L g1023 ( .A1(n_883), .A2(n_942), .B(n_931), .Y(n_1023) );
OA21x2_ASAP7_75t_L g1024 ( .A1(n_935), .A2(n_857), .B(n_946), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_860), .B(n_945), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_902), .Y(n_1026) );
OAI21xp5_ASAP7_75t_L g1027 ( .A1(n_876), .A2(n_884), .B(n_907), .Y(n_1027) );
OR2x6_ASAP7_75t_L g1028 ( .A(n_928), .B(n_887), .Y(n_1028) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_916), .A2(n_908), .B(n_858), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_811), .Y(n_1030) );
OR2x6_ASAP7_75t_L g1031 ( .A(n_928), .B(n_887), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_853), .B(n_820), .Y(n_1032) );
OAI21xp5_ASAP7_75t_L g1033 ( .A1(n_842), .A2(n_888), .B(n_871), .Y(n_1033) );
INVx1_ASAP7_75t_SL g1034 ( .A(n_917), .Y(n_1034) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_858), .A2(n_921), .B(n_922), .Y(n_1035) );
BUFx2_ASAP7_75t_L g1036 ( .A(n_929), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_824), .Y(n_1037) );
AO21x1_ASAP7_75t_L g1038 ( .A1(n_822), .A2(n_926), .B(n_920), .Y(n_1038) );
AND2x4_ASAP7_75t_L g1039 ( .A(n_932), .B(n_917), .Y(n_1039) );
A2O1A1Ixp33_ASAP7_75t_L g1040 ( .A1(n_881), .A2(n_938), .B(n_936), .C(n_813), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_854), .B(n_885), .Y(n_1041) );
AO31x2_ASAP7_75t_L g1042 ( .A1(n_896), .A2(n_898), .A3(n_861), .B(n_867), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_866), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g1044 ( .A1(n_864), .A2(n_944), .B(n_939), .Y(n_1044) );
NAND4xp25_ASAP7_75t_L g1045 ( .A(n_862), .B(n_868), .C(n_880), .D(n_866), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_854), .B(n_892), .Y(n_1046) );
AOI21xp33_ASAP7_75t_SL g1047 ( .A1(n_943), .A2(n_854), .B(n_831), .Y(n_1047) );
OAI22xp33_ASAP7_75t_SL g1048 ( .A1(n_831), .A2(n_901), .B1(n_892), .B2(n_885), .Y(n_1048) );
AO21x2_ASAP7_75t_L g1049 ( .A1(n_831), .A2(n_885), .B(n_892), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_909), .Y(n_1050) );
OAI21x1_ASAP7_75t_SL g1051 ( .A1(n_930), .A2(n_812), .B(n_900), .Y(n_1051) );
INVx2_ASAP7_75t_SL g1052 ( .A(n_930), .Y(n_1052) );
OR2x2_ASAP7_75t_L g1053 ( .A(n_956), .B(n_610), .Y(n_1053) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_817), .Y(n_1054) );
AO31x2_ASAP7_75t_L g1055 ( .A1(n_952), .A2(n_791), .A3(n_788), .B(n_836), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_956), .Y(n_1056) );
INVx1_ASAP7_75t_L g1057 ( .A(n_956), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_956), .B(n_953), .Y(n_1058) );
AO21x2_ASAP7_75t_L g1059 ( .A1(n_809), .A2(n_819), .B(n_814), .Y(n_1059) );
BUFx6f_ASAP7_75t_L g1060 ( .A(n_848), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_958), .A2(n_626), .B1(n_707), .B2(n_555), .Y(n_1061) );
OAI21xp5_ASAP7_75t_L g1062 ( .A1(n_952), .A2(n_809), .B(n_814), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_956), .Y(n_1063) );
NOR2xp33_ASAP7_75t_L g1064 ( .A(n_956), .B(n_807), .Y(n_1064) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_807), .B(n_956), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_956), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_956), .B(n_610), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_956), .Y(n_1068) );
AOI21xp5_ASAP7_75t_L g1069 ( .A1(n_952), .A2(n_729), .B(n_684), .Y(n_1069) );
OAI21xp33_ASAP7_75t_SL g1070 ( .A1(n_812), .A2(n_900), .B(n_819), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1071 ( .A(n_956), .B(n_610), .Y(n_1071) );
INVx3_ASAP7_75t_L g1072 ( .A(n_874), .Y(n_1072) );
AO21x2_ASAP7_75t_L g1073 ( .A1(n_809), .A2(n_819), .B(n_814), .Y(n_1073) );
A2O1A1Ixp33_ASAP7_75t_L g1074 ( .A1(n_959), .A2(n_918), .B(n_812), .C(n_681), .Y(n_1074) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_956), .Y(n_1075) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_913), .A2(n_610), .B1(n_626), .B2(n_590), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_807), .B(n_956), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_807), .B(n_956), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_956), .Y(n_1079) );
A2O1A1Ixp33_ASAP7_75t_L g1080 ( .A1(n_959), .A2(n_918), .B(n_812), .C(n_681), .Y(n_1080) );
AO21x2_ASAP7_75t_L g1081 ( .A1(n_809), .A2(n_819), .B(n_814), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_807), .Y(n_1082) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_956), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1084 ( .A(n_807), .B(n_956), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1077), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1082), .B(n_1004), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1077), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1078), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g1089 ( .A(n_1054), .Y(n_1089) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_1009), .Y(n_1090) );
OA21x2_ASAP7_75t_L g1091 ( .A1(n_1062), .A2(n_1010), .B(n_1029), .Y(n_1091) );
INVx3_ASAP7_75t_L g1092 ( .A(n_1002), .Y(n_1092) );
AO21x2_ASAP7_75t_L g1093 ( .A1(n_1047), .A2(n_1010), .B(n_1051), .Y(n_1093) );
OR2x6_ASAP7_75t_L g1094 ( .A(n_1009), .B(n_1000), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_971), .B(n_962), .Y(n_1095) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_962), .B(n_1078), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_969), .B(n_965), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1064), .B(n_1065), .Y(n_1098) );
OR2x2_ASAP7_75t_L g1099 ( .A(n_972), .B(n_973), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_989), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_1056), .Y(n_1101) );
AO21x2_ASAP7_75t_L g1102 ( .A1(n_1047), .A2(n_1062), .B(n_1006), .Y(n_1102) );
AO21x2_ASAP7_75t_L g1103 ( .A1(n_1069), .A2(n_1080), .B(n_1074), .Y(n_1103) );
INVx5_ASAP7_75t_L g1104 ( .A(n_1060), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1105 ( .A(n_1012), .B(n_969), .Y(n_1105) );
BUFx3_ASAP7_75t_L g1106 ( .A(n_966), .Y(n_1106) );
AO21x2_ASAP7_75t_L g1107 ( .A1(n_1013), .A2(n_1046), .B(n_1041), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1084), .B(n_1058), .Y(n_1108) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_1072), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_974), .B(n_1016), .Y(n_1110) );
BUFx2_ASAP7_75t_L g1111 ( .A(n_1014), .Y(n_1111) );
OA21x2_ASAP7_75t_L g1112 ( .A1(n_1030), .A2(n_1037), .B(n_1046), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_964), .Y(n_1113) );
AOI21x1_ASAP7_75t_L g1114 ( .A1(n_1028), .A2(n_1031), .B(n_1026), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_967), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1075), .B(n_1083), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1016), .B(n_975), .Y(n_1117) );
BUFx6f_ASAP7_75t_L g1118 ( .A(n_1052), .Y(n_1118) );
BUFx6f_ASAP7_75t_L g1119 ( .A(n_1039), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1049), .Y(n_1120) );
AND2x4_ASAP7_75t_L g1121 ( .A(n_1039), .B(n_1050), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_960), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1057), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1014), .B(n_1025), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_975), .B(n_979), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_980), .B(n_995), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1063), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1066), .Y(n_1128) );
AO21x2_ASAP7_75t_L g1129 ( .A1(n_982), .A2(n_1035), .B(n_992), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1068), .Y(n_1130) );
AOI22xp5_ASAP7_75t_L g1131 ( .A1(n_1076), .A2(n_1001), .B1(n_977), .B2(n_1015), .Y(n_1131) );
OR2x2_ASAP7_75t_L g1132 ( .A(n_1001), .B(n_1053), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_992), .B(n_1020), .Y(n_1133) );
INVx11_ASAP7_75t_L g1134 ( .A(n_999), .Y(n_1134) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1067), .B(n_1071), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_1079), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_986), .B(n_994), .Y(n_1137) );
OA21x2_ASAP7_75t_L g1138 ( .A1(n_968), .A2(n_1027), .B(n_1043), .Y(n_1138) );
INVx4_ASAP7_75t_L g1139 ( .A(n_1011), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_994), .B(n_988), .Y(n_1140) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_998), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1018), .B(n_1003), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_991), .B(n_1061), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_996), .B(n_1005), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1005), .B(n_1021), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g1146 ( .A(n_984), .Y(n_1146) );
AND2x4_ASAP7_75t_L g1147 ( .A(n_1008), .B(n_983), .Y(n_1147) );
BUFx2_ASAP7_75t_L g1148 ( .A(n_1034), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1055), .Y(n_1149) );
INVx3_ASAP7_75t_L g1150 ( .A(n_1028), .Y(n_1150) );
INVx2_ASAP7_75t_L g1151 ( .A(n_1055), .Y(n_1151) );
INVx3_ASAP7_75t_L g1152 ( .A(n_1031), .Y(n_1152) );
OA21x2_ASAP7_75t_L g1153 ( .A1(n_1027), .A2(n_1044), .B(n_981), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1019), .B(n_985), .Y(n_1154) );
OR2x6_ASAP7_75t_L g1155 ( .A(n_990), .B(n_978), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_987), .Y(n_1156) );
CKINVDCx5p33_ASAP7_75t_R g1157 ( .A(n_999), .Y(n_1157) );
OR2x6_ASAP7_75t_L g1158 ( .A(n_976), .B(n_978), .Y(n_1158) );
BUFx2_ASAP7_75t_L g1159 ( .A(n_1034), .Y(n_1159) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1021), .B(n_1081), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_1032), .A2(n_1038), .B1(n_1045), .B2(n_1073), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1036), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1059), .B(n_1081), .Y(n_1163) );
INVx4_ASAP7_75t_SL g1164 ( .A(n_1042), .Y(n_1164) );
OA21x2_ASAP7_75t_L g1165 ( .A1(n_1033), .A2(n_1007), .B(n_1040), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1022), .Y(n_1166) );
OR2x6_ASAP7_75t_L g1167 ( .A(n_961), .B(n_963), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_1045), .A2(n_1070), .B1(n_1017), .B2(n_993), .Y(n_1168) );
INVx3_ASAP7_75t_L g1169 ( .A(n_1042), .Y(n_1169) );
NOR2x1_ASAP7_75t_L g1170 ( .A(n_1090), .B(n_1023), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1096), .B(n_1070), .Y(n_1171) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1101), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1133), .B(n_997), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1133), .B(n_997), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1160), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1099), .B(n_997), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1160), .Y(n_1177) );
INVx2_ASAP7_75t_SL g1178 ( .A(n_1104), .Y(n_1178) );
INVx4_ASAP7_75t_L g1179 ( .A(n_1104), .Y(n_1179) );
INVx3_ASAP7_75t_L g1180 ( .A(n_1114), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1142), .B(n_1024), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1099), .Y(n_1182) );
CKINVDCx5p33_ASAP7_75t_R g1183 ( .A(n_1134), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1144), .B(n_1024), .Y(n_1184) );
BUFx3_ASAP7_75t_L g1185 ( .A(n_1090), .Y(n_1185) );
INVxp67_ASAP7_75t_SL g1186 ( .A(n_1111), .Y(n_1186) );
NOR2xp33_ASAP7_75t_L g1187 ( .A(n_1105), .B(n_970), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1144), .B(n_1048), .Y(n_1188) );
INVxp67_ASAP7_75t_SL g1189 ( .A(n_1111), .Y(n_1189) );
OAI21xp5_ASAP7_75t_L g1190 ( .A1(n_1131), .A2(n_1048), .B(n_1161), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1117), .B(n_1165), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1132), .B(n_1124), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1117), .B(n_1165), .Y(n_1193) );
BUFx2_ASAP7_75t_L g1194 ( .A(n_1148), .Y(n_1194) );
NOR2xp67_ASAP7_75t_L g1195 ( .A(n_1150), .B(n_1152), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1132), .B(n_1124), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1165), .B(n_1145), .Y(n_1197) );
INVx2_ASAP7_75t_SL g1198 ( .A(n_1104), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1112), .Y(n_1199) );
AOI22xp33_ASAP7_75t_SL g1200 ( .A1(n_1150), .A2(n_1152), .B1(n_1162), .B2(n_1146), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1145), .B(n_1097), .Y(n_1201) );
HB1xp67_ASAP7_75t_L g1202 ( .A(n_1136), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1110), .B(n_1155), .Y(n_1203) );
OR2x4_ASAP7_75t_L g1204 ( .A(n_1140), .B(n_1119), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1112), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1155), .B(n_1086), .Y(n_1206) );
AND2x4_ASAP7_75t_L g1207 ( .A(n_1164), .B(n_1155), .Y(n_1207) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1095), .B(n_1085), .Y(n_1208) );
BUFx3_ASAP7_75t_L g1209 ( .A(n_1104), .Y(n_1209) );
BUFx3_ASAP7_75t_L g1210 ( .A(n_1104), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1163), .B(n_1125), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1163), .B(n_1125), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1095), .B(n_1087), .Y(n_1213) );
BUFx2_ASAP7_75t_L g1214 ( .A(n_1159), .Y(n_1214) );
OR2x6_ASAP7_75t_L g1215 ( .A(n_1158), .B(n_1119), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1088), .B(n_1137), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1137), .B(n_1140), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_1154), .A2(n_1168), .B1(n_1098), .B2(n_1105), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1149), .B(n_1151), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1151), .B(n_1158), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1158), .B(n_1113), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1126), .B(n_1166), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1199), .Y(n_1223) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_1207), .B(n_1164), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1211), .B(n_1102), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1192), .B(n_1135), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1212), .B(n_1102), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1212), .B(n_1102), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1191), .B(n_1138), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1191), .B(n_1138), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1193), .B(n_1138), .Y(n_1231) );
NAND2x1_ASAP7_75t_L g1232 ( .A(n_1207), .B(n_1120), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_1202), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1193), .B(n_1169), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1192), .B(n_1135), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1171), .B(n_1126), .Y(n_1236) );
BUFx3_ASAP7_75t_L g1237 ( .A(n_1209), .Y(n_1237) );
INVx1_ASAP7_75t_SL g1238 ( .A(n_1185), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1197), .B(n_1169), .Y(n_1239) );
AND2x4_ASAP7_75t_SL g1240 ( .A(n_1179), .B(n_1119), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1205), .Y(n_1241) );
HB1xp67_ASAP7_75t_L g1242 ( .A(n_1172), .Y(n_1242) );
INVx1_ASAP7_75t_SL g1243 ( .A(n_1185), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1205), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_1175), .B(n_1115), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1188), .B(n_1153), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1188), .B(n_1129), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1196), .B(n_1129), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1173), .B(n_1107), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1174), .B(n_1107), .Y(n_1250) );
AOI21xp5_ASAP7_75t_L g1251 ( .A1(n_1170), .A2(n_1103), .B(n_1093), .Y(n_1251) );
OR2x2_ASAP7_75t_L g1252 ( .A(n_1177), .B(n_1116), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1174), .B(n_1091), .Y(n_1253) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_1204), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1203), .B(n_1091), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1203), .B(n_1103), .Y(n_1256) );
BUFx2_ASAP7_75t_L g1257 ( .A(n_1204), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1181), .B(n_1103), .Y(n_1258) );
NAND4xp25_ASAP7_75t_L g1259 ( .A(n_1218), .B(n_1139), .C(n_1108), .D(n_1143), .Y(n_1259) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_1194), .Y(n_1260) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1252), .B(n_1176), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1247), .B(n_1182), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1223), .Y(n_1263) );
OAI32xp33_ASAP7_75t_L g1264 ( .A1(n_1259), .A2(n_1139), .A3(n_1187), .B1(n_1089), .B2(n_1179), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1236), .B(n_1217), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1223), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1252), .B(n_1176), .Y(n_1267) );
NAND2x1p5_ASAP7_75t_L g1268 ( .A(n_1237), .B(n_1179), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1246), .B(n_1184), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1246), .B(n_1206), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1233), .B(n_1201), .Y(n_1271) );
AND2x4_ASAP7_75t_L g1272 ( .A(n_1224), .B(n_1234), .Y(n_1272) );
AOI22xp5_ASAP7_75t_SL g1273 ( .A1(n_1254), .A2(n_1157), .B1(n_1183), .B2(n_1139), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1241), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1255), .B(n_1221), .Y(n_1275) );
NAND3xp33_ASAP7_75t_L g1276 ( .A(n_1242), .B(n_1141), .C(n_1190), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1225), .B(n_1221), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1225), .B(n_1220), .Y(n_1278) );
INVx2_ASAP7_75t_SL g1279 ( .A(n_1237), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1227), .B(n_1220), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1241), .Y(n_1281) );
AND2x4_ASAP7_75t_SL g1282 ( .A(n_1224), .B(n_1215), .Y(n_1282) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1248), .B(n_1214), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1228), .B(n_1219), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1226), .B(n_1222), .Y(n_1285) );
BUFx3_ASAP7_75t_L g1286 ( .A(n_1240), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1253), .B(n_1219), .Y(n_1287) );
NAND2x1p5_ASAP7_75t_L g1288 ( .A(n_1254), .B(n_1209), .Y(n_1288) );
INVxp67_ASAP7_75t_SL g1289 ( .A(n_1260), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1244), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1244), .Y(n_1291) );
NOR2xp67_ASAP7_75t_L g1292 ( .A(n_1251), .B(n_1180), .Y(n_1292) );
NOR2xp33_ASAP7_75t_R g1293 ( .A(n_1286), .B(n_1157), .Y(n_1293) );
OR2x6_ASAP7_75t_L g1294 ( .A(n_1268), .B(n_1257), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1263), .Y(n_1295) );
NAND2xp33_ASAP7_75t_L g1296 ( .A(n_1268), .B(n_1089), .Y(n_1296) );
OAI21xp5_ASAP7_75t_L g1297 ( .A1(n_1276), .A2(n_1189), .B(n_1186), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1266), .Y(n_1298) );
NAND2xp5_ASAP7_75t_SL g1299 ( .A(n_1273), .B(n_1238), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1270), .B(n_1275), .Y(n_1300) );
AOI32xp33_ASAP7_75t_L g1301 ( .A1(n_1272), .A2(n_1243), .A3(n_1200), .B1(n_1256), .B2(n_1106), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1262), .B(n_1249), .Y(n_1302) );
NAND3xp33_ASAP7_75t_L g1303 ( .A(n_1289), .B(n_1123), .C(n_1122), .Y(n_1303) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1271), .B(n_1226), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1262), .B(n_1250), .Y(n_1305) );
NOR2xp33_ASAP7_75t_L g1306 ( .A(n_1285), .B(n_1235), .Y(n_1306) );
NOR2x1_ASAP7_75t_L g1307 ( .A(n_1286), .B(n_1106), .Y(n_1307) );
OR2x6_ASAP7_75t_L g1308 ( .A(n_1268), .B(n_1232), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1265), .B(n_1250), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1295), .Y(n_1310) );
NAND2xp5_ASAP7_75t_SL g1311 ( .A(n_1301), .B(n_1288), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1306), .B(n_1269), .Y(n_1312) );
A2O1A1Ixp33_ASAP7_75t_L g1313 ( .A1(n_1296), .A2(n_1264), .B(n_1282), .C(n_1286), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1300), .B(n_1269), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1298), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1309), .B(n_1284), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1302), .B(n_1284), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1305), .B(n_1277), .Y(n_1318) );
AOI21xp33_ASAP7_75t_SL g1319 ( .A1(n_1299), .A2(n_1288), .B(n_1279), .Y(n_1319) );
OAI21xp5_ASAP7_75t_L g1320 ( .A1(n_1307), .A2(n_1303), .B(n_1297), .Y(n_1320) );
NAND2xp33_ASAP7_75t_SL g1321 ( .A(n_1293), .B(n_1232), .Y(n_1321) );
OAI21xp5_ASAP7_75t_L g1322 ( .A1(n_1320), .A2(n_1294), .B(n_1308), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1314), .B(n_1278), .Y(n_1323) );
OAI221xp5_ASAP7_75t_L g1324 ( .A1(n_1321), .A2(n_1294), .B1(n_1308), .B2(n_1304), .C(n_1261), .Y(n_1324) );
OAI221xp5_ASAP7_75t_L g1325 ( .A1(n_1313), .A2(n_1308), .B1(n_1267), .B2(n_1292), .C(n_1283), .Y(n_1325) );
AOI21xp33_ASAP7_75t_L g1326 ( .A1(n_1311), .A2(n_1245), .B(n_1128), .Y(n_1326) );
OAI21xp5_ASAP7_75t_L g1327 ( .A1(n_1319), .A2(n_1195), .B(n_1178), .Y(n_1327) );
AOI222xp33_ASAP7_75t_L g1328 ( .A1(n_1312), .A2(n_1222), .B1(n_1130), .B2(n_1127), .C1(n_1280), .C2(n_1287), .Y(n_1328) );
AOI222xp33_ASAP7_75t_L g1329 ( .A1(n_1310), .A2(n_1229), .B1(n_1230), .B2(n_1231), .C1(n_1258), .C2(n_1239), .Y(n_1329) );
NAND4xp25_ASAP7_75t_L g1330 ( .A(n_1318), .B(n_1216), .C(n_1208), .D(n_1213), .Y(n_1330) );
AOI221xp5_ASAP7_75t_L g1331 ( .A1(n_1315), .A2(n_1291), .B1(n_1290), .B2(n_1281), .C(n_1274), .Y(n_1331) );
NAND3xp33_ASAP7_75t_L g1332 ( .A(n_1316), .B(n_1291), .C(n_1281), .Y(n_1332) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1317), .Y(n_1333) );
AOI211x1_ASAP7_75t_L g1334 ( .A1(n_1322), .A2(n_1326), .B(n_1324), .C(n_1325), .Y(n_1334) );
OAI311xp33_ASAP7_75t_L g1335 ( .A1(n_1328), .A2(n_1329), .A3(n_1330), .B1(n_1327), .C1(n_1331), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_1333), .B(n_1332), .Y(n_1336) );
NAND3xp33_ASAP7_75t_L g1337 ( .A(n_1334), .B(n_1100), .C(n_1109), .Y(n_1337) );
XNOR2x1_ASAP7_75t_L g1338 ( .A(n_1335), .B(n_1167), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1336), .B(n_1323), .Y(n_1339) );
OR2x6_ASAP7_75t_L g1340 ( .A(n_1337), .B(n_1167), .Y(n_1340) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1338), .Y(n_1341) );
NOR3x1_ASAP7_75t_L g1342 ( .A(n_1339), .B(n_1198), .C(n_1156), .Y(n_1342) );
CKINVDCx16_ASAP7_75t_R g1343 ( .A(n_1341), .Y(n_1343) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1342), .Y(n_1344) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_1343), .A2(n_1340), .B1(n_1180), .B2(n_1094), .Y(n_1345) );
OAI21xp33_ASAP7_75t_L g1346 ( .A1(n_1344), .A2(n_1340), .B(n_1209), .Y(n_1346) );
OAI21xp33_ASAP7_75t_L g1347 ( .A1(n_1346), .A2(n_1094), .B(n_1210), .Y(n_1347) );
NAND3xp33_ASAP7_75t_L g1348 ( .A(n_1347), .B(n_1345), .C(n_1118), .Y(n_1348) );
AOI21xp33_ASAP7_75t_SL g1349 ( .A1(n_1348), .A2(n_1147), .B(n_1180), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_1349), .A2(n_1180), .B1(n_1121), .B2(n_1214), .Y(n_1350) );
AOI21xp33_ASAP7_75t_SL g1351 ( .A1(n_1350), .A2(n_1121), .B(n_1092), .Y(n_1351) );
endmodule