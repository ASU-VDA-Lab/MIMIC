module fake_aes_8804_n_34 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
XNOR2xp5_ASAP7_75t_L g15 ( .A(n_6), .B(n_0), .Y(n_15) );
INVxp67_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_12), .B(n_11), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_7), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_10), .Y(n_19) );
NAND2xp33_ASAP7_75t_SL g20 ( .A(n_14), .B(n_1), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_16), .B(n_2), .Y(n_22) );
CKINVDCx6p67_ASAP7_75t_R g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVxp67_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
AOI211xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_20), .B(n_26), .C(n_15), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
NAND4xp25_ASAP7_75t_SL g31 ( .A(n_29), .B(n_17), .C(n_21), .D(n_19), .Y(n_31) );
HB1xp67_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_32), .Y(n_33) );
AOI322xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_31), .A3(n_4), .B1(n_5), .B2(n_8), .C1(n_9), .C2(n_13), .Y(n_34) );
endmodule