module fake_jpeg_3730_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_31),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_38),
.B1(n_19),
.B2(n_26),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_33),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_59),
.Y(n_82)
);

BUFx2_ASAP7_75t_SL g57 ( 
.A(n_36),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_22),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_18),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_14),
.B(n_13),
.C(n_16),
.Y(n_74)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_22),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_28),
.B1(n_19),
.B2(n_17),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_74),
.B1(n_83),
.B2(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_78),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_27),
.B(n_31),
.C(n_14),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_51),
.B1(n_34),
.B2(n_13),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_87),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

XNOR2x1_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_27),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_92),
.C(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_52),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_27),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_98),
.B1(n_80),
.B2(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_34),
.B1(n_47),
.B2(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_80),
.B1(n_68),
.B2(n_84),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_65),
.B(n_60),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_99),
.Y(n_110)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_70),
.B(n_9),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_108),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_94),
.C(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_109),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_84),
.C(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_93),
.B1(n_86),
.B2(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_100),
.Y(n_116)
);

OA21x2_ASAP7_75t_SL g119 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_79),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_117),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_124),
.C(n_104),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_109),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_126),
.C(n_13),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_112),
.C(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_103),
.B(n_108),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_129),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_72),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_121),
.B1(n_124),
.B2(n_72),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_16),
.B1(n_8),
.B2(n_3),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_0),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_133),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_4),
.B(n_5),
.C(n_10),
.D(n_12),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_136),
.B(n_4),
.C(n_5),
.Y(n_137)
);

NOR2x1p5_ASAP7_75t_SL g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_132),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_140),
.B(n_135),
.CI(n_2),
.CON(n_141),
.SN(n_141)
);


endmodule