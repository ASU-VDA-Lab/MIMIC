module real_jpeg_4714_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_2),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_2),
.A2(n_47),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_2),
.A2(n_47),
.B1(n_117),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_2),
.A2(n_47),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_2),
.B(n_150),
.C(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_2),
.B(n_249),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_2),
.A2(n_256),
.B(n_258),
.C(n_259),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_2),
.B(n_269),
.C(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_2),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_2),
.B(n_215),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_2),
.B(n_26),
.Y(n_295)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_4),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_4),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_4),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_5),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_13)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_6),
.Y(n_238)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_9),
.Y(n_130)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_9),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_10),
.A2(n_51),
.B1(n_55),
.B2(n_58),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_43),
.B1(n_58),
.B2(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_10),
.A2(n_58),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_10),
.A2(n_58),
.B1(n_76),
.B2(n_188),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_11),
.A2(n_85),
.B1(n_89),
.B2(n_92),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_92),
.B1(n_116),
.B2(n_119),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_92),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_11),
.A2(n_92),
.B1(n_163),
.B2(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_12),
.Y(n_114)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_366),
.B(n_368),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_138),
.B(n_365),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_133),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_22),
.B(n_133),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_121),
.C(n_132),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_23),
.A2(n_24),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_49),
.C(n_93),
.Y(n_24)
);

XNOR2x1_ASAP7_75t_L g145 ( 
.A(n_25),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_25),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_203),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_25),
.A2(n_180),
.B1(n_181),
.B2(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_25),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_25),
.A2(n_222),
.B1(n_252),
.B2(n_262),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_25),
.B(n_172),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_25),
.A2(n_222),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_25),
.A2(n_180),
.B(n_218),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_25),
.A2(n_222),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_25),
.A2(n_222),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

OA21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B(n_45),
.Y(n_25)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_26),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_32),
.Y(n_149)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_37)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_38),
.Y(n_135)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_47),
.A2(n_73),
.B(n_76),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_49),
.A2(n_93),
.B1(n_94),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_49),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_59),
.B1(n_72),
.B2(n_84),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_50),
.A2(n_59),
.B1(n_72),
.B2(n_147),
.Y(n_343)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_72),
.B(n_84),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AO21x2_ASAP7_75t_SL g146 ( 
.A1(n_60),
.A2(n_72),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_61)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_62),
.Y(n_257)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_72),
.Y(n_249)
);

OA22x2_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_78),
.B2(n_81),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_91),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_93),
.A2(n_94),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_94),
.B(n_222),
.C(n_343),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_104),
.B(n_115),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_95),
.B(n_104),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_95),
.A2(n_104),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

NAND2x1_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_104),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_103),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_99),
.Y(n_270)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_110),
.B2(n_114),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_105),
.B(n_279),
.Y(n_278)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_115),
.Y(n_214)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g271 ( 
.A(n_118),
.Y(n_271)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_121),
.B(n_132),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_131),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_124),
.B1(n_131),
.B2(n_134),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g367 ( 
.A1(n_123),
.A2(n_131),
.B(n_134),
.Y(n_367)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_133),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_133),
.B(n_367),
.Y(n_369)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_359),
.B(n_364),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_337),
.B(n_356),
.Y(n_139)
);

OAI211xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_242),
.B(n_331),
.C(n_336),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_224),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_142),
.A2(n_224),
.B(n_332),
.C(n_335),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_206),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_143),
.B(n_206),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_179),
.C(n_191),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_144),
.B(n_179),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_151),
.B1(n_177),
.B2(n_178),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_145),
.B(n_192),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_145),
.A2(n_177),
.B1(n_231),
.B2(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_146),
.B(n_212),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_146),
.A2(n_205),
.B(n_222),
.C(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_146),
.A2(n_172),
.B1(n_203),
.B2(n_228),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_146),
.A2(n_203),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_151),
.A2(n_202),
.B(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_172),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_152),
.A2(n_172),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_159),
.B1(n_165),
.B2(n_169),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_157),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_159),
.B1(n_194),
.B2(n_200),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_155),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_169),
.B(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_172),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_172),
.A2(n_228),
.B1(n_248),
.B2(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_172),
.A2(n_228),
.B1(n_266),
.B2(n_267),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_172),
.A2(n_228),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_172),
.A2(n_203),
.B(n_254),
.C(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_172),
.B(n_203),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_172),
.A2(n_193),
.B1(n_228),
.B2(n_322),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_190),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_184),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_195),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_187),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_212)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_202),
.B(n_204),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_193),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_203),
.A2(n_211),
.B(n_216),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_203),
.B(n_239),
.C(n_294),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AND3x1_ASAP7_75t_L g324 ( 
.A(n_205),
.B(n_301),
.C(n_325),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_223),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_210),
.B(n_217),
.C(n_223),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

FAx1_ASAP7_75t_L g339 ( 
.A(n_216),
.B(n_340),
.CI(n_345),
.CON(n_339),
.SN(n_339)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_222),
.B(n_351),
.C(n_355),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_240),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_225),
.B(n_240),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.C(n_230),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_226),
.B(n_227),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_248),
.C(n_250),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_228),
.B(n_291),
.C(n_298),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_230),
.B(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_231),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_232),
.A2(n_233),
.B1(n_239),
.B2(n_250),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_239),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_250),
.B1(n_255),
.B2(n_261),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_239),
.A2(n_250),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_239),
.B(n_255),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_313),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_303),
.B(n_312),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_289),
.B(n_302),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_263),
.B(n_288),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_250),
.B(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_262),
.Y(n_251)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_275),
.B(n_287),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_272),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_285),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_283),
.Y(n_276)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_299),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_299),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_305),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_309),
.C(n_310),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_316),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_323),
.B2(n_324),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_323),
.C(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_326),
.A2(n_333),
.B(n_334),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_329),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_347),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_346),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_339),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_346),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_348),
.Y(n_358)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_343),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_347),
.A2(n_357),
.B(n_358),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_355),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_363),
.Y(n_364)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_369),
.Y(n_368)
);


endmodule