module real_jpeg_2416_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_1),
.A2(n_42),
.B1(n_48),
.B2(n_64),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_1),
.A2(n_44),
.B1(n_55),
.B2(n_64),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_1),
.A2(n_64),
.B1(n_71),
.B2(n_73),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_1),
.A2(n_28),
.B1(n_36),
.B2(n_64),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_42),
.B1(n_48),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_71),
.B1(n_73),
.B2(n_77),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_3),
.A2(n_28),
.B1(n_36),
.B2(n_77),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_4),
.A2(n_44),
.B1(n_55),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_42),
.B1(n_48),
.B2(n_60),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_60),
.B1(n_71),
.B2(n_73),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_4),
.A2(n_28),
.B1(n_36),
.B2(n_60),
.Y(n_206)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_11),
.A2(n_71),
.B1(n_73),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_11),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_11),
.A2(n_28),
.B1(n_36),
.B2(n_91),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_11),
.A2(n_42),
.B1(n_48),
.B2(n_91),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_12),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_12),
.A2(n_37),
.B1(n_71),
.B2(n_73),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_13),
.A2(n_44),
.B1(n_55),
.B2(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_42),
.B1(n_48),
.B2(n_58),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_13),
.A2(n_58),
.B1(n_71),
.B2(n_73),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_13),
.A2(n_28),
.B1(n_36),
.B2(n_58),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_14),
.A2(n_55),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_14),
.B(n_48),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_28),
.C(n_85),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_14),
.A2(n_46),
.B1(n_71),
.B2(n_73),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_14),
.B(n_78),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_14),
.B(n_32),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_14),
.B(n_92),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g222 ( 
.A1(n_14),
.A2(n_48),
.B(n_171),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_28),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_15),
.A2(n_39),
.B1(n_71),
.B2(n_73),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_20),
.B(n_111),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.C(n_101),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_21),
.A2(n_22),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_50),
.B2(n_51),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_52),
.C(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_25),
.A2(n_26),
.B1(n_40),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_38),
.Y(n_26)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_27),
.B(n_106),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_27),
.A2(n_117),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_27),
.A2(n_32),
.B1(n_46),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_27),
.A2(n_32),
.B1(n_203),
.B2(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_28),
.A2(n_36),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_28),
.B(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_31),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_31),
.A2(n_35),
.B(n_120),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_31),
.A2(n_103),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_32),
.B(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_38),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_40),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.C(n_47),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_44),
.B1(n_49),
.B2(n_55),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_56)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_48),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_42),
.B(n_69),
.C(n_73),
.Y(n_172)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_48),
.C(n_49),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_61),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_56),
.B1(n_57),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_53),
.A2(n_56),
.B1(n_59),
.B2(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_56),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B(n_74),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_78),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_65),
.A2(n_76),
.B(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_65),
.A2(n_70),
.B1(n_99),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_65),
.A2(n_70),
.B1(n_152),
.B2(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_67),
.A2(n_71),
.B(n_170),
.C(n_172),
.Y(n_169)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_73),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_71),
.B(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_78),
.B(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_79),
.A2(n_80),
.B1(n_101),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_93),
.C(n_96),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_81),
.A2(n_96),
.B1(n_97),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_88),
.B(n_89),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_108),
.B1(n_109),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_82),
.A2(n_108),
.B1(n_166),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_90),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_83),
.A2(n_165),
.B(n_167),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_83),
.A2(n_92),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_83),
.A2(n_92),
.B1(n_189),
.B2(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_87),
.B(n_88),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_107),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_103),
.A2(n_105),
.B(n_118),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B(n_110),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_121),
.B2(n_122),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_132),
.B2(n_133),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_157),
.B(n_232),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_153),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_138),
.B(n_153),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_145),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_140),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_145),
.B1(n_146),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.C(n_151),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_178),
.B(n_231),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_174),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_160),
.B(n_174),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_168),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_161),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_164),
.B(n_168),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_173),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_226),
.B(n_230),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_216),
.B(n_225),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_197),
.B(n_215),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_194),
.C(n_196),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_209),
.B(n_214),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_204),
.B(n_208),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_207),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_213),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_221),
.C(n_223),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_229),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);


endmodule