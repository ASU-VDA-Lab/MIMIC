module real_jpeg_12744_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_357, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_357;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_2),
.B(n_67),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_2),
.B(n_81),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_2),
.B(n_62),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_2),
.B(n_45),
.Y(n_295)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_5),
.B(n_81),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_5),
.B(n_53),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_5),
.B(n_62),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_5),
.B(n_31),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_6),
.B(n_27),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_6),
.B(n_62),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_6),
.B(n_67),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_81),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_6),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_6),
.B(n_45),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_6),
.B(n_31),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_6),
.B(n_35),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_7),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_7),
.B(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_7),
.B(n_45),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_7),
.B(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_7),
.B(n_27),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_7),
.B(n_62),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_10),
.B(n_62),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_10),
.B(n_45),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_10),
.B(n_27),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_10),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_10),
.B(n_31),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_12),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_12),
.B(n_62),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_12),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_12),
.B(n_31),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_12),
.B(n_53),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_12),
.B(n_67),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_13),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_13),
.B(n_45),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_13),
.B(n_67),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_14),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_14),
.B(n_31),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_14),
.B(n_27),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_53),
.Y(n_185)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_147),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_20),
.B(n_121),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_107),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_21),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_64),
.C(n_76),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_22),
.A2(n_23),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_24),
.B(n_41),
.C(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_26),
.B(n_30),
.C(n_33),
.Y(n_106)
);

INVx5_ASAP7_75t_SL g173 ( 
.A(n_27),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_34),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_34),
.B(n_49),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_34),
.B(n_204),
.Y(n_275)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_37),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_37),
.B(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_57),
.B2(n_58),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_56),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_44),
.B(n_52),
.C(n_54),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_48),
.A2(n_54),
.B1(n_140),
.B2(n_141),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_SL g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_50),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_50),
.B(n_91),
.Y(n_293)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_66),
.C(n_70),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_55),
.B1(n_66),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_52),
.A2(n_55),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_52),
.B(n_165),
.Y(n_181)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_53),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_54),
.B(n_140),
.C(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_59),
.A2(n_61),
.B1(n_137),
.B2(n_315),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_59),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_60),
.B(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_61),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_64),
.B(n_76),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_72),
.C(n_74),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_66),
.A2(n_79),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_66),
.B(n_232),
.Y(n_264)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_68),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_68),
.B(n_204),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_74),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_74),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_117),
.C(n_119),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_73),
.B(n_99),
.C(n_103),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_73),
.A2(n_74),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_74),
.B(n_185),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.C(n_82),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_77),
.B(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_80),
.A2(n_82),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_80),
.Y(n_326)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_82),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_83),
.B(n_107),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_95),
.B2(n_96),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_97),
.C(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_94),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_89),
.C(n_92),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_90),
.B(n_161),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_93),
.B(n_163),
.Y(n_271)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_105),
.B2(n_106),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_99),
.A2(n_104),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_99),
.B(n_287),
.C(n_288),
.Y(n_317)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_102),
.A2(n_103),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_102),
.A2(n_103),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_103),
.B(n_225),
.C(n_227),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_112),
.C(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_120),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_119),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_121),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.CI(n_145),
.CON(n_121),
.SN(n_121)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_135),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

AOI321xp33_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_333),
.A3(n_343),
.B1(n_347),
.B2(n_352),
.C(n_357),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_278),
.C(n_328),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_249),
.B(n_277),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_219),
.B(n_248),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_188),
.B(n_218),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_167),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_153),
.B(n_167),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.C(n_164),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_170),
.B1(n_171),
.B2(n_179),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_215),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.CI(n_157),
.CON(n_154),
.SN(n_154)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_162),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_163),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_180),
.B2(n_187),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_179),
.C(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_175),
.C(n_178),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_181),
.B(n_183),
.C(n_184),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_185),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_185),
.A2(n_186),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_185),
.B(n_301),
.C(n_304),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_212),
.B(n_217),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_201),
.B(n_211),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_191),
.B(n_196),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_199),
.C(n_200),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_206),
.B(n_210),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_220),
.B(n_221),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_234),
.B2(n_235),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_236),
.C(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_230),
.C(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_246),
.B2(n_247),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_245),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_242),
.C(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_241),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_251),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_267),
.B2(n_276),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_266),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_254),
.B(n_266),
.C(n_276),
.Y(n_329)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_262),
.B2(n_263),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_264),
.C(n_265),
.Y(n_297)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_258),
.Y(n_353)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.CI(n_261),
.CON(n_258),
.SN(n_258)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_306)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_267),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.CI(n_273),
.CON(n_267),
.SN(n_267)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_268),
.B(n_269),
.C(n_273),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B(n_272),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_272),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_272),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g348 ( 
.A1(n_279),
.A2(n_349),
.B(n_350),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_310),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_280),
.B(n_310),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_298),
.C(n_309),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_297),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_290),
.C(n_297),
.Y(n_327)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_286),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_287),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_294),
.C(n_296),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_298),
.A2(n_299),
.B1(n_309),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_306),
.C(n_308),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_309),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_327),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_319),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_319),
.C(n_327),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_317),
.C(n_318),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_322),
.C(n_323),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_330),
.Y(n_349)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_334),
.A2(n_348),
.B(n_351),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_335),
.B(n_336),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_339),
.C(n_342),
.Y(n_344)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_345),
.Y(n_352)
);


endmodule