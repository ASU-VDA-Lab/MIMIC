module real_jpeg_30499_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_366;
wire n_149;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_0),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g458 ( 
.A(n_0),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_1),
.A2(n_42),
.B1(n_44),
.B2(n_48),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_1),
.A2(n_48),
.B1(n_87),
.B2(n_269),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_2),
.A2(n_30),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_3),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_3),
.A2(n_136),
.B1(n_219),
.B2(n_223),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_3),
.A2(n_136),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_3),
.A2(n_136),
.B1(n_502),
.B2(n_506),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_4),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_4),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_4),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_5),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_5),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_6),
.Y(n_420)
);

AOI22x1_ASAP7_75t_SL g121 ( 
.A1(n_7),
.A2(n_122),
.B1(n_125),
.B2(n_130),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_7),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_7),
.A2(n_130),
.B1(n_318),
.B2(n_320),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_7),
.A2(n_87),
.B1(n_130),
.B2(n_431),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_7),
.A2(n_130),
.B1(n_446),
.B2(n_448),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_8),
.A2(n_183),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_8),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_8),
.A2(n_230),
.B1(n_349),
.B2(n_352),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_8),
.A2(n_230),
.B1(n_392),
.B2(n_395),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_8),
.A2(n_230),
.B1(n_440),
.B2(n_444),
.Y(n_439)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_9),
.A2(n_252),
.B1(n_255),
.B2(n_258),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_9),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_10),
.A2(n_76),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_10),
.A2(n_81),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_10),
.A2(n_81),
.B1(n_362),
.B2(n_366),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_11),
.B(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_11),
.A2(n_201),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_11),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_11),
.B(n_173),
.Y(n_427)
);

OAI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_11),
.A2(n_35),
.B1(n_439),
.B2(n_457),
.Y(n_456)
);

OAI32xp33_ASAP7_75t_L g476 ( 
.A1(n_11),
.A2(n_143),
.A3(n_477),
.B1(n_481),
.B2(n_485),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_11),
.A2(n_370),
.B1(n_498),
.B2(n_499),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_12),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_14),
.Y(n_405)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_15),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_15),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_15),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_15),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_16),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_16),
.A2(n_90),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_16),
.A2(n_90),
.B1(n_292),
.B2(n_295),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_17),
.A2(n_164),
.B1(n_169),
.B2(n_170),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_17),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_17),
.A2(n_169),
.B1(n_284),
.B2(n_287),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_17),
.A2(n_169),
.B1(n_332),
.B2(n_335),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_17),
.A2(n_169),
.B1(n_208),
.B2(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_303),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_300),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_259),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_22),
.B(n_259),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_180),
.C(n_235),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2x1_ASAP7_75t_L g340 ( 
.A(n_24),
.B(n_235),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_94),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_25),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_53),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_26),
.B(n_53),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_35),
.B1(n_41),
.B2(n_49),
.Y(n_26)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_27),
.Y(n_212)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_29),
.Y(n_208)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_29),
.Y(n_368)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_34),
.Y(n_443)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_35),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_35),
.A2(n_41),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_35),
.B(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_35),
.A2(n_439),
.B1(n_445),
.B2(n_452),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_38),
.Y(n_360)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_40),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_46),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_47),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_47),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_47),
.Y(n_365)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_47),
.Y(n_451)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_50),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_464)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_75),
.B1(n_85),
.B2(n_86),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_54),
.A2(n_85),
.B1(n_86),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_54),
.A2(n_85),
.B1(n_237),
.B2(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_54),
.A2(n_75),
.B1(n_85),
.B2(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_54),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_54),
.A2(n_85),
.B1(n_429),
.B2(n_430),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_54),
.A2(n_523),
.B(n_524),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_62),
.B(n_69),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_61),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_61),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_61),
.Y(n_432)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_61),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_62),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_63),
.Y(n_241)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g505 ( 
.A(n_65),
.Y(n_505)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_70),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_70),
.Y(n_425)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_74),
.Y(n_210)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_80),
.Y(n_244)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_85),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_85),
.B(n_370),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_89),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_93),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_140),
.B1(n_141),
.B2(n_179),
.Y(n_94)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_95),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_121),
.B1(n_131),
.B2(n_132),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_97),
.A2(n_228),
.B1(n_233),
.B2(n_234),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_97),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_280)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_97),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_110),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_106),
.B2(n_108),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_102),
.Y(n_286)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_106),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_117),
.B2(n_120),
.Y(n_110)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_112),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_113),
.Y(n_351)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_119),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_119),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_119),
.Y(n_356)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_121),
.Y(n_233)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_128),
.Y(n_287)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_131),
.Y(n_234)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_131),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_131),
.A2(n_229),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

NOR2x1_ASAP7_75t_R g369 ( 
.A(n_131),
.B(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_132),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_140),
.Y(n_263)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22x1_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_163),
.B1(n_172),
.B2(n_174),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_142),
.A2(n_163),
.B1(n_172),
.B2(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_142),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_142),
.A2(n_172),
.B1(n_218),
.B2(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_142),
.A2(n_172),
.B1(n_317),
.B2(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_142),
.A2(n_172),
.B1(n_348),
.B2(n_497),
.Y(n_496)
);

AO21x2_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_150),
.B(n_155),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_161),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_157),
.Y(n_395)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22x1_ASAP7_75t_L g288 ( 
.A1(n_173),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_174),
.Y(n_290)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_179),
.Y(n_262)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_180),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_215),
.C(n_226),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_181),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_205),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_182),
.A2(n_205),
.B1(n_206),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_182),
.Y(n_372)
);

OAI32xp33_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_185),
.A3(n_186),
.B1(n_191),
.B2(n_200),
.Y(n_182)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_SL g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_207),
.A2(n_211),
.B1(n_359),
.B2(n_361),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_210),
.Y(n_401)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_211),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_211),
.A2(n_361),
.B1(n_424),
.B2(n_490),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_217),
.B(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_222),
.Y(n_319)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_222),
.Y(n_480)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_227),
.Y(n_310)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_231),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2x2_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_245),
.Y(n_278)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_244),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

INVx3_ASAP7_75t_SL g276 ( 
.A(n_247),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_250),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_250),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_250),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_256),
.Y(n_444)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_277),
.Y(n_264)
);

XNOR2x2_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.Y(n_279)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_292),
.Y(n_498)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_295),
.Y(n_499)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_375),
.B(n_537),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_341),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_338),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_307),
.B(n_338),
.C(n_539),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_308),
.B(n_374),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_314),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_324),
.C(n_329),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_330),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_331),
.Y(n_525)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_334),
.Y(n_488)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_334),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_373),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_343),
.B(n_373),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_346),
.C(n_371),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_344),
.B(n_534),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_346),
.B(n_371),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_357),
.C(n_369),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_347),
.B(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_357),
.A2(n_358),
.B1(n_369),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_369),
.Y(n_519)
);

OAI21xp33_ASAP7_75t_SL g384 ( 
.A1(n_370),
.A2(n_385),
.B(n_387),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_388),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_370),
.B(n_452),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_370),
.B(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

AOI21x1_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_532),
.B(n_536),
.Y(n_376)
);

OAI21x1_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_515),
.B(n_531),
.Y(n_377)
);

AOI21x1_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_472),
.B(n_514),
.Y(n_378)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_435),
.B(n_471),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_411),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_381),
.B(n_411),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_397),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_382),
.A2(n_383),
.B1(n_397),
.B2(n_398),
.Y(n_463)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_390),
.B1(n_391),
.B2(n_396),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_387),
.Y(n_406)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_390),
.A2(n_396),
.B1(n_501),
.B2(n_511),
.Y(n_500)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_396),
.B(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_406),
.B1(n_407),
.B2(n_410),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_426),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_412),
.B(n_428),
.C(n_433),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_414),
.B1(n_421),
.B2(n_423),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_413),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_433),
.B2(n_434),
.Y(n_426)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_427),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_428),
.Y(n_434)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_430),
.Y(n_511)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI31xp33_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_462),
.A3(n_468),
.B(n_470),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_455),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_454),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_438),
.B(n_454),
.Y(n_469)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_444),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_445),
.Y(n_465)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx8_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

INVx8_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_464),
.Y(n_470)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_SL g514 ( 
.A(n_473),
.B(n_474),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_495),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_475),
.B(n_500),
.C(n_513),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_489),
.B1(n_493),
.B2(n_494),
.Y(n_475)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_476),
.B(n_494),
.Y(n_521)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_489),
.Y(n_494)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_500),
.B1(n_512),
.B2(n_513),
.Y(n_495)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_496),
.Y(n_513)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_501),
.Y(n_523)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_530),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_530),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_520),
.B1(n_528),
.B2(n_529),
.Y(n_516)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_517),
.Y(n_529)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_520),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_521),
.A2(n_522),
.B1(n_526),
.B2(n_527),
.Y(n_520)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_521),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_522),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_526),
.C(n_529),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_533),
.B(n_535),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_535),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);


endmodule