module real_jpeg_14329_n_17 (n_329, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_329;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_286;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_1),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_1),
.A2(n_35),
.B1(n_53),
.B2(n_54),
.Y(n_323)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_4),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_159),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_159),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_159),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_6),
.A2(n_39),
.B1(n_57),
.B2(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_6),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_9),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_9),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_77),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_77),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_77),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g248 ( 
.A(n_11),
.B(n_58),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_12),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_30),
.C(n_44),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_12),
.B(n_75),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_12),
.A2(n_110),
.B(n_163),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_57),
.B(n_74),
.C(n_190),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_147),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_12),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_12),
.B(n_53),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_13),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_55),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_66),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_66),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_66),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_15),
.A2(n_53),
.B1(n_54),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_15),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_119),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_119),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_119),
.Y(n_238)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_320),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_307),
.B(n_319),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_135),
.B(n_304),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_122),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_97),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_22),
.B(n_97),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_67),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_68),
.C(n_83),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B(n_51),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_24),
.A2(n_25),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_26),
.A2(n_27),
.B1(n_51),
.B2(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_26),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_33),
.Y(n_27)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_28),
.A2(n_32),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_28),
.B(n_164),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_28),
.A2(n_32),
.B1(n_109),
.B2(n_252),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_29),
.B(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_32),
.B(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_34),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_47),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_38),
.A2(n_42),
.B1(n_50),
.B2(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_41),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_40),
.B(n_151),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_41),
.A2(n_73),
.B(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_42),
.A2(n_50),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_42),
.B(n_149),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_42),
.A2(n_50),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_42),
.A2(n_50),
.B1(n_114),
.B2(n_241),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_48),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_46),
.A2(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_46),
.B(n_147),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_46),
.A2(n_160),
.B(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_50),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_60),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_56),
.B1(n_62),
.B2(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_54),
.A2(n_62),
.B(n_147),
.C(n_234),
.Y(n_233)
);

AOI32xp33_ASAP7_75t_L g247 ( 
.A1(n_54),
.A2(n_57),
.A3(n_59),
.B1(n_235),
.B2(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_65),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_56),
.A2(n_62),
.B1(n_95),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_56),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_56),
.A2(n_60),
.B(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_56),
.A2(n_62),
.B1(n_118),
.B2(n_262),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_58),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_61),
.A2(n_215),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_61),
.A2(n_215),
.B1(n_314),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_62),
.A2(n_118),
.B(n_120),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_83),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_69),
.B(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_80),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_78),
.B1(n_88),
.B2(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_70),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_70),
.A2(n_78),
.B1(n_210),
.B2(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_70),
.A2(n_196),
.B(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_75),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_71),
.B(n_197),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_71),
.A2(n_75),
.B(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_75),
.B(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_78),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_78),
.A2(n_116),
.B(n_211),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_81),
.A2(n_146),
.B(n_148),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_81),
.A2(n_148),
.B(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_85),
.B(n_90),
.C(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_90),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_90),
.B(n_127),
.C(n_131),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_94),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_94),
.B(n_126),
.C(n_133),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.C(n_104),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_103),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_104),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.C(n_117),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_105),
.A2(n_106),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_107),
.A2(n_112),
.B1(n_113),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_107),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_110),
.A2(n_111),
.B1(n_192),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_110),
.A2(n_111),
.B1(n_218),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_111),
.A2(n_169),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_111),
.B(n_147),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_111),
.A2(n_177),
.B(n_192),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_115),
.B(n_117),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_121),
.B(n_233),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_122),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_134),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_123),
.B(n_134),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_133),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_128),
.Y(n_313)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_132),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_298),
.B(n_303),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_286),
.B(n_297),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_254),
.A3(n_279),
.B1(n_284),
.B2(n_285),
.C(n_329),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_227),
.B(n_253),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_204),
.B(n_226),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_185),
.B(n_203),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_165),
.B(n_184),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_143),
.B(n_152),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_145),
.B1(n_150),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_161),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_157),
.C(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_162),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_173),
.B(n_183),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_167),
.B(n_171),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_178),
.B(n_182),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_176),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_186),
.B(n_187),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_198),
.C(n_202),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_191),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_205),
.B(n_206),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_219),
.B2(n_220),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_222),
.C(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_213),
.C(n_217),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_229),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_243),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_230),
.B(n_244),
.C(n_245),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_236),
.B2(n_242),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_237),
.C(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_250),
.Y(n_264)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_269),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_269),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.C(n_268),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_257),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_264),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_263),
.C(n_264),
.Y(n_278)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_265),
.B(n_268),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_267),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_278),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_273),
.C(n_278),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_276),
.C(n_277),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_296),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_291),
.C(n_292),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_318),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_318),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_317),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_312),
.B1(n_315),
.B2(n_316),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_315),
.C(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_322),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_324),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);


endmodule