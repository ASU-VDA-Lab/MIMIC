module fake_jpeg_2378_n_118 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_49),
.B1(n_45),
.B2(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_59),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_42),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_41),
.B1(n_37),
.B2(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_37),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_46),
.B1(n_49),
.B2(n_40),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_57),
.B1(n_39),
.B2(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_69),
.B(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_48),
.B1(n_1),
.B2(n_2),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_54),
.B1(n_36),
.B2(n_50),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_38),
.Y(n_82)
);

NOR4xp25_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_50),
.C(n_1),
.D(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_61),
.B1(n_71),
.B2(n_58),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_70),
.C(n_58),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_77),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_91),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_76),
.C(n_3),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_97),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_98),
.C(n_15),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_102),
.B1(n_86),
.B2(n_93),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_0),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_9),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_83),
.B(n_81),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_107),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_110),
.B1(n_107),
.B2(n_104),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_108),
.C(n_103),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_113),
.A3(n_98),
.B1(n_16),
.B2(n_96),
.C1(n_10),
.C2(n_13),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_14),
.Y(n_116)
);

OA21x2_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_11),
.B(n_12),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_14),
.Y(n_118)
);


endmodule