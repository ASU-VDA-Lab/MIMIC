module fake_jpeg_18180_n_204 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_0),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_12),
.B(n_22),
.C(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_30),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_20),
.C(n_17),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_27),
.C(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_28),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_27),
.B1(n_28),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_52),
.B1(n_25),
.B2(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_55),
.Y(n_67)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_54),
.Y(n_59)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_28),
.B1(n_25),
.B2(n_29),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_30),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_30),
.B(n_22),
.C(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_15),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_18),
.B(n_15),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_13),
.B(n_14),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_25),
.B1(n_33),
.B2(n_34),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_56),
.B1(n_45),
.B2(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_14),
.Y(n_72)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_25),
.B(n_29),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_52),
.B1(n_26),
.B2(n_29),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_51),
.B1(n_41),
.B2(n_29),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_86),
.B1(n_49),
.B2(n_61),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_80),
.B1(n_85),
.B2(n_69),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_84),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_50),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_85),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_62),
.C(n_22),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_13),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_55),
.B1(n_37),
.B2(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_49),
.B1(n_44),
.B2(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_88),
.B(n_89),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_14),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_69),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NAND4xp25_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_53),
.C(n_70),
.D(n_44),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_66),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_110),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_66),
.B(n_59),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_61),
.B(n_74),
.Y(n_121)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_59),
.B1(n_71),
.B2(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_104),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_65),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_60),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_74),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_78),
.B1(n_57),
.B2(n_60),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_114),
.B1(n_116),
.B2(n_129),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_90),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_119),
.C(n_21),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_97),
.B1(n_109),
.B2(n_105),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_78),
.B1(n_74),
.B2(n_73),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_74),
.C(n_65),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_24),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_116),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_70),
.B(n_1),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_103),
.B1(n_101),
.B2(n_95),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_101),
.B1(n_93),
.B2(n_91),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_40),
.Y(n_141)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_13),
.B1(n_20),
.B2(n_17),
.C(n_21),
.Y(n_132)
);

AOI322xp5_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_21),
.A3(n_24),
.B1(n_23),
.B2(n_19),
.C1(n_16),
.C2(n_26),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_131),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_126),
.B(n_7),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_135),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_137),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_17),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_138),
.B(n_144),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_115),
.B(n_124),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_20),
.B1(n_21),
.B2(n_10),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_148),
.B1(n_128),
.B2(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_20),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_26),
.B1(n_21),
.B2(n_16),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_53),
.C(n_24),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_120),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_26),
.B1(n_23),
.B2(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_158),
.B1(n_111),
.B2(n_129),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_121),
.B(n_117),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_130),
.B(n_125),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_160),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_139),
.B1(n_117),
.B2(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_143),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_137),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_170),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_166),
.A2(n_172),
.B1(n_7),
.B2(n_6),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_169),
.B(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_147),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_8),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_151),
.A2(n_136),
.B1(n_113),
.B2(n_138),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_162),
.B1(n_150),
.B2(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_174),
.B(n_175),
.Y(n_183)
);

OAI221xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_153),
.B1(n_155),
.B2(n_159),
.C(n_7),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_176),
.B(n_6),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_179),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_23),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_189),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_164),
.B(n_172),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_2),
.B(n_3),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_19),
.C(n_23),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_19),
.C(n_1),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_185),
.B(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_192),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_177),
.B(n_19),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_2),
.C(n_3),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_197),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_4),
.C(n_5),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_4),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_201),
.A2(n_196),
.B(n_198),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule