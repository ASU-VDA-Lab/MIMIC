module fake_jpeg_4868_n_300 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_287;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_53),
.Y(n_72)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_47),
.B1(n_59),
.B2(n_24),
.Y(n_74)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_65),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_61),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_69),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_23),
.B(n_1),
.CON(n_63),
.SN(n_63)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_28),
.Y(n_93)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_67),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_26),
.B1(n_25),
.B2(n_23),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_98),
.B1(n_38),
.B2(n_41),
.Y(n_121)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_26),
.B1(n_36),
.B2(n_25),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_80),
.A2(n_96),
.B1(n_109),
.B2(n_41),
.Y(n_134)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_88),
.Y(n_119)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_90),
.Y(n_120)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_93),
.Y(n_123)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_100),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_27),
.B1(n_29),
.B2(n_37),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_46),
.A2(n_37),
.B1(n_39),
.B2(n_20),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_107),
.B1(n_1),
.B2(n_2),
.Y(n_122)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_47),
.A2(n_59),
.B1(n_19),
.B2(n_39),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_20),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_111),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_55),
.A2(n_38),
.B1(n_19),
.B2(n_58),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_132),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_60),
.C(n_43),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_131),
.C(n_82),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_70),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_128),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_121),
.A2(n_137),
.B1(n_143),
.B2(n_7),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_141),
.B(n_5),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_77),
.B(n_110),
.Y(n_124)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_138),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_86),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_134),
.C(n_5),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_60),
.C(n_43),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_60),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_43),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_146),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_81),
.A2(n_43),
.B1(n_41),
.B2(n_30),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_142),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_93),
.A2(n_41),
.B(n_4),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_71),
.B(n_2),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_87),
.A2(n_16),
.B1(n_15),
.B2(n_6),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_2),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_101),
.B1(n_113),
.B2(n_75),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_151),
.A2(n_179),
.B1(n_155),
.B2(n_149),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_168),
.B1(n_9),
.B2(n_10),
.Y(n_205)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_145),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_79),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_79),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_74),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_115),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_5),
.Y(n_165)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_101),
.B1(n_103),
.B2(n_88),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_175),
.B1(n_180),
.B2(n_139),
.Y(n_198)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_132),
.A2(n_133),
.B(n_123),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_127),
.B(n_149),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_85),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_129),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_136),
.A2(n_95),
.B1(n_85),
.B2(n_84),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_119),
.Y(n_176)
);

INVx6_ASAP7_75t_SL g193 ( 
.A(n_176),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_116),
.Y(n_178)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_178),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_126),
.B1(n_144),
.B2(n_138),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_13),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_142),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_187),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_148),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_84),
.B(n_95),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_190),
.A2(n_193),
.B(n_198),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_194),
.A2(n_200),
.B(n_201),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_148),
.C(n_127),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_197),
.C(n_207),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_202),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_210),
.B1(n_211),
.B2(n_182),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_161),
.A2(n_147),
.B(n_10),
.C(n_12),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_147),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_9),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_162),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_173),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_145),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_153),
.A2(n_167),
.B1(n_163),
.B2(n_175),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_151),
.A2(n_179),
.B1(n_174),
.B2(n_168),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_212),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_220),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_219),
.B1(n_227),
.B2(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_156),
.B1(n_171),
.B2(n_169),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_185),
.B(n_159),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_194),
.A2(n_181),
.B(n_170),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_200),
.B(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_170),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_170),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_15),
.B1(n_16),
.B2(n_166),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_14),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_184),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_SL g230 ( 
.A(n_183),
.B(n_193),
.C(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_202),
.B(n_188),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_232),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_185),
.B(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_191),
.B(n_195),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_249),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_228),
.A2(n_190),
.B1(n_203),
.B2(n_197),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_207),
.C(n_206),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_244),
.Y(n_255)
);

AO21x1_ASAP7_75t_L g243 ( 
.A1(n_235),
.A2(n_190),
.B(n_201),
.Y(n_243)
);

NOR3xp33_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_246),
.C(n_213),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_207),
.C(n_192),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_192),
.C(n_209),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_250),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_SL g246 ( 
.A(n_234),
.B(n_189),
.C(n_212),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_189),
.B1(n_195),
.B2(n_191),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_184),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_221),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_213),
.B1(n_225),
.B2(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_253),
.B(n_254),
.Y(n_267)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_266),
.C(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_264),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_241),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_271),
.Y(n_279)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_255),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_240),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_251),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_241),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_276),
.B(n_238),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_249),
.B(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

OAI31xp33_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_264),
.A3(n_259),
.B(n_256),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_278),
.A2(n_280),
.B(n_281),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_276),
.A2(n_256),
.B(n_230),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_267),
.B(n_248),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_255),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_285),
.A2(n_232),
.B(n_274),
.C(n_233),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_292),
.B(n_283),
.Y(n_295)
);

NOR4xp25_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_279),
.C(n_289),
.D(n_287),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_232),
.B(n_227),
.C(n_222),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_215),
.B1(n_222),
.B2(n_284),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_279),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_294),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_295),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_296),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_297),
.Y(n_300)
);


endmodule