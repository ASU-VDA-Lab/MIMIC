module real_jpeg_3513_n_27 (n_17, n_8, n_0, n_21, n_141, n_2, n_142, n_143, n_10, n_9, n_12, n_147, n_24, n_146, n_6, n_151, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_145, n_144, n_5, n_4, n_150, n_1, n_26, n_20, n_19, n_148, n_149, n_16, n_15, n_13, n_27);

input n_17;
input n_8;
input n_0;
input n_21;
input n_141;
input n_2;
input n_142;
input n_143;
input n_10;
input n_9;
input n_12;
input n_147;
input n_24;
input n_146;
input n_6;
input n_151;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_145;
input n_144;
input n_5;
input n_4;
input n_150;
input n_1;
input n_26;
input n_20;
input n_19;
input n_148;
input n_149;
input n_16;
input n_15;
input n_13;

output n_27;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_139;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_0),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_2),
.Y(n_109)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_3),
.A2(n_65),
.B1(n_68),
.B2(n_78),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_5),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_6),
.B(n_64),
.C(n_79),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_7),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_9),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_10),
.B(n_62),
.C(n_87),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_11),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_12),
.A2(n_60),
.B1(n_93),
.B2(n_96),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_12),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_13),
.A2(n_135),
.B1(n_136),
.B2(n_139),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_13),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_16),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_18),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_20),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_21),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_21),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_22),
.B(n_42),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_24),
.A2(n_70),
.B(n_74),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_26),
.B(n_55),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_134),
.Y(n_27)
);

MAJx2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_130),
.C(n_131),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_39),
.B(n_129),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_38),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_31),
.B(n_38),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_34),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_34),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_34),
.B(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_34),
.Y(n_138)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx6p67_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_37),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_37),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_45),
.C(n_128),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

MAJx2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_124),
.C(n_125),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_123),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_48),
.B(n_52),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_92),
.Y(n_91)
);

OAI221xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B1(n_59),
.B2(n_99),
.C(n_113),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_56),
.B(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_89),
.C(n_90),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_82),
.C(n_83),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_75),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.C(n_77),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_74),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_108),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_114),
.A3(n_115),
.B1(n_118),
.B2(n_119),
.C1(n_122),
.C2(n_151),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.C(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_141),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_142),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_143),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_144),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_145),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_146),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_147),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_148),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_149),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_150),
.Y(n_112)
);


endmodule