module fake_jpeg_19130_n_58 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_24),
.B(n_6),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_41),
.B(n_44),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_23),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_3),
.C(n_7),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_45),
.B(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_10),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_51),
.B(n_16),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_15),
.C(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_18),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_19),
.B(n_20),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_21),
.Y(n_58)
);


endmodule