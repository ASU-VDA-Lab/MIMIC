module fake_aes_1277_n_682 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_682);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_682;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_70), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_76), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_4), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_41), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_26), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_39), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_62), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_75), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_46), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_29), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_13), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_59), .Y(n_91) );
INVx1_ASAP7_75t_SL g92 ( .A(n_5), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_32), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_73), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_20), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_71), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g97 ( .A(n_65), .B(n_22), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_60), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_51), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_21), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_53), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_72), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_6), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_23), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_68), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_27), .Y(n_106) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_7), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_61), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_48), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_69), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_55), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_42), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_58), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_66), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_50), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_15), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_44), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_52), .Y(n_121) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_28), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_37), .Y(n_123) );
BUFx2_ASAP7_75t_SL g124 ( .A(n_3), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_19), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_43), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_8), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_109), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_110), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_95), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_110), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_103), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_90), .B(n_0), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_88), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_115), .Y(n_141) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_111), .Y(n_143) );
NAND2xp33_ASAP7_75t_SL g144 ( .A(n_80), .B(n_0), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_127), .B(n_1), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_107), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_126), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_99), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
BUFx8_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_119), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_91), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_79), .B(n_2), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_91), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_93), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_93), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_94), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_79), .B(n_4), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_94), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_96), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_112), .B(n_6), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_100), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_112), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_116), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_167), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_168), .B(n_104), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_167), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_168), .B(n_100), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_157), .B(n_92), .Y(n_175) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_167), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_128), .B(n_98), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
NOR2x1p5_ASAP7_75t_L g179 ( .A(n_149), .B(n_104), .Y(n_179) );
NAND3xp33_ASAP7_75t_L g180 ( .A(n_162), .B(n_105), .C(n_123), .Y(n_180) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_145), .A2(n_97), .B(n_116), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_135), .B(n_105), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_153), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_141), .B(n_124), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_132), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_133), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_170), .Y(n_188) );
INVxp67_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
AOI22x1_ASAP7_75t_L g190 ( .A1(n_170), .A2(n_123), .B1(n_106), .B2(n_102), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_170), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_165), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_163), .Y(n_193) );
NAND2xp33_ASAP7_75t_SL g194 ( .A(n_163), .B(n_84), .Y(n_194) );
AO22x2_ASAP7_75t_L g195 ( .A1(n_138), .A2(n_82), .B1(n_85), .B2(n_121), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_148), .B(n_89), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_153), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_152), .A2(n_107), .B1(n_122), .B2(n_118), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_169), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_138), .B(n_120), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_155), .B(n_125), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_139), .B(n_86), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_156), .B(n_83), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_165), .Y(n_205) );
OR2x2_ASAP7_75t_SL g206 ( .A(n_136), .B(n_117), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_166), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_130), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
AND2x6_ASAP7_75t_L g210 ( .A(n_139), .B(n_101), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_166), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_158), .B(n_122), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_153), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_140), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_169), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_140), .B(n_118), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_159), .B(n_113), .Y(n_217) );
AND2x6_ASAP7_75t_L g218 ( .A(n_160), .B(n_34), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_161), .B(n_7), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_129), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_152), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_129), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_130), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_131), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_152), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_154), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_131), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_164), .B(n_8), .Y(n_229) );
NOR3xp33_ASAP7_75t_L g230 ( .A(n_144), .B(n_9), .C(n_10), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_154), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_134), .B(n_36), .Y(n_232) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_143), .A2(n_38), .B(n_77), .Y(n_233) );
INVx4_ASAP7_75t_L g234 ( .A(n_130), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_143), .B(n_10), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_188), .Y(n_236) );
BUFx4f_ASAP7_75t_SL g237 ( .A(n_226), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_189), .B(n_147), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_188), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_188), .Y(n_240) );
INVx5_ASAP7_75t_L g241 ( .A(n_218), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_229), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_191), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_212), .B(n_146), .Y(n_244) );
INVx2_ASAP7_75t_SL g245 ( .A(n_176), .Y(n_245) );
BUFx4f_ASAP7_75t_L g246 ( .A(n_218), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_193), .Y(n_247) );
INVx1_ASAP7_75t_SL g248 ( .A(n_174), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_195), .A2(n_169), .B1(n_146), .B2(n_151), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_229), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_195), .A2(n_169), .B1(n_151), .B2(n_150), .Y(n_251) );
INVx5_ASAP7_75t_L g252 ( .A(n_218), .Y(n_252) );
INVx1_ASAP7_75t_SL g253 ( .A(n_172), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_193), .Y(n_255) );
BUFx12f_ASAP7_75t_SL g256 ( .A(n_184), .Y(n_256) );
INVx5_ASAP7_75t_L g257 ( .A(n_218), .Y(n_257) );
BUFx12f_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_186), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_201), .B(n_150), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_201), .B(n_137), .Y(n_261) );
NOR2xp67_ASAP7_75t_L g262 ( .A(n_199), .B(n_11), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_185), .Y(n_263) );
INVx5_ASAP7_75t_L g264 ( .A(n_218), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_187), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_185), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_223), .Y(n_267) );
AND3x1_ASAP7_75t_L g268 ( .A(n_230), .B(n_144), .C(n_12), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_201), .B(n_137), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_223), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_196), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_203), .B(n_197), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_189), .A2(n_137), .B1(n_130), .B2(n_154), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_208), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_208), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_210), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_202), .B(n_137), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_183), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_210), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_183), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_220), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_195), .A2(n_154), .B1(n_137), .B2(n_130), .Y(n_283) );
BUFx8_ASAP7_75t_L g284 ( .A(n_216), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_222), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_175), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_183), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_221), .Y(n_288) );
INVx5_ASAP7_75t_L g289 ( .A(n_210), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_210), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_176), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_183), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_178), .B(n_11), .Y(n_293) );
INVx5_ASAP7_75t_L g294 ( .A(n_210), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_175), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_196), .Y(n_296) );
AOI22x1_ASAP7_75t_L g297 ( .A1(n_234), .A2(n_40), .B1(n_74), .B2(n_67), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_198), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_198), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_213), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_182), .B(n_33), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_213), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_227), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_204), .B(n_12), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_245), .B(n_179), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_236), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_295), .B(n_194), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_284), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_289), .B(n_203), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_247), .B(n_226), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_238), .A2(n_203), .B1(n_171), .B2(n_173), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_286), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_277), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_265), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_236), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_277), .Y(n_317) );
BUFx8_ASAP7_75t_SL g318 ( .A(n_258), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
NAND2x1p5_ASAP7_75t_L g320 ( .A(n_280), .B(n_219), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_239), .Y(n_321) );
NAND2xp5_ASAP7_75t_SL g322 ( .A(n_289), .B(n_214), .Y(n_322) );
BUFx4f_ASAP7_75t_L g323 ( .A(n_258), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_238), .A2(n_216), .B1(n_230), .B2(n_190), .Y(n_324) );
AOI21x1_ASAP7_75t_L g325 ( .A1(n_250), .A2(n_192), .B(n_211), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_242), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_260), .Y(n_327) );
BUFx8_ASAP7_75t_SL g328 ( .A(n_288), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_245), .B(n_180), .Y(n_329) );
AND2x6_ASAP7_75t_SL g330 ( .A(n_237), .B(n_177), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_253), .B(n_206), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_239), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_243), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_290), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_278), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_282), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_291), .B(n_217), .Y(n_337) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_261), .A2(n_233), .B(n_181), .Y(n_338) );
INVx5_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_248), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_278), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_278), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_255), .A2(n_194), .B1(n_177), .B2(n_207), .C(n_205), .Y(n_343) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_246), .B(n_232), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_289), .B(n_234), .Y(n_345) );
INVx6_ASAP7_75t_L g346 ( .A(n_284), .Y(n_346) );
INVx6_ASAP7_75t_L g347 ( .A(n_284), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_256), .Y(n_348) );
CKINVDCx8_ASAP7_75t_R g349 ( .A(n_288), .Y(n_349) );
HAxp5_ASAP7_75t_L g350 ( .A(n_256), .B(n_181), .CON(n_350), .SN(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_242), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_238), .B(n_216), .Y(n_352) );
OR2x6_ASAP7_75t_SL g353 ( .A(n_272), .B(n_216), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_274), .Y(n_354) );
INVx3_ASAP7_75t_SL g355 ( .A(n_304), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_304), .Y(n_356) );
AND2x6_ASAP7_75t_L g357 ( .A(n_290), .B(n_224), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_306), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_307), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_346), .B(n_242), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_314), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_339), .B(n_289), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_333), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_336), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_352), .B(n_291), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_328), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_314), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_315), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_328), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_336), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_356), .A2(n_254), .B1(n_251), .B2(n_249), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_316), .Y(n_376) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_321), .A2(n_246), .B(n_301), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_331), .A2(n_262), .B1(n_304), .B2(n_293), .C1(n_244), .C2(n_216), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_325), .A2(n_297), .B(n_283), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_331), .A2(n_240), .B1(n_285), .B2(n_301), .Y(n_380) );
OAI22xp33_ASAP7_75t_SL g381 ( .A1(n_355), .A2(n_268), .B1(n_246), .B2(n_264), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_312), .A2(n_337), .B1(n_343), .B2(n_311), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_312), .B(n_249), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_321), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_355), .A2(n_251), .B1(n_283), .B2(n_257), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_313), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_327), .B(n_228), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_337), .A2(n_274), .B1(n_275), .B2(n_276), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_320), .A2(n_257), .B1(n_264), .B2(n_252), .Y(n_390) );
AND2x4_ASAP7_75t_SL g391 ( .A(n_360), .B(n_305), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g392 ( .A1(n_378), .A2(n_308), .B(n_324), .Y(n_392) );
AOI222xp33_ASAP7_75t_L g393 ( .A1(n_382), .A2(n_323), .B1(n_324), .B2(n_305), .C1(n_348), .C2(n_341), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_383), .A2(n_347), .B1(n_346), .B2(n_329), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_383), .A2(n_347), .B1(n_346), .B2(n_329), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_358), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_360), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_372), .Y(n_399) );
AOI211xp5_ASAP7_75t_L g400 ( .A1(n_381), .A2(n_342), .B(n_309), .C(n_235), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_364), .A2(n_353), .B1(n_320), .B2(n_344), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_387), .B(n_350), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_387), .B(n_350), .Y(n_403) );
AO31x2_ASAP7_75t_L g404 ( .A1(n_364), .A2(n_227), .A3(n_332), .B(n_269), .Y(n_404) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_380), .A2(n_273), .B(n_344), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_375), .A2(n_326), .B(n_351), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_365), .Y(n_407) );
CKINVDCx14_ASAP7_75t_R g408 ( .A(n_369), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_370), .A2(n_309), .B(n_351), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_365), .A2(n_347), .B1(n_326), .B2(n_349), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_368), .A2(n_323), .B1(n_354), .B2(n_318), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_368), .A2(n_354), .B1(n_318), .B2(n_338), .Y(n_412) );
OAI211xp5_ASAP7_75t_L g413 ( .A1(n_386), .A2(n_310), .B(n_234), .C(n_322), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_368), .A2(n_338), .B1(n_310), .B2(n_357), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_367), .A2(n_357), .B1(n_264), .B2(n_257), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_388), .A2(n_330), .B1(n_275), .B2(n_274), .C(n_276), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_374), .A2(n_357), .B1(n_241), .B2(n_252), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_396), .Y(n_418) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_396), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_L g420 ( .A1(n_392), .A2(n_385), .B(n_376), .C(n_384), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_393), .A2(n_360), .B1(n_389), .B2(n_377), .C(n_384), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_407), .Y(n_422) );
NAND4xp25_ASAP7_75t_L g423 ( .A(n_411), .B(n_209), .C(n_200), .D(n_215), .Y(n_423) );
AND2x4_ASAP7_75t_SL g424 ( .A(n_398), .B(n_360), .Y(n_424) );
AOI31xp33_ASAP7_75t_L g425 ( .A1(n_408), .A2(n_369), .A3(n_373), .B(n_363), .Y(n_425) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_408), .A2(n_373), .A3(n_376), .B1(n_13), .B2(n_14), .C1(n_358), .C2(n_366), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_402), .B(n_366), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_402), .A2(n_362), .B1(n_241), .B2(n_252), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_394), .A2(n_362), .B1(n_252), .B2(n_241), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_403), .A2(n_275), .B1(n_276), .B2(n_209), .C(n_200), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_404), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_403), .B(n_371), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_397), .A2(n_209), .B1(n_215), .B2(n_361), .C(n_371), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_407), .B(n_361), .Y(n_434) );
OA21x2_ASAP7_75t_L g435 ( .A1(n_406), .A2(n_379), .B(n_322), .Y(n_435) );
AOI33xp33_ASAP7_75t_L g436 ( .A1(n_399), .A2(n_14), .A3(n_298), .B1(n_303), .B2(n_271), .B3(n_302), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
AND2x4_ASAP7_75t_SL g439 ( .A(n_398), .B(n_395), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_391), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_404), .Y(n_441) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_405), .A2(n_379), .B(n_390), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_412), .B(n_371), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_400), .B(n_361), .C(n_225), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_401), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_409), .A2(n_241), .B1(n_233), .B2(n_334), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_410), .A2(n_241), .B1(n_319), .B2(n_334), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_416), .A2(n_231), .B1(n_225), .B2(n_345), .C(n_270), .Y(n_449) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_413), .A2(n_345), .B(n_263), .Y(n_450) );
AOI21xp33_ASAP7_75t_L g451 ( .A1(n_414), .A2(n_334), .B(n_319), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_391), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_427), .B(n_17), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_427), .B(n_415), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_422), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_422), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_424), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_437), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_443), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_445), .B(n_363), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_443), .Y(n_461) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_445), .A2(n_296), .B(n_303), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_431), .Y(n_463) );
OAI31xp33_ASAP7_75t_L g464 ( .A1(n_421), .A2(n_446), .A3(n_439), .B(n_426), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_437), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_438), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_418), .B(n_18), .Y(n_468) );
NAND2xp33_ASAP7_75t_SL g469 ( .A(n_440), .B(n_417), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_438), .Y(n_470) );
AOI33xp33_ASAP7_75t_L g471 ( .A1(n_439), .A2(n_296), .A3(n_298), .B1(n_299), .B2(n_271), .B3(n_300), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_418), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_441), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_432), .B(n_24), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_440), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_446), .A2(n_319), .B(n_317), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_441), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_434), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_432), .B(n_25), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_419), .B(n_30), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_435), .Y(n_482) );
INVx5_ASAP7_75t_L g483 ( .A(n_452), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_435), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_444), .B(n_231), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_434), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_442), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_444), .B(n_231), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_452), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_425), .B(n_299), .C(n_300), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_451), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_420), .A2(n_319), .B1(n_317), .B2(n_314), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_442), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_449), .A2(n_294), .B(n_317), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_436), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_450), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_442), .B(n_31), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_433), .B(n_231), .C(n_225), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_423), .B(n_314), .Y(n_501) );
OAI31xp33_ASAP7_75t_SL g502 ( .A1(n_448), .A2(n_35), .A3(n_45), .B(n_47), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_487), .B(n_450), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_478), .B(n_442), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_487), .B(n_447), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_456), .B(n_428), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_465), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_455), .B(n_429), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_455), .B(n_430), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_458), .B(n_49), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_467), .B(n_225), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_467), .B(n_54), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_458), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_467), .B(n_470), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_464), .B(n_270), .C(n_267), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_470), .B(n_56), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_477), .B(n_63), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_473), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_459), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_473), .Y(n_520) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_497), .A2(n_302), .B(n_263), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_477), .B(n_64), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_472), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_490), .B(n_78), .Y(n_524) );
NAND4xp25_ASAP7_75t_SL g525 ( .A(n_464), .B(n_339), .C(n_294), .D(n_317), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_477), .B(n_267), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_472), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_472), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_466), .B(n_267), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_466), .B(n_267), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_457), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_497), .B(n_270), .Y(n_532) );
BUFx2_ASAP7_75t_SL g533 ( .A(n_475), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_453), .B(n_270), .Y(n_534) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_459), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_460), .A2(n_294), .B(n_339), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_459), .B(n_266), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_500), .A2(n_294), .B(n_279), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_461), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_461), .Y(n_540) );
NAND5xp2_ASAP7_75t_L g541 ( .A(n_502), .B(n_294), .C(n_279), .D(n_281), .E(n_287), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_461), .B(n_279), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_454), .B(n_281), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_453), .B(n_281), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_475), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_490), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_479), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_490), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_469), .B(n_287), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
NOR3xp33_ASAP7_75t_SL g551 ( .A(n_501), .B(n_292), .C(n_492), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_463), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_491), .A2(n_292), .B1(n_480), .B2(n_474), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_531), .B(n_483), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_513), .Y(n_555) );
NAND2x1p5_ASAP7_75t_L g556 ( .A(n_524), .B(n_483), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_518), .B(n_463), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_533), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_520), .Y(n_559) );
AND4x1_ASAP7_75t_L g560 ( .A(n_515), .B(n_471), .C(n_500), .D(n_480), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_514), .B(n_489), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_553), .A2(n_483), .B(n_499), .C(n_468), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_545), .B(n_483), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_539), .B(n_485), .Y(n_564) );
XOR2x2_ASAP7_75t_L g565 ( .A(n_524), .B(n_468), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_550), .B(n_483), .Y(n_566) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_551), .B(n_483), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_535), .B(n_484), .Y(n_568) );
NOR2x1_ASAP7_75t_L g569 ( .A(n_541), .B(n_462), .Y(n_569) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_525), .A2(n_499), .B(n_496), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_505), .B(n_479), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_546), .B(n_486), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_548), .B(n_476), .Y(n_573) );
NOR2xp67_ASAP7_75t_SL g574 ( .A(n_517), .B(n_495), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_552), .B(n_482), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_507), .Y(n_576) );
INVx4_ASAP7_75t_SL g577 ( .A(n_524), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_509), .B(n_482), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_507), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_523), .Y(n_580) );
AOI32xp33_ASAP7_75t_L g581 ( .A1(n_510), .A2(n_493), .A3(n_498), .B1(n_486), .B2(n_484), .Y(n_581) );
OAI31xp33_ASAP7_75t_L g582 ( .A1(n_510), .A2(n_498), .A3(n_484), .B(n_486), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_527), .B(n_494), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_528), .B(n_494), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_506), .B(n_462), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_552), .B(n_494), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_519), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_519), .B(n_488), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_540), .B(n_488), .Y(n_589) );
CKINVDCx16_ASAP7_75t_R g590 ( .A(n_534), .Y(n_590) );
INVx2_ASAP7_75t_SL g591 ( .A(n_529), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_510), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_530), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_540), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_503), .B(n_488), .Y(n_595) );
INVx2_ASAP7_75t_SL g596 ( .A(n_537), .Y(n_596) );
INVx2_ASAP7_75t_SL g597 ( .A(n_537), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_590), .B(n_526), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_565), .A2(n_532), .B1(n_549), .B2(n_521), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_568), .Y(n_600) );
AOI21xp33_ASAP7_75t_L g601 ( .A1(n_585), .A2(n_549), .B(n_516), .Y(n_601) );
NAND2x1_ASAP7_75t_L g602 ( .A(n_569), .B(n_512), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_571), .A2(n_504), .B(n_508), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_558), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_559), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_555), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_558), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_593), .B(n_543), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_575), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_580), .Y(n_610) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_567), .B(n_516), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_577), .B(n_547), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_557), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_596), .Y(n_614) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_573), .A2(n_512), .B(n_522), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_595), .B(n_511), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_593), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_581), .A2(n_517), .B(n_522), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_554), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_561), .B(n_544), .Y(n_620) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_556), .Y(n_621) );
INVx4_ASAP7_75t_L g622 ( .A(n_577), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_572), .Y(n_623) );
NAND2x1_ASAP7_75t_L g624 ( .A(n_586), .B(n_538), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_591), .B(n_542), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_576), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_563), .B(n_536), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_579), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_592), .A2(n_597), .B1(n_566), .B2(n_564), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_570), .A2(n_574), .B1(n_582), .B2(n_586), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_594), .Y(n_631) );
NAND2xp33_ASAP7_75t_SL g632 ( .A(n_560), .B(n_570), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_589), .B(n_583), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_584), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_560), .B(n_587), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_588), .Y(n_636) );
XNOR2x1_ASAP7_75t_L g637 ( .A(n_582), .B(n_562), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_556), .Y(n_638) );
O2A1O1Ixp5_ASAP7_75t_L g639 ( .A1(n_566), .A2(n_585), .B(n_554), .C(n_578), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_559), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_558), .B(n_569), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_558), .B(n_569), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_558), .B(n_569), .Y(n_643) );
XNOR2x1_ASAP7_75t_L g644 ( .A(n_565), .B(n_408), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_569), .A2(n_464), .B1(n_403), .B2(n_402), .Y(n_645) );
OAI21xp33_ASAP7_75t_SL g646 ( .A1(n_641), .A2(n_642), .B(n_643), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_632), .A2(n_637), .B(n_644), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_623), .Y(n_648) );
XNOR2x1_ASAP7_75t_L g649 ( .A(n_604), .B(n_611), .Y(n_649) );
XNOR2x1_ASAP7_75t_L g650 ( .A(n_604), .B(n_617), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_607), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_645), .A2(n_630), .B(n_635), .C(n_622), .Y(n_652) );
NOR2xp67_ASAP7_75t_L g653 ( .A(n_622), .B(n_630), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_617), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_634), .B(n_636), .Y(n_655) );
AOI331xp33_ASAP7_75t_L g656 ( .A1(n_645), .A2(n_613), .A3(n_605), .B1(n_606), .B2(n_640), .B3(n_610), .C1(n_608), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_639), .B(n_629), .C(n_602), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_633), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_629), .A2(n_603), .B1(n_618), .B2(n_601), .C(n_619), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_647), .A2(n_621), .B(n_624), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_656), .B(n_628), .Y(n_661) );
NOR2x1p5_ASAP7_75t_L g662 ( .A(n_646), .B(n_638), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_649), .A2(n_614), .B1(n_638), .B2(n_599), .Y(n_663) );
OAI22x1_ASAP7_75t_L g664 ( .A1(n_651), .A2(n_612), .B1(n_600), .B2(n_598), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_657), .A2(n_627), .B1(n_601), .B2(n_615), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_652), .B(n_626), .C(n_631), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_653), .A2(n_612), .B1(n_609), .B2(n_620), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_666), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_663), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_664), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_661), .B(n_650), .Y(n_671) );
INVxp67_ASAP7_75t_SL g672 ( .A(n_662), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_669), .A2(n_665), .B1(n_660), .B2(n_667), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_670), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_668), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_673), .A2(n_671), .B1(n_672), .B2(n_668), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_674), .Y(n_677) );
OR2x6_ASAP7_75t_L g678 ( .A(n_677), .B(n_675), .Y(n_678) );
NOR3x1_ASAP7_75t_L g679 ( .A(n_676), .B(n_655), .C(n_648), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_678), .A2(n_659), .B1(n_654), .B2(n_655), .Y(n_680) );
XNOR2xp5_ASAP7_75t_L g681 ( .A(n_680), .B(n_679), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_658), .B1(n_625), .B2(n_616), .Y(n_682) );
endmodule