module fake_jpeg_25759_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_18),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_46),
.B(n_62),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_32),
.B1(n_16),
.B2(n_26),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_36),
.B1(n_20),
.B2(n_26),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_28),
.C(n_33),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_22),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_60),
.B1(n_66),
.B2(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_61),
.B(n_65),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2x1_ASAP7_75t_R g65 ( 
.A(n_41),
.B(n_28),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_16),
.B1(n_28),
.B2(n_30),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_22),
.B1(n_34),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_17),
.B1(n_30),
.B2(n_21),
.Y(n_69)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_69),
.A2(n_75),
.B1(n_101),
.B2(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_73),
.C(n_84),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_72),
.B(n_80),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_55),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_76),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_95),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_81),
.B(n_86),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_96),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_87),
.A2(n_89),
.B1(n_102),
.B2(n_104),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

AO22x2_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_39),
.B1(n_36),
.B2(n_44),
.Y(n_89)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_25),
.A3(n_27),
.B1(n_31),
.B2(n_34),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_17),
.Y(n_114)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_27),
.Y(n_94)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_52),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_17),
.B1(n_26),
.B2(n_24),
.Y(n_111)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_25),
.B1(n_31),
.B2(n_22),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_54),
.B1(n_57),
.B2(n_51),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_49),
.A2(n_44),
.B1(n_17),
.B2(n_21),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_59),
.A2(n_19),
.B1(n_29),
.B2(n_35),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_39),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_40),
.C(n_36),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_33),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_83),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_20),
.B(n_24),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_117),
.A2(n_20),
.B(n_24),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_72),
.B(n_26),
.CI(n_20),
.CON(n_125),
.SN(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_103),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_19),
.B1(n_29),
.B2(n_35),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_92),
.B1(n_29),
.B2(n_19),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_75),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_134),
.B(n_100),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_26),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_138),
.C(n_107),
.Y(n_150)
);

AOI22x1_ASAP7_75t_L g136 ( 
.A1(n_89),
.A2(n_40),
.B1(n_36),
.B2(n_26),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_89),
.B1(n_87),
.B2(n_102),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_40),
.C(n_36),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_139),
.B(n_147),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_141),
.A2(n_167),
.B1(n_135),
.B2(n_118),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_145),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_146),
.B1(n_149),
.B2(n_164),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_144),
.A2(n_152),
.B(n_158),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_70),
.B1(n_75),
.B2(n_84),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_73),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_153),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_115),
.A2(n_84),
.B1(n_73),
.B2(n_77),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_151),
.C(n_161),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_91),
.C(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_35),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_155),
.B(n_159),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_162),
.Y(n_178)
);

AOI32xp33_ASAP7_75t_L g158 ( 
.A1(n_114),
.A2(n_99),
.A3(n_98),
.B1(n_95),
.B2(n_88),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_78),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_124),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_88),
.C(n_40),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_119),
.A2(n_85),
.B1(n_100),
.B2(n_90),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_126),
.B(n_90),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_155),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_136),
.B1(n_116),
.B2(n_117),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_131),
.B1(n_121),
.B2(n_112),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_145),
.B1(n_143),
.B2(n_170),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_140),
.B(n_144),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_85),
.B1(n_76),
.B2(n_71),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_110),
.B1(n_121),
.B2(n_112),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

OAI22x1_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_110),
.B1(n_131),
.B2(n_122),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_174),
.A2(n_200),
.B1(n_0),
.B2(n_2),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_175),
.A2(n_198),
.B(n_203),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_181),
.B1(n_184),
.B2(n_197),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_187),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_182),
.B1(n_150),
.B2(n_168),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_134),
.B1(n_120),
.B2(n_79),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_167),
.A2(n_105),
.B1(n_26),
.B2(n_24),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_24),
.B1(n_20),
.B2(n_33),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_20),
.B1(n_24),
.B2(n_33),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_185),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_230)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_189),
.B(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_195),
.B(n_201),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_144),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_36),
.C(n_23),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_154),
.C(n_163),
.Y(n_211)
);

OAI22x1_ASAP7_75t_L g200 ( 
.A1(n_151),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_157),
.B(n_148),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_191),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_222),
.B1(n_223),
.B2(n_226),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_147),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_219),
.C(n_227),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_139),
.B1(n_1),
.B2(n_2),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_8),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_15),
.C(n_13),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_187),
.A2(n_172),
.B1(n_192),
.B2(n_179),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_221),
.B1(n_230),
.B2(n_210),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_182),
.A2(n_200),
.B1(n_180),
.B2(n_195),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_0),
.B(n_2),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_172),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_176),
.B1(n_193),
.B2(n_178),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_0),
.B(n_3),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_184),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_12),
.C(n_10),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_189),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

AOI21x1_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_203),
.B(n_196),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_225),
.B(n_209),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_217),
.B1(n_213),
.B2(n_205),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_199),
.C(n_176),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_249),
.C(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_241),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_224),
.Y(n_269)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_252),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_197),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_251),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_183),
.C(n_202),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_202),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_208),
.Y(n_252)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_9),
.C(n_10),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_254),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_256),
.C(n_259),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_231),
.C(n_220),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_261),
.B(n_234),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_222),
.C(n_227),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_219),
.C(n_210),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_263),
.Y(n_287)
);

NOR2x1p5_ASAP7_75t_SL g261 ( 
.A(n_251),
.B(n_209),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_262),
.A2(n_272),
.B1(n_234),
.B2(n_257),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_247),
.B(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_249),
.B(n_216),
.Y(n_268)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_239),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_223),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_216),
.C(n_230),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_240),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_254),
.B1(n_237),
.B2(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_285),
.B(n_4),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_246),
.B1(n_244),
.B2(n_240),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_250),
.C(n_235),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_286),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_248),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_282),
.C(n_284),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_242),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_242),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_270),
.A2(n_252),
.B1(n_238),
.B2(n_241),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_288),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_258),
.B(n_264),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_282),
.B(n_284),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_256),
.CI(n_273),
.CON(n_293),
.SN(n_293)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_277),
.Y(n_301)
);

OAI32xp33_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_269),
.A3(n_260),
.B1(n_259),
.B2(n_7),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_280),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_6),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_286),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_288),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_303),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_306),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_296),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_277),
.B(n_281),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_292),
.B(n_307),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_299),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_291),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_315),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_290),
.C(n_291),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_312),
.B1(n_310),
.B2(n_297),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_293),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_314),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_SL g321 ( 
.A(n_319),
.B(n_320),
.C(n_317),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_321),
.A2(n_320),
.B(n_290),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_322),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_323),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_309),
.Y(n_325)
);


endmodule