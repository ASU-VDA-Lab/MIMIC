module fake_netlist_6_1687_n_1295 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1295);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1295;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g315 ( 
.A(n_79),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_291),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_212),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_214),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_63),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_192),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_13),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_243),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_139),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_280),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_65),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_76),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_167),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_92),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_74),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_211),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_242),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_181),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_141),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_123),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_82),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_275),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_25),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_142),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_262),
.B(n_22),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_303),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_220),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_161),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_271),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_14),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_108),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_76),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_114),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_1),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_230),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_111),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_250),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_131),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_160),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_238),
.B(n_53),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_196),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_189),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_81),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_208),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_124),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_16),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_93),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_82),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_72),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_236),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_56),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_19),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_182),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_263),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_170),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_137),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_72),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_191),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_281),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_54),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_132),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_98),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_54),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_194),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_150),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_152),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_62),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_201),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_148),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_255),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_277),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_292),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_297),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_284),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_92),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_195),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_144),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_166),
.B(n_254),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_268),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_8),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_27),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_36),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_184),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_104),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_256),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_293),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_52),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_163),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_8),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_143),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_12),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_229),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_215),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_6),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_75),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_157),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_30),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_279),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_133),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_221),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_190),
.B(n_172),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_155),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_200),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_239),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_289),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_217),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_67),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_186),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_247),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_17),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_197),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_267),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_314),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_14),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_162),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_106),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_29),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_50),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_126),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_219),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_251),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_35),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_171),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_210),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_296),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_88),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_122),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_25),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_113),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_115),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_147),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_282),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_300),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_273),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_51),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_52),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_95),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_299),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_110),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_75),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_164),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_33),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_53),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_116),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_261),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_231),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_91),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_13),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_209),
.Y(n_466)
);

BUFx8_ASAP7_75t_L g467 ( 
.A(n_459),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_335),
.B(n_0),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_374),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_324),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_324),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_457),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_324),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_335),
.B(n_0),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_374),
.B(n_1),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_377),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_324),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_315),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_414),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_322),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_322),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_320),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_328),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_342),
.B(n_2),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_330),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_331),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_370),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_370),
.Y(n_491)
);

OAI22x1_ASAP7_75t_L g492 ( 
.A1(n_439),
.A2(n_366),
.B1(n_408),
.B2(n_369),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_409),
.B(n_3),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_364),
.Y(n_494)
);

OA21x2_ASAP7_75t_L g495 ( 
.A1(n_318),
.A2(n_4),
.B(n_5),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_399),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_367),
.A2(n_107),
.B(n_105),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_349),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_366),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_409),
.B(n_4),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_327),
.Y(n_501)
);

OA21x2_ASAP7_75t_L g502 ( 
.A1(n_321),
.A2(n_5),
.B(n_6),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_404),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_424),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_370),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_342),
.B(n_7),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_368),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_434),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_373),
.B(n_9),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_370),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_373),
.B(n_11),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_343),
.B(n_11),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_401),
.B(n_12),
.Y(n_514)
);

CKINVDCx6p67_ASAP7_75t_R g515 ( 
.A(n_376),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_343),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_453),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_316),
.B(n_15),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_336),
.B(n_15),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_375),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_465),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_353),
.B(n_16),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_380),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_353),
.B(n_17),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_375),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_372),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_450),
.B(n_18),
.Y(n_527)
);

AND2x2_ASAP7_75t_SL g528 ( 
.A(n_429),
.B(n_18),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_338),
.B(n_19),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_394),
.B(n_20),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_372),
.Y(n_531)
);

BUFx12f_ASAP7_75t_L g532 ( 
.A(n_385),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_392),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_398),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_375),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_386),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_412),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_516),
.B(n_378),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_469),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_472),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_482),
.B(n_427),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_475),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_493),
.B(n_341),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_471),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_516),
.B(n_386),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_501),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_481),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_501),
.Y(n_549)
);

CKINVDCx6p67_ASAP7_75t_R g550 ( 
.A(n_515),
.Y(n_550)
);

CKINVDCx6p67_ASAP7_75t_R g551 ( 
.A(n_532),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_510),
.B(n_512),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_L g553 ( 
.A(n_487),
.B(n_375),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_528),
.B(n_433),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_485),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_528),
.A2(n_439),
.B1(n_445),
.B2(n_452),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_486),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_473),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_488),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_473),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_474),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_474),
.Y(n_562)
);

AND2x6_ASAP7_75t_L g563 ( 
.A(n_507),
.B(n_393),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_489),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_476),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_478),
.B(n_441),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_L g567 ( 
.A1(n_508),
.A2(n_384),
.B1(n_411),
.B2(n_379),
.Y(n_567)
);

INVx6_ASAP7_75t_L g568 ( 
.A(n_525),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_476),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_476),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_480),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_496),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_526),
.B(n_410),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_468),
.B(n_410),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_470),
.B(n_444),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_531),
.B(n_428),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_478),
.B(n_385),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_536),
.B(n_428),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_490),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_490),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_491),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_491),
.Y(n_584)
);

NOR2x1p5_ASAP7_75t_L g585 ( 
.A(n_470),
.B(n_395),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_552),
.B(n_520),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_543),
.A2(n_502),
.B1(n_495),
.B2(n_468),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_547),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_556),
.B(n_512),
.C(n_510),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_566),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_576),
.B(n_520),
.Y(n_591)
);

NOR2xp67_ASAP7_75t_L g592 ( 
.A(n_549),
.B(n_520),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_541),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_548),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_525),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_539),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_576),
.B(n_477),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_550),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_556),
.B(n_566),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_579),
.B(n_514),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_568),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_558),
.B(n_477),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_560),
.Y(n_603)
);

AND2x6_ASAP7_75t_SL g604 ( 
.A(n_543),
.B(n_493),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_557),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_543),
.B(n_479),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_559),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_562),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_579),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_554),
.B(n_527),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_545),
.B(n_484),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_564),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_538),
.B(n_484),
.Y(n_614)
);

NOR3x1_ASAP7_75t_L g615 ( 
.A(n_554),
.B(n_500),
.C(n_518),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_585),
.B(n_500),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_569),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_575),
.B(n_418),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_573),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_574),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_539),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_567),
.A2(n_508),
.B1(n_483),
.B2(n_518),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_569),
.B(n_513),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_578),
.A2(n_530),
.B(n_483),
.C(n_529),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_570),
.B(n_513),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_553),
.A2(n_502),
.B1(n_495),
.B2(n_522),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_570),
.B(n_522),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_568),
.B(n_519),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_580),
.B(n_499),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_567),
.B(n_393),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_571),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_540),
.B(n_393),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_561),
.Y(n_633)
);

AND2x6_ASAP7_75t_SL g634 ( 
.A(n_551),
.B(n_530),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_581),
.B(n_524),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_581),
.B(n_491),
.Y(n_636)
);

AND2x6_ASAP7_75t_SL g637 ( 
.A(n_551),
.B(n_357),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_582),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_553),
.A2(n_519),
.B1(n_529),
.B2(n_499),
.Y(n_639)
);

O2A1O1Ixp5_ASAP7_75t_L g640 ( 
.A1(n_542),
.A2(n_505),
.B(n_509),
.C(n_504),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_584),
.B(n_506),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_546),
.B(n_523),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_544),
.B(n_568),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_572),
.B(n_506),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_572),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_542),
.A2(n_357),
.B1(n_419),
.B2(n_329),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_561),
.B(n_393),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_561),
.B(n_523),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_595),
.A2(n_565),
.B(n_561),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_598),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_597),
.A2(n_591),
.B(n_602),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_590),
.B(n_467),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_648),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_589),
.A2(n_497),
.B(n_323),
.C(n_332),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_594),
.B(n_503),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_605),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_590),
.A2(n_396),
.B1(n_455),
.B2(n_344),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_593),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_610),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_596),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_623),
.A2(n_583),
.B(n_535),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_606),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_628),
.B(n_563),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_608),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_611),
.A2(n_563),
.B1(n_492),
.B2(n_440),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_625),
.A2(n_583),
.B(n_535),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_627),
.A2(n_583),
.B(n_535),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_628),
.B(n_612),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_612),
.B(n_467),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_596),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_635),
.A2(n_511),
.B(n_430),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_607),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_624),
.A2(n_333),
.B(n_334),
.C(n_325),
.Y(n_673)
);

O2A1O1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_624),
.A2(n_630),
.B(n_611),
.C(n_600),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_587),
.A2(n_563),
.B(n_340),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_614),
.B(n_563),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_614),
.B(n_600),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_613),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_588),
.A2(n_419),
.B1(n_466),
.B2(n_461),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_621),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_630),
.A2(n_521),
.B(n_517),
.C(n_533),
.Y(n_681)
);

BUFx4_ASAP7_75t_SL g682 ( 
.A(n_637),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_587),
.A2(n_354),
.B1(n_355),
.B2(n_350),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_626),
.B(n_356),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_643),
.A2(n_359),
.B(n_358),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_626),
.A2(n_362),
.B(n_361),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_619),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_646),
.B(n_337),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_620),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_639),
.B(n_387),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_632),
.A2(n_391),
.B(n_389),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_615),
.B(n_405),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_632),
.A2(n_413),
.B(n_407),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_642),
.Y(n_694)
);

OR2x6_ASAP7_75t_SL g695 ( 
.A(n_622),
.B(n_339),
.Y(n_695)
);

BUFx12f_ASAP7_75t_L g696 ( 
.A(n_604),
.Y(n_696)
);

NOR2x1_ASAP7_75t_L g697 ( 
.A(n_616),
.B(n_422),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_640),
.A2(n_425),
.B(n_426),
.C(n_423),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_636),
.A2(n_436),
.B(n_432),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_618),
.B(n_534),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_622),
.A2(n_537),
.B(n_438),
.C(n_442),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_640),
.A2(n_446),
.B(n_447),
.C(n_437),
.Y(n_702)
);

BUFx12f_ASAP7_75t_L g703 ( 
.A(n_634),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_SL g704 ( 
.A(n_618),
.B(n_443),
.C(n_351),
.Y(n_704)
);

NOR2x1_ASAP7_75t_L g705 ( 
.A(n_592),
.B(n_451),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_631),
.A2(n_462),
.B(n_463),
.C(n_458),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_645),
.Y(n_707)
);

A2O1A1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_638),
.A2(n_319),
.B(n_326),
.C(n_317),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_644),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_603),
.B(n_347),
.Y(n_710)
);

OR2x6_ASAP7_75t_SL g711 ( 
.A(n_609),
.B(n_360),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_617),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_647),
.A2(n_403),
.B1(n_365),
.B2(n_397),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_647),
.A2(n_403),
.B1(n_406),
.B2(n_363),
.Y(n_714)
);

OA22x2_ASAP7_75t_L g715 ( 
.A1(n_641),
.A2(n_454),
.B1(n_460),
.B2(n_435),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_SL g716 ( 
.A1(n_633),
.A2(n_498),
.B(n_403),
.C(n_464),
.Y(n_716)
);

NAND2x1_ASAP7_75t_L g717 ( 
.A(n_626),
.B(n_498),
.Y(n_717)
);

INVx4_ASAP7_75t_L g718 ( 
.A(n_601),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_599),
.A2(n_346),
.B(n_348),
.C(n_345),
.Y(n_719)
);

AOI22x1_ASAP7_75t_L g720 ( 
.A1(n_610),
.A2(n_371),
.B1(n_381),
.B2(n_352),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_629),
.B(n_382),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_596),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_588),
.B(n_109),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_593),
.Y(n_724)
);

A2O1A1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_589),
.A2(n_388),
.B(n_390),
.C(n_383),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_589),
.A2(n_456),
.B1(n_400),
.B2(n_402),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_590),
.A2(n_416),
.B1(n_417),
.B2(n_415),
.Y(n_727)
);

BUFx8_ASAP7_75t_L g728 ( 
.A(n_593),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_595),
.A2(n_421),
.B(n_420),
.Y(n_729)
);

OAI21xp5_ASAP7_75t_L g730 ( 
.A1(n_586),
.A2(n_449),
.B(n_448),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_628),
.B(n_112),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_589),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_732)
);

BUFx4f_ASAP7_75t_L g733 ( 
.A(n_616),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_599),
.A2(n_24),
.B(n_21),
.C(n_23),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_593),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_590),
.A2(n_118),
.B1(n_119),
.B2(n_117),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_610),
.B(n_23),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_656),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_660),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_660),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_L g741 ( 
.A1(n_684),
.A2(n_121),
.B(n_120),
.Y(n_741)
);

INVx6_ASAP7_75t_L g742 ( 
.A(n_728),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_664),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_668),
.A2(n_127),
.B1(n_128),
.B2(n_125),
.Y(n_744)
);

AOI21x1_ASAP7_75t_L g745 ( 
.A1(n_663),
.A2(n_130),
.B(n_129),
.Y(n_745)
);

AO31x2_ASAP7_75t_L g746 ( 
.A1(n_654),
.A2(n_673),
.A3(n_686),
.B(n_698),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_651),
.A2(n_649),
.B(n_717),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_683),
.B(n_26),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_687),
.Y(n_749)
);

AOI31xp67_ASAP7_75t_L g750 ( 
.A1(n_692),
.A2(n_670),
.A3(n_722),
.B(n_680),
.Y(n_750)
);

AO31x2_ASAP7_75t_L g751 ( 
.A1(n_702),
.A2(n_31),
.A3(n_28),
.B(n_29),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_689),
.Y(n_752)
);

INVx6_ASAP7_75t_SL g753 ( 
.A(n_700),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_675),
.A2(n_135),
.B(n_134),
.Y(n_754)
);

NAND3x1_ASAP7_75t_L g755 ( 
.A(n_669),
.B(n_679),
.C(n_688),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_653),
.B(n_136),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_657),
.B(n_28),
.C(n_31),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_676),
.A2(n_140),
.B(n_138),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_658),
.Y(n_759)
);

AO32x2_ASAP7_75t_L g760 ( 
.A1(n_726),
.A2(n_701),
.A3(n_690),
.B1(n_734),
.B2(n_695),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_721),
.B(n_32),
.Y(n_761)
);

AO32x2_ASAP7_75t_L g762 ( 
.A1(n_718),
.A2(n_36),
.A3(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_719),
.A2(n_146),
.B(n_145),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_724),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_662),
.Y(n_765)
);

O2A1O1Ixp5_ASAP7_75t_L g766 ( 
.A1(n_730),
.A2(n_151),
.B(n_153),
.C(n_149),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_655),
.Y(n_767)
);

BUFx4f_ASAP7_75t_L g768 ( 
.A(n_696),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_709),
.B(n_37),
.Y(n_769)
);

AND2x2_ASAP7_75t_SL g770 ( 
.A(n_733),
.B(n_38),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_L g771 ( 
.A(n_665),
.B(n_39),
.C(n_40),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_650),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_655),
.B(n_154),
.Y(n_773)
);

NAND3x1_ASAP7_75t_L g774 ( 
.A(n_697),
.B(n_41),
.C(n_42),
.Y(n_774)
);

AO31x2_ASAP7_75t_L g775 ( 
.A1(n_725),
.A2(n_45),
.A3(n_43),
.B(n_44),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_672),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_661),
.A2(n_667),
.B(n_666),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_678),
.B(n_46),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_694),
.B(n_46),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_712),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_707),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_SL g782 ( 
.A(n_659),
.B(n_47),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_685),
.A2(n_158),
.B(n_156),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_710),
.B(n_48),
.Y(n_784)
);

NOR2x1_ASAP7_75t_SL g785 ( 
.A(n_700),
.B(n_159),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_681),
.Y(n_786)
);

AO31x2_ASAP7_75t_L g787 ( 
.A1(n_732),
.A2(n_50),
.A3(n_48),
.B(n_49),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_735),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_733),
.B(n_165),
.Y(n_789)
);

OR2x6_ASAP7_75t_SL g790 ( 
.A(n_682),
.B(n_49),
.Y(n_790)
);

OR2x6_ASAP7_75t_L g791 ( 
.A(n_703),
.B(n_51),
.Y(n_791)
);

AO31x2_ASAP7_75t_L g792 ( 
.A1(n_708),
.A2(n_58),
.A3(n_55),
.B(n_57),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_737),
.Y(n_793)
);

OAI21xp33_ASAP7_75t_L g794 ( 
.A1(n_652),
.A2(n_55),
.B(n_57),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_723),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_727),
.B(n_58),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_729),
.A2(n_169),
.B(n_168),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_713),
.B(n_59),
.Y(n_798)
);

BUFx4f_ASAP7_75t_SL g799 ( 
.A(n_728),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_714),
.B(n_59),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_720),
.B(n_60),
.Y(n_801)
);

CKINVDCx6p67_ASAP7_75t_R g802 ( 
.A(n_711),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_705),
.B(n_736),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_715),
.Y(n_804)
);

AOI221x1_ASAP7_75t_L g805 ( 
.A1(n_704),
.A2(n_225),
.B1(n_313),
.B2(n_312),
.C(n_311),
.Y(n_805)
);

AO31x2_ASAP7_75t_L g806 ( 
.A1(n_706),
.A2(n_62),
.A3(n_60),
.B(n_61),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_691),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_716),
.Y(n_808)
);

AO22x1_ASAP7_75t_L g809 ( 
.A1(n_693),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_809)
);

NOR4xp25_ASAP7_75t_L g810 ( 
.A(n_699),
.B(n_67),
.C(n_68),
.D(n_69),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_671),
.B(n_68),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_656),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_684),
.A2(n_174),
.B(n_173),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_668),
.B(n_69),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_662),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_658),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_660),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_668),
.B(n_70),
.Y(n_818)
);

OAI21x1_ASAP7_75t_SL g819 ( 
.A1(n_674),
.A2(n_176),
.B(n_175),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_683),
.B(n_177),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_668),
.B(n_70),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_656),
.Y(n_822)
);

AOI21x1_ASAP7_75t_L g823 ( 
.A1(n_663),
.A2(n_179),
.B(n_178),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_653),
.B(n_180),
.Y(n_824)
);

NAND2x1_ASAP7_75t_SL g825 ( 
.A(n_679),
.B(n_71),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_658),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_668),
.B(n_71),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_656),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_668),
.B(n_73),
.Y(n_829)
);

O2A1O1Ixp5_ASAP7_75t_SL g830 ( 
.A1(n_730),
.A2(n_73),
.B(n_74),
.C(n_77),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_684),
.A2(n_185),
.B(n_183),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_668),
.B(n_77),
.Y(n_832)
);

OAI21x1_ASAP7_75t_SL g833 ( 
.A1(n_674),
.A2(n_188),
.B(n_187),
.Y(n_833)
);

XOR2xp5_ASAP7_75t_L g834 ( 
.A(n_650),
.B(n_193),
.Y(n_834)
);

AOI211x1_ASAP7_75t_L g835 ( 
.A1(n_692),
.A2(n_78),
.B(n_79),
.C(n_80),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_656),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_658),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_658),
.Y(n_838)
);

AOI221x1_ASAP7_75t_L g839 ( 
.A1(n_673),
.A2(n_244),
.B1(n_310),
.B2(n_309),
.C(n_308),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_684),
.A2(n_199),
.B(n_198),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_668),
.B(n_80),
.Y(n_841)
);

AO21x1_ASAP7_75t_L g842 ( 
.A1(n_677),
.A2(n_81),
.B(n_83),
.Y(n_842)
);

AO31x2_ASAP7_75t_L g843 ( 
.A1(n_654),
.A2(n_83),
.A3(n_84),
.B(n_85),
.Y(n_843)
);

AO31x2_ASAP7_75t_L g844 ( 
.A1(n_654),
.A2(n_85),
.A3(n_86),
.B(n_87),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_658),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_660),
.Y(n_846)
);

OAI21x1_ASAP7_75t_SL g847 ( 
.A1(n_674),
.A2(n_246),
.B(n_307),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_668),
.B(n_88),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_658),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_668),
.B(n_89),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_658),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_660),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_684),
.A2(n_248),
.B(n_305),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_653),
.B(n_202),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_684),
.A2(n_249),
.B(n_304),
.Y(n_855)
);

AOI211x1_ASAP7_75t_L g856 ( 
.A1(n_692),
.A2(n_90),
.B(n_91),
.C(n_93),
.Y(n_856)
);

OA21x2_ASAP7_75t_L g857 ( 
.A1(n_747),
.A2(n_245),
.B(n_302),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_763),
.A2(n_813),
.B(n_741),
.Y(n_858)
);

OA21x2_ASAP7_75t_L g859 ( 
.A1(n_831),
.A2(n_853),
.B(n_840),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_739),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_814),
.B(n_90),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_767),
.B(n_203),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_829),
.B(n_94),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_SL g864 ( 
.A1(n_770),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_864)
);

NAND2x1p5_ASAP7_75t_L g865 ( 
.A(n_765),
.B(n_204),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_761),
.B(n_96),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_772),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_765),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_740),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_816),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_817),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_816),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_815),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_846),
.Y(n_874)
);

INVxp33_ASAP7_75t_L g875 ( 
.A(n_837),
.Y(n_875)
);

XOR2xp5_ASAP7_75t_L g876 ( 
.A(n_834),
.B(n_205),
.Y(n_876)
);

AO31x2_ASAP7_75t_L g877 ( 
.A1(n_839),
.A2(n_97),
.A3(n_98),
.B(n_99),
.Y(n_877)
);

OAI21xp33_ASAP7_75t_SL g878 ( 
.A1(n_841),
.A2(n_97),
.B(n_99),
.Y(n_878)
);

NOR2xp67_ASAP7_75t_L g879 ( 
.A(n_795),
.B(n_784),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_850),
.B(n_100),
.Y(n_880)
);

AOI22x1_ASAP7_75t_L g881 ( 
.A1(n_808),
.A2(n_252),
.B1(n_301),
.B2(n_298),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_852),
.Y(n_882)
);

AO21x2_ASAP7_75t_L g883 ( 
.A1(n_855),
.A2(n_241),
.B(n_295),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_738),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_743),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_749),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_752),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_826),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_786),
.A2(n_240),
.B(n_294),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_826),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_776),
.B(n_838),
.Y(n_891)
);

AO21x1_ASAP7_75t_L g892 ( 
.A1(n_754),
.A2(n_100),
.B(n_101),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_812),
.Y(n_893)
);

OAI21x1_ASAP7_75t_SL g894 ( 
.A1(n_785),
.A2(n_237),
.B(n_290),
.Y(n_894)
);

AO21x2_ASAP7_75t_L g895 ( 
.A1(n_758),
.A2(n_235),
.B(n_288),
.Y(n_895)
);

NOR2x1_ASAP7_75t_SL g896 ( 
.A(n_789),
.B(n_306),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_773),
.Y(n_897)
);

OAI21x1_ASAP7_75t_SL g898 ( 
.A1(n_819),
.A2(n_234),
.B(n_285),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_759),
.B(n_233),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_849),
.B(n_101),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_851),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_821),
.B(n_102),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_851),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_822),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_828),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_788),
.B(n_102),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_773),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_827),
.B(n_103),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_836),
.Y(n_909)
);

AO21x2_ASAP7_75t_L g910 ( 
.A1(n_833),
.A2(n_232),
.B(n_206),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_799),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_845),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_781),
.Y(n_913)
);

AO21x1_ASAP7_75t_L g914 ( 
.A1(n_832),
.A2(n_103),
.B(n_207),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_750),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_764),
.B(n_213),
.Y(n_916)
);

INVx8_ASAP7_75t_L g917 ( 
.A(n_756),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_745),
.A2(n_216),
.B(n_218),
.Y(n_918)
);

AO21x2_ASAP7_75t_L g919 ( 
.A1(n_847),
.A2(n_222),
.B(n_223),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_779),
.Y(n_920)
);

AOI21x1_ASAP7_75t_L g921 ( 
.A1(n_823),
.A2(n_224),
.B(n_226),
.Y(n_921)
);

OA21x2_ASAP7_75t_L g922 ( 
.A1(n_766),
.A2(n_227),
.B(n_228),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_843),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_848),
.A2(n_253),
.B(n_257),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_742),
.B(n_258),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_843),
.Y(n_926)
);

AO21x2_ASAP7_75t_L g927 ( 
.A1(n_797),
.A2(n_259),
.B(n_260),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_844),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_793),
.B(n_264),
.Y(n_929)
);

AO31x2_ASAP7_75t_L g930 ( 
.A1(n_842),
.A2(n_265),
.A3(n_266),
.B(n_269),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_787),
.Y(n_931)
);

AO21x2_ASAP7_75t_L g932 ( 
.A1(n_783),
.A2(n_270),
.B(n_272),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_756),
.B(n_286),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_753),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_811),
.Y(n_935)
);

OA21x2_ASAP7_75t_L g936 ( 
.A1(n_805),
.A2(n_274),
.B(n_276),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_780),
.B(n_769),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_751),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_751),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_746),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_804),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_804),
.B(n_796),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_824),
.Y(n_943)
);

AOI21xp33_ASAP7_75t_SL g944 ( 
.A1(n_757),
.A2(n_794),
.B(n_798),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_807),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_824),
.B(n_854),
.Y(n_946)
);

OA21x2_ASAP7_75t_L g947 ( 
.A1(n_778),
.A2(n_801),
.B(n_748),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_746),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_800),
.A2(n_820),
.B1(n_803),
.B2(n_854),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_775),
.Y(n_950)
);

INVx8_ASAP7_75t_L g951 ( 
.A(n_803),
.Y(n_951)
);

NOR2xp67_ASAP7_75t_L g952 ( 
.A(n_771),
.B(n_744),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_760),
.B(n_802),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_830),
.A2(n_755),
.B(n_774),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_825),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_760),
.A2(n_792),
.B(n_753),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_782),
.B(n_856),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_806),
.A2(n_809),
.B(n_810),
.Y(n_958)
);

INVx6_ASAP7_75t_L g959 ( 
.A(n_742),
.Y(n_959)
);

OAI21x1_ASAP7_75t_SL g960 ( 
.A1(n_762),
.A2(n_835),
.B(n_806),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_791),
.B(n_790),
.Y(n_961)
);

OA21x2_ASAP7_75t_L g962 ( 
.A1(n_762),
.A2(n_791),
.B(n_768),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_762),
.A2(n_747),
.B(n_777),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_761),
.B(n_629),
.Y(n_964)
);

AO21x2_ASAP7_75t_L g965 ( 
.A1(n_763),
.A2(n_731),
.B(n_741),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_772),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_818),
.A2(n_668),
.B(n_677),
.C(n_599),
.Y(n_967)
);

BUFx12f_ASAP7_75t_L g968 ( 
.A(n_742),
.Y(n_968)
);

NOR2x1_ASAP7_75t_SL g969 ( 
.A(n_765),
.B(n_789),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_816),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_816),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_739),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_765),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_816),
.Y(n_974)
);

NOR2x1_ASAP7_75t_SL g975 ( 
.A(n_765),
.B(n_789),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_739),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_814),
.B(n_668),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_765),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_739),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_814),
.B(n_668),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_765),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_765),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_970),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_977),
.B(n_980),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_971),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_888),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_884),
.Y(n_987)
);

AO21x2_ASAP7_75t_L g988 ( 
.A1(n_858),
.A2(n_965),
.B(n_915),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_964),
.B(n_946),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_967),
.A2(n_963),
.B(n_952),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_884),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_920),
.B(n_870),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_966),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_901),
.B(n_903),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_885),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_885),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_886),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_891),
.B(n_942),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_893),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_887),
.Y(n_1000)
);

AO21x2_ASAP7_75t_L g1001 ( 
.A1(n_858),
.A2(n_965),
.B(n_915),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_887),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_904),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_904),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_905),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_905),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_909),
.Y(n_1007)
);

NAND2x1p5_ASAP7_75t_L g1008 ( 
.A(n_981),
.B(n_907),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_872),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_968),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_941),
.B(n_866),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_SL g1012 ( 
.A(n_945),
.B(n_935),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_912),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_940),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_940),
.Y(n_1015)
);

BUFx2_ASAP7_75t_SL g1016 ( 
.A(n_867),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_890),
.B(n_974),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_959),
.Y(n_1018)
);

BUFx4f_ASAP7_75t_L g1019 ( 
.A(n_959),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_897),
.B(n_943),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_948),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_868),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_935),
.B(n_949),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_981),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_913),
.B(n_875),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_981),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_860),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_869),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_907),
.B(n_944),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_868),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_911),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_868),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_951),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_952),
.A2(n_859),
.B(n_948),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_951),
.B(n_917),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_871),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_882),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_944),
.B(n_937),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_897),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_978),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_972),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_938),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_976),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_978),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_973),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_979),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_939),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_861),
.B(n_863),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_859),
.A2(n_954),
.B(n_956),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_874),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_874),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_917),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_934),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_880),
.B(n_902),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_931),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_864),
.A2(n_892),
.B1(n_962),
.B2(n_914),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_908),
.B(n_955),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_862),
.B(n_982),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_900),
.B(n_906),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_916),
.B(n_953),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_873),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_925),
.B(n_876),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_925),
.B(n_879),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_923),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_899),
.Y(n_1065)
);

INVxp67_ASAP7_75t_SL g1066 ( 
.A(n_926),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_928),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_929),
.B(n_947),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_950),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_865),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_958),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_957),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_960),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_933),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_969),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_998),
.B(n_878),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_987),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_989),
.B(n_962),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_991),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_1014),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1059),
.B(n_1060),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_1066),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1011),
.B(n_975),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_984),
.B(n_961),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1057),
.B(n_930),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1054),
.B(n_930),
.Y(n_1086)
);

AND2x4_ASAP7_75t_SL g1087 ( 
.A(n_993),
.B(n_896),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1038),
.A2(n_924),
.B1(n_927),
.B2(n_883),
.Y(n_1088)
);

NOR4xp25_ASAP7_75t_SL g1089 ( 
.A(n_1072),
.B(n_936),
.C(n_877),
.D(n_927),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1048),
.B(n_930),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1038),
.A2(n_883),
.B1(n_932),
.B2(n_895),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_995),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_996),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_994),
.B(n_877),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1000),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1015),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1002),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1003),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1021),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1058),
.B(n_910),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1063),
.B(n_910),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1004),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_997),
.B(n_919),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_999),
.B(n_919),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_983),
.B(n_895),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1005),
.Y(n_1106)
);

AND2x4_ASAP7_75t_SL g1107 ( 
.A(n_993),
.B(n_898),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_983),
.B(n_932),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_985),
.B(n_918),
.Y(n_1109)
);

INVxp67_ASAP7_75t_SL g1110 ( 
.A(n_1066),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1006),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_985),
.B(n_921),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_1035),
.B(n_894),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1035),
.B(n_889),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1013),
.B(n_922),
.Y(n_1115)
);

INVx4_ASAP7_75t_R g1116 ( 
.A(n_1018),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1013),
.B(n_922),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_992),
.B(n_857),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_1017),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1007),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1025),
.B(n_881),
.Y(n_1121)
);

INVxp67_ASAP7_75t_SL g1122 ( 
.A(n_1042),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1035),
.B(n_1033),
.Y(n_1123)
);

BUFx2_ASAP7_75t_SL g1124 ( 
.A(n_986),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1074),
.B(n_1023),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1027),
.B(n_1028),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_1052),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_1032),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1061),
.Y(n_1129)
);

OAI21xp33_ASAP7_75t_SL g1130 ( 
.A1(n_1029),
.A2(n_1056),
.B(n_1075),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1032),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_1040),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1047),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1056),
.A2(n_1029),
.B1(n_1065),
.B2(n_990),
.Y(n_1134)
);

AO22x1_ASAP7_75t_L g1135 ( 
.A1(n_1065),
.A2(n_1070),
.B1(n_1062),
.B2(n_1020),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1064),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1016),
.B(n_1036),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1041),
.B(n_1037),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1012),
.B(n_1068),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1052),
.B(n_1039),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_1052),
.B(n_1039),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1055),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1078),
.B(n_1073),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_1129),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1125),
.B(n_1046),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1125),
.B(n_1043),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1142),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1086),
.B(n_1049),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1080),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1080),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1119),
.B(n_1070),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1119),
.B(n_1068),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1099),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1099),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_1094),
.B(n_988),
.Y(n_1155)
);

OR2x2_ASAP7_75t_L g1156 ( 
.A(n_1139),
.B(n_988),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1090),
.B(n_1067),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1082),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_1082),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1110),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1110),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1085),
.B(n_1108),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1084),
.B(n_1081),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1130),
.B(n_1051),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1131),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1105),
.B(n_1069),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1077),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1076),
.B(n_1050),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1079),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1092),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1093),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1095),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1096),
.B(n_1034),
.Y(n_1173)
);

OR2x2_ASAP7_75t_L g1174 ( 
.A(n_1139),
.B(n_1001),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1097),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1128),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1138),
.B(n_1126),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1128),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1098),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1083),
.B(n_1009),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1102),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1106),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1132),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1137),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_1118),
.B(n_1001),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1111),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1120),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1162),
.B(n_1071),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1147),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1162),
.B(n_1101),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1152),
.B(n_1122),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1180),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1166),
.B(n_1100),
.Y(n_1193)
);

AND2x4_ASAP7_75t_SL g1194 ( 
.A(n_1144),
.B(n_1123),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1167),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1169),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1170),
.Y(n_1197)
);

NAND5xp2_ASAP7_75t_L g1198 ( 
.A(n_1164),
.B(n_1088),
.C(n_1134),
.D(n_1091),
.E(n_990),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1171),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1166),
.B(n_1109),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1172),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1184),
.B(n_1112),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1164),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1175),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1155),
.B(n_1115),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1158),
.B(n_1161),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1143),
.B(n_1134),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1179),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1143),
.B(n_1103),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1181),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1182),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1155),
.B(n_1117),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1186),
.Y(n_1213)
);

NAND2x1p5_ASAP7_75t_L g1214 ( 
.A(n_1158),
.B(n_1114),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1148),
.B(n_1133),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1159),
.B(n_1133),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1160),
.B(n_1136),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1187),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1149),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1148),
.B(n_1104),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1150),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1153),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1154),
.Y(n_1223)
);

NAND3xp33_ASAP7_75t_L g1224 ( 
.A(n_1203),
.B(n_1088),
.C(n_1121),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1220),
.B(n_1156),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1189),
.Y(n_1226)
);

OAI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1192),
.A2(n_1146),
.B1(n_1145),
.B2(n_1163),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1189),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1213),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1202),
.B(n_1165),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1203),
.A2(n_1113),
.B1(n_1107),
.B2(n_1087),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1213),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1190),
.B(n_1157),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1200),
.B(n_1174),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1205),
.B(n_1185),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1220),
.B(n_1174),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1212),
.B(n_1185),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1206),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1218),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1218),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1195),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1193),
.B(n_1157),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1209),
.B(n_1176),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1196),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1188),
.B(n_1215),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1197),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1188),
.B(n_1173),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1199),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1227),
.A2(n_1198),
.B(n_1151),
.C(n_1168),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1224),
.A2(n_1207),
.B1(n_1113),
.B2(n_1107),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1231),
.A2(n_1113),
.B1(n_1198),
.B2(n_1214),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1225),
.B(n_1191),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1230),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1225),
.B(n_1206),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1246),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1245),
.B(n_1236),
.Y(n_1256)
);

AO22x1_ASAP7_75t_L g1257 ( 
.A1(n_1238),
.A2(n_1201),
.B1(n_1210),
.B2(n_1211),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1243),
.Y(n_1258)
);

AOI222xp33_ASAP7_75t_L g1259 ( 
.A1(n_1227),
.A2(n_1177),
.B1(n_1135),
.B2(n_1204),
.C1(n_1208),
.C2(n_1191),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1233),
.B(n_1219),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1246),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1234),
.B(n_1221),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1238),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1242),
.B(n_1123),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1235),
.B(n_1053),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1251),
.A2(n_1114),
.B(n_1216),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1249),
.A2(n_1087),
.B(n_1248),
.C(n_1244),
.Y(n_1267)
);

AOI222xp33_ASAP7_75t_L g1268 ( 
.A1(n_1258),
.A2(n_1241),
.B1(n_1183),
.B2(n_1178),
.C1(n_1222),
.C2(n_1223),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1259),
.A2(n_1194),
.B1(n_1247),
.B2(n_1237),
.Y(n_1269)
);

OAI31xp33_ASAP7_75t_L g1270 ( 
.A1(n_1253),
.A2(n_1214),
.A3(n_1194),
.B(n_1239),
.Y(n_1270)
);

NOR2x1_ASAP7_75t_L g1271 ( 
.A(n_1261),
.B(n_1226),
.Y(n_1271)
);

AOI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1257),
.A2(n_1240),
.B(n_1232),
.Y(n_1272)
);

AOI211xp5_ASAP7_75t_L g1273 ( 
.A1(n_1267),
.A2(n_1265),
.B(n_1250),
.C(n_1264),
.Y(n_1273)
);

AOI21xp33_ASAP7_75t_L g1274 ( 
.A1(n_1269),
.A2(n_1263),
.B(n_1262),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1271),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1266),
.B(n_1010),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1270),
.A2(n_1260),
.B1(n_1252),
.B2(n_1255),
.C(n_1228),
.Y(n_1277)
);

OAI211xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1274),
.A2(n_1268),
.B(n_1255),
.C(n_1256),
.Y(n_1278)
);

NAND5xp2_ASAP7_75t_L g1279 ( 
.A(n_1276),
.B(n_1272),
.C(n_1254),
.D(n_1091),
.E(n_1008),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1277),
.B(n_1247),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_L g1281 ( 
.A(n_1275),
.B(n_1217),
.C(n_1216),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1273),
.B(n_1229),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1282),
.B(n_1281),
.C(n_1278),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_SL g1284 ( 
.A(n_1280),
.B(n_1031),
.C(n_1089),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1279),
.B(n_1053),
.Y(n_1285)
);

OAI211xp5_ASAP7_75t_L g1286 ( 
.A1(n_1283),
.A2(n_1284),
.B(n_1285),
.C(n_1031),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1283),
.B(n_1124),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1287),
.B(n_1229),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1288),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1289),
.A2(n_1286),
.B1(n_1019),
.B2(n_1127),
.Y(n_1290)
);

AO22x2_ASAP7_75t_L g1291 ( 
.A1(n_1290),
.A2(n_1026),
.B1(n_1024),
.B2(n_1116),
.Y(n_1291)
);

XNOR2x1_ASAP7_75t_L g1292 ( 
.A(n_1291),
.B(n_1019),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1292),
.B(n_1022),
.C(n_1045),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1293),
.A2(n_1044),
.B(n_1140),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1294),
.A2(n_1140),
.B1(n_1141),
.B2(n_1030),
.Y(n_1295)
);


endmodule