module fake_jpeg_4130_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_15),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_22),
.B1(n_11),
.B2(n_23),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_40),
.B1(n_14),
.B2(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_24),
.Y(n_50)
);

NAND2x1_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_18),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_19),
.C(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_16),
.B1(n_12),
.B2(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_16),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_27),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_17),
.B(n_20),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_12),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_53),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_54),
.B(n_56),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_55),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_34),
.B1(n_27),
.B2(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_71),
.B(n_78),
.Y(n_82)
);

OAI322xp33_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_41),
.A3(n_44),
.B1(n_43),
.B2(n_54),
.C1(n_48),
.C2(n_26),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_77),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_47),
.B(n_26),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_68),
.B(n_63),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_67),
.A3(n_68),
.B1(n_59),
.B2(n_60),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_62),
.B(n_64),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_53),
.B(n_17),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_52),
.C(n_17),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_75),
.B1(n_76),
.B2(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_82),
.B(n_7),
.Y(n_93)
);

FAx1_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_5),
.CI(n_10),
.CON(n_97),
.SN(n_97)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_87),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_1),
.B(n_2),
.Y(n_96)
);

NAND5xp2_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_88),
.C(n_8),
.D(n_5),
.E(n_9),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_97),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_4),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_4),
.C(n_100),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_99),
.B(n_4),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_99),
.Y(n_104)
);


endmodule