module fake_jpeg_23847_n_193 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_193);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_27),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_40),
.Y(n_77)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_1),
.C(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_32),
.B1(n_31),
.B2(n_5),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_2),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_3),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_64),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_17),
.B1(n_16),
.B2(n_22),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_54),
.B1(n_73),
.B2(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_27),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_31),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_65),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_69),
.C(n_6),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_31),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_31),
.B(n_26),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_3),
.B(n_4),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_75),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_35),
.A2(n_25),
.B1(n_29),
.B2(n_20),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_35),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_4),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_97),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_75),
.B(n_8),
.Y(n_109)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_12),
.A3(n_11),
.B1(n_10),
.B2(n_7),
.Y(n_90)
);

NOR4xp25_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_8),
.C(n_9),
.D(n_64),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_98),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_5),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_6),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_11),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_7),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_54),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_62),
.B(n_53),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_123),
.B1(n_102),
.B2(n_97),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_110),
.B1(n_100),
.B2(n_83),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_114),
.B(n_120),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_70),
.B1(n_63),
.B2(n_56),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_125),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_121),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_54),
.B(n_49),
.Y(n_120)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_95),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_138),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_79),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_134),
.Y(n_152)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_95),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_132),
.B(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_123),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_78),
.B(n_88),
.C(n_82),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_111),
.B1(n_93),
.B2(n_86),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_98),
.C(n_87),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_141),
.C(n_116),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_121),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_101),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_84),
.C(n_78),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_128),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_120),
.B(n_109),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_111),
.C(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_157),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_106),
.B1(n_105),
.B2(n_103),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_155),
.B1(n_122),
.B2(n_113),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_106),
.B1(n_105),
.B2(n_82),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_55),
.C(n_118),
.Y(n_157)
);

XOR2x1_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_129),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_152),
.C(n_148),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_134),
.B1(n_126),
.B2(n_135),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_160),
.A2(n_162),
.B1(n_122),
.B2(n_151),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_149),
.C(n_157),
.Y(n_171)
);

OAI322xp33_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_139),
.A3(n_132),
.B1(n_144),
.B2(n_141),
.C1(n_137),
.C2(n_140),
.Y(n_163)
);

AOI31xp33_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_166),
.A3(n_152),
.B(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_168),
.B1(n_72),
.B2(n_133),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_139),
.B1(n_126),
.B2(n_118),
.C(n_112),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_174),
.B(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_172),
.C(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_176),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_159),
.A2(n_133),
.B(n_72),
.C(n_64),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_156),
.C(n_92),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_72),
.C(n_8),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_162),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_164),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_187),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_178),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_189),
.B(n_181),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_170),
.B1(n_181),
.B2(n_171),
.Y(n_189)
);

HAxp5_ASAP7_75t_SL g193 ( 
.A(n_191),
.B(n_192),
.CON(n_193),
.SN(n_193)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_184),
.B(n_9),
.Y(n_192)
);


endmodule