module fake_netlist_1_418_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_30;
wire n_26;
wire n_16;
wire n_33;
wire n_13;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
INVx3_ASAP7_75t_L g10 ( .A(n_3), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_9), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_0), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_11), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_10), .B(n_1), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_10), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_10), .B(n_1), .Y(n_20) );
INVx3_ASAP7_75t_L g21 ( .A(n_10), .Y(n_21) );
BUFx3_ASAP7_75t_L g22 ( .A(n_12), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
CKINVDCx16_ASAP7_75t_R g25 ( .A(n_22), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_17), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_20), .B1(n_18), .B2(n_19), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_23), .A2(n_20), .B1(n_18), .B2(n_19), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_25), .B(n_20), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_26), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_29), .B(n_23), .Y(n_31) );
AOI22xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_20), .B1(n_28), .B2(n_27), .Y(n_32) );
INVx3_ASAP7_75t_SL g33 ( .A(n_31), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_31), .A2(n_22), .B(n_21), .Y(n_34) );
NAND3xp33_ASAP7_75t_SL g35 ( .A(n_32), .B(n_15), .C(n_14), .Y(n_35) );
NOR3xp33_ASAP7_75t_L g36 ( .A(n_34), .B(n_16), .C(n_21), .Y(n_36) );
OAI211xp5_ASAP7_75t_L g37 ( .A1(n_33), .A2(n_16), .B(n_21), .C(n_19), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_35), .B(n_21), .Y(n_38) );
AOI221xp5_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_21), .B1(n_19), .B2(n_22), .C(n_13), .Y(n_39) );
AOI22xp33_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_39), .B1(n_37), .B2(n_5), .Y(n_40) );
AOI22xp33_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_2), .B1(n_7), .B2(n_8), .Y(n_41) );
endmodule