module real_aes_6799_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g484 ( .A1(n_0), .A2(n_188), .B(n_485), .C(n_488), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_1), .B(n_479), .Y(n_490) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g237 ( .A(n_3), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_4), .B(n_176), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_5), .A2(n_463), .B(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g760 ( .A1(n_6), .A2(n_9), .B1(n_446), .B2(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_6), .Y(n_761) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_7), .A2(n_193), .B(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_8), .A2(n_39), .B1(n_149), .B2(n_161), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_9), .A2(n_133), .B1(n_134), .B2(n_446), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_9), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_10), .B(n_193), .Y(n_226) );
AND2x6_ASAP7_75t_L g164 ( .A(n_11), .B(n_165), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_12), .A2(n_164), .B(n_466), .C(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_13), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_14), .B(n_40), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_14), .B(n_40), .Y(n_123) );
INVx1_ASAP7_75t_L g145 ( .A(n_15), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_16), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g231 ( .A(n_17), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_18), .B(n_176), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_19), .B(n_191), .Y(n_209) );
AO32x2_ASAP7_75t_L g185 ( .A1(n_20), .A2(n_186), .A3(n_190), .B1(n_192), .B2(n_193), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_21), .A2(n_100), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_21), .Y(n_128) );
AND2x2_ASAP7_75t_L g527 ( .A(n_22), .B(n_141), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_23), .B(n_149), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_24), .B(n_191), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_25), .A2(n_55), .B1(n_149), .B2(n_161), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g202 ( .A1(n_26), .A2(n_81), .B1(n_149), .B2(n_153), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_27), .B(n_149), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_28), .A2(n_192), .B(n_466), .C(n_468), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_29), .A2(n_192), .B(n_466), .C(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_30), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_31), .B(n_141), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_32), .A2(n_463), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_33), .B(n_141), .Y(n_183) );
INVx2_ASAP7_75t_L g151 ( .A(n_34), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_35), .A2(n_497), .B(n_498), .C(n_502), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_36), .B(n_149), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_37), .B(n_141), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_38), .B(n_156), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_41), .B(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_42), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_43), .B(n_176), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_44), .B(n_463), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_45), .A2(n_497), .B(n_502), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_46), .B(n_149), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_47), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g486 ( .A(n_48), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_49), .A2(n_90), .B1(n_161), .B2(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g525 ( .A(n_50), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_51), .B(n_149), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_52), .B(n_149), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_53), .B(n_463), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_54), .B(n_224), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g213 ( .A1(n_56), .A2(n_60), .B1(n_149), .B2(n_153), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_57), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_58), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_59), .B(n_149), .Y(n_250) );
INVx1_ASAP7_75t_L g165 ( .A(n_61), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_62), .B(n_463), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_63), .B(n_479), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_64), .A2(n_224), .B(n_234), .C(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_65), .B(n_149), .Y(n_238) );
INVx1_ASAP7_75t_L g144 ( .A(n_66), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_67), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_68), .B(n_176), .Y(n_500) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_69), .A2(n_192), .A3(n_193), .B1(n_199), .B2(n_203), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_70), .B(n_177), .Y(n_556) );
INVx1_ASAP7_75t_L g249 ( .A(n_71), .Y(n_249) );
INVx1_ASAP7_75t_L g174 ( .A(n_72), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_73), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_74), .B(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_75), .A2(n_466), .B(n_502), .C(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_76), .B(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_76), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_77), .B(n_153), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_78), .Y(n_534) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_80), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_82), .B(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_83), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_84), .B(n_153), .Y(n_180) );
INVx2_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_86), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_87), .B(n_163), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_88), .B(n_153), .Y(n_220) );
INVx2_ASAP7_75t_L g112 ( .A(n_89), .Y(n_112) );
OR2x2_ASAP7_75t_L g120 ( .A(n_89), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g449 ( .A(n_89), .B(n_122), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_91), .A2(n_101), .B1(n_153), .B2(n_154), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_92), .B(n_463), .Y(n_495) );
INVx1_ASAP7_75t_L g499 ( .A(n_93), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_94), .A2(n_103), .B1(n_116), .B2(n_766), .Y(n_102) );
INVxp67_ASAP7_75t_L g537 ( .A(n_95), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_96), .B(n_153), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_97), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g512 ( .A(n_98), .Y(n_512) );
INVx1_ASAP7_75t_L g552 ( .A(n_99), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_100), .Y(n_127) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g766 ( .A(n_105), .Y(n_766) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .C(n_113), .Y(n_110) );
AND2x2_ASAP7_75t_L g122 ( .A(n_111), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g743 ( .A(n_112), .B(n_122), .Y(n_743) );
NOR2x2_ASAP7_75t_L g751 ( .A(n_112), .B(n_121), .Y(n_751) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_124), .Y(n_117) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g765 ( .A(n_120), .Y(n_765) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI32xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_748), .A3(n_752), .B1(n_753), .B2(n_756), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_744), .B2(n_745), .Y(n_125) );
INVx1_ASAP7_75t_L g744 ( .A(n_126), .Y(n_744) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22x1_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_447), .B1(n_450), .B2(n_741), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_132), .A2(n_451), .B1(n_741), .B2(n_747), .Y(n_746) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_133), .A2(n_134), .B1(n_759), .B2(n_760), .Y(n_758) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_368), .Y(n_134) );
NAND5xp2_ASAP7_75t_L g135 ( .A(n_136), .B(n_287), .C(n_302), .D(n_328), .E(n_350), .Y(n_135) );
NOR2xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_267), .Y(n_136) );
OAI221xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_204), .B1(n_240), .B2(n_256), .C(n_257), .Y(n_137) );
NOR2xp33_ASAP7_75t_SL g138 ( .A(n_139), .B(n_194), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_139), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g444 ( .A(n_139), .Y(n_444) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_167), .Y(n_139) );
INVx1_ASAP7_75t_L g284 ( .A(n_140), .Y(n_284) );
AND2x2_ASAP7_75t_L g286 ( .A(n_140), .B(n_185), .Y(n_286) );
AND2x2_ASAP7_75t_L g296 ( .A(n_140), .B(n_184), .Y(n_296) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_140), .Y(n_314) );
INVx1_ASAP7_75t_L g324 ( .A(n_140), .Y(n_324) );
OR2x2_ASAP7_75t_L g362 ( .A(n_140), .B(n_261), .Y(n_362) );
INVx2_ASAP7_75t_L g412 ( .A(n_140), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_140), .B(n_260), .Y(n_429) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_146), .B(n_166), .Y(n_140) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_141), .A2(n_171), .B(n_183), .Y(n_170) );
INVx2_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
INVx1_ASAP7_75t_L g476 ( .A(n_141), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_141), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_141), .A2(n_522), .B(n_523), .Y(n_521) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_L g191 ( .A(n_142), .B(n_143), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_158), .B(n_164), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_152), .B(n_155), .Y(n_147) );
INVx3_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_149), .Y(n_514) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
BUFx3_ASAP7_75t_L g201 ( .A(n_150), .Y(n_201) );
AND2x6_ASAP7_75t_L g466 ( .A(n_150), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
INVx1_ASAP7_75t_L g225 ( .A(n_151), .Y(n_225) );
INVx2_ASAP7_75t_L g232 ( .A(n_153), .Y(n_232) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_157), .Y(n_163) );
INVx3_ASAP7_75t_L g177 ( .A(n_157), .Y(n_177) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
AND2x2_ASAP7_75t_L g464 ( .A(n_157), .B(n_225), .Y(n_464) );
INVx1_ASAP7_75t_L g467 ( .A(n_157), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_162), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_L g248 ( .A1(n_162), .A2(n_236), .B(n_249), .C(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_163), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g199 ( .A1(n_163), .A2(n_177), .B1(n_200), .B2(n_202), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_163), .A2(n_188), .B1(n_212), .B2(n_213), .Y(n_211) );
INVx4_ASAP7_75t_L g487 ( .A(n_163), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_164), .A2(n_172), .B(n_178), .Y(n_171) );
BUFx3_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_164), .A2(n_218), .B(n_221), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_164), .A2(n_230), .B(n_235), .Y(n_229) );
AND2x4_ASAP7_75t_L g463 ( .A(n_164), .B(n_464), .Y(n_463) );
INVx4_ASAP7_75t_SL g489 ( .A(n_164), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g553 ( .A(n_164), .B(n_464), .Y(n_553) );
NOR2xp67_ASAP7_75t_L g167 ( .A(n_168), .B(n_184), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_169), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_169), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_169), .B(n_284), .Y(n_344) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_170), .Y(n_196) );
INVx2_ASAP7_75t_L g261 ( .A(n_170), .Y(n_261) );
OR2x2_ASAP7_75t_L g323 ( .A(n_170), .B(n_324), .Y(n_323) );
O2A1O1Ixp5_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_176), .Y(n_172) );
INVx2_ASAP7_75t_L g188 ( .A(n_176), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_176), .A2(n_219), .B(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_176), .A2(n_246), .B(n_247), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_176), .B(n_537), .Y(n_536) );
INVx5_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
INVx1_ASAP7_75t_L g234 ( .A(n_181), .Y(n_234) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g470 ( .A(n_182), .Y(n_470) );
AND2x2_ASAP7_75t_L g262 ( .A(n_184), .B(n_198), .Y(n_262) );
AND2x2_ASAP7_75t_L g279 ( .A(n_184), .B(n_259), .Y(n_279) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g197 ( .A(n_185), .B(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g282 ( .A(n_185), .Y(n_282) );
AND2x2_ASAP7_75t_L g411 ( .A(n_185), .B(n_412), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_188), .A2(n_222), .B(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_188), .A2(n_236), .B(n_237), .C(n_238), .Y(n_235) );
INVx2_ASAP7_75t_L g228 ( .A(n_190), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_190), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_191), .Y(n_193) );
NAND3xp33_ASAP7_75t_L g210 ( .A(n_192), .B(n_211), .C(n_214), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_192), .A2(n_245), .B(n_248), .Y(n_244) );
INVx4_ASAP7_75t_L g214 ( .A(n_193), .Y(n_214) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_193), .A2(n_217), .B(n_226), .Y(n_216) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_193), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_193), .A2(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g256 ( .A(n_194), .Y(n_256) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_197), .Y(n_194) );
AND2x2_ASAP7_75t_L g374 ( .A(n_195), .B(n_262), .Y(n_374) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g375 ( .A(n_196), .B(n_286), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g342 ( .A1(n_197), .A2(n_343), .B(n_345), .C(n_347), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_197), .B(n_343), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_197), .A2(n_273), .B1(n_416), .B2(n_417), .C(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g259 ( .A(n_198), .Y(n_259) );
INVx1_ASAP7_75t_L g295 ( .A(n_198), .Y(n_295) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_198), .Y(n_304) );
INVx2_ASAP7_75t_L g488 ( .A(n_201), .Y(n_488) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_201), .Y(n_501) );
INVx1_ASAP7_75t_L g473 ( .A(n_203), .Y(n_473) );
INVx1_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_215), .Y(n_205) );
AND2x2_ASAP7_75t_L g321 ( .A(n_206), .B(n_266), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_206), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_207), .B(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g413 ( .A(n_207), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g445 ( .A(n_207), .Y(n_445) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx3_ASAP7_75t_L g275 ( .A(n_208), .Y(n_275) );
AND2x2_ASAP7_75t_L g301 ( .A(n_208), .B(n_255), .Y(n_301) );
NOR2x1_ASAP7_75t_L g310 ( .A(n_208), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g317 ( .A(n_208), .B(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g253 ( .A(n_209), .Y(n_253) );
AO21x1_ASAP7_75t_L g252 ( .A1(n_211), .A2(n_214), .B(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g479 ( .A(n_214), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_214), .B(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_214), .A2(n_509), .B(n_516), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_214), .B(n_517), .Y(n_516) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_214), .A2(n_551), .B(n_558), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_215), .B(n_357), .Y(n_392) );
INVx1_ASAP7_75t_SL g396 ( .A(n_215), .Y(n_396) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_227), .Y(n_215) );
INVx3_ASAP7_75t_L g255 ( .A(n_216), .Y(n_255) );
AND2x2_ASAP7_75t_L g266 ( .A(n_216), .B(n_243), .Y(n_266) );
AND2x2_ASAP7_75t_L g288 ( .A(n_216), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g333 ( .A(n_216), .B(n_327), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_216), .B(n_265), .Y(n_414) );
INVx2_ASAP7_75t_L g236 ( .A(n_224), .Y(n_236) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g254 ( .A(n_227), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_227), .B(n_243), .Y(n_290) );
AND2x2_ASAP7_75t_L g326 ( .A(n_227), .B(n_327), .Y(n_326) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_239), .Y(n_227) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_228), .A2(n_244), .B(n_251), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .C(n_234), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_232), .A2(n_546), .B(n_547), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_232), .A2(n_556), .B(n_557), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_234), .A2(n_512), .B(n_513), .C(n_514), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_236), .A2(n_469), .B(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_254), .Y(n_241) );
INVx1_ASAP7_75t_L g306 ( .A(n_242), .Y(n_306) );
AND2x2_ASAP7_75t_L g348 ( .A(n_242), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_242), .B(n_269), .Y(n_354) );
AOI21xp5_ASAP7_75t_SL g428 ( .A1(n_242), .A2(n_260), .B(n_283), .Y(n_428) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_252), .Y(n_242) );
OR2x2_ASAP7_75t_L g271 ( .A(n_243), .B(n_252), .Y(n_271) );
AND2x2_ASAP7_75t_L g318 ( .A(n_243), .B(n_255), .Y(n_318) );
INVx2_ASAP7_75t_L g327 ( .A(n_243), .Y(n_327) );
INVx1_ASAP7_75t_L g433 ( .A(n_243), .Y(n_433) );
AND2x2_ASAP7_75t_L g357 ( .A(n_252), .B(n_327), .Y(n_357) );
INVx1_ASAP7_75t_L g382 ( .A(n_252), .Y(n_382) );
AND2x2_ASAP7_75t_L g291 ( .A(n_254), .B(n_275), .Y(n_291) );
AND2x2_ASAP7_75t_L g303 ( .A(n_254), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_SL g421 ( .A(n_254), .Y(n_421) );
INVx2_ASAP7_75t_L g311 ( .A(n_255), .Y(n_311) );
AND2x2_ASAP7_75t_L g349 ( .A(n_255), .B(n_265), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_255), .B(n_433), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_262), .B(n_263), .Y(n_257) );
AND2x2_ASAP7_75t_L g364 ( .A(n_258), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g418 ( .A(n_258), .Y(n_418) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g338 ( .A(n_259), .Y(n_338) );
BUFx2_ASAP7_75t_L g437 ( .A(n_259), .Y(n_437) );
BUFx2_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
AND2x2_ASAP7_75t_L g410 ( .A(n_260), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g393 ( .A(n_261), .Y(n_393) );
AND2x4_ASAP7_75t_L g320 ( .A(n_262), .B(n_283), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g356 ( .A(n_262), .B(n_344), .Y(n_356) );
AOI32xp33_ASAP7_75t_L g280 ( .A1(n_263), .A2(n_281), .A3(n_283), .B1(n_285), .B2(n_286), .Y(n_280) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
INVx3_ASAP7_75t_L g269 ( .A(n_264), .Y(n_269) );
OR2x2_ASAP7_75t_L g405 ( .A(n_264), .B(n_361), .Y(n_405) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g274 ( .A(n_265), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g381 ( .A(n_265), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g273 ( .A(n_266), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g285 ( .A(n_266), .B(n_275), .Y(n_285) );
INVx1_ASAP7_75t_L g406 ( .A(n_266), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_266), .B(n_381), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_272), .B(n_276), .C(n_280), .Y(n_267) );
OAI322xp33_ASAP7_75t_L g376 ( .A1(n_268), .A2(n_313), .A3(n_377), .B1(n_379), .B2(n_383), .C1(n_384), .C2(n_388), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVxp67_ASAP7_75t_L g341 ( .A(n_269), .Y(n_341) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g395 ( .A(n_271), .B(n_396), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_271), .B(n_311), .Y(n_442) );
INVxp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g334 ( .A(n_274), .Y(n_334) );
OR2x2_ASAP7_75t_L g420 ( .A(n_275), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_278), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g329 ( .A(n_279), .B(n_308), .Y(n_329) );
AND2x2_ASAP7_75t_L g400 ( .A(n_279), .B(n_313), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_279), .B(n_387), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g287 ( .A1(n_281), .A2(n_288), .B1(n_291), .B2(n_292), .C(n_297), .Y(n_287) );
OR2x2_ASAP7_75t_L g298 ( .A(n_281), .B(n_294), .Y(n_298) );
AND2x2_ASAP7_75t_L g386 ( .A(n_281), .B(n_387), .Y(n_386) );
AOI32xp33_ASAP7_75t_L g425 ( .A1(n_281), .A2(n_311), .A3(n_426), .B1(n_427), .B2(n_430), .Y(n_425) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_282), .B(n_318), .C(n_341), .Y(n_359) );
AND2x2_ASAP7_75t_L g385 ( .A(n_282), .B(n_378), .Y(n_385) );
INVxp67_ASAP7_75t_L g365 ( .A(n_283), .Y(n_365) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_286), .B(n_338), .Y(n_394) );
INVx2_ASAP7_75t_L g404 ( .A(n_286), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_286), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g373 ( .A(n_289), .Y(n_373) );
OR2x2_ASAP7_75t_L g299 ( .A(n_290), .B(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_292), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_295), .Y(n_378) );
AND2x2_ASAP7_75t_L g337 ( .A(n_296), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g383 ( .A(n_296), .Y(n_383) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_296), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AOI21xp33_ASAP7_75t_SL g322 ( .A1(n_298), .A2(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g416 ( .A(n_301), .B(n_326), .Y(n_416) );
AOI211xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_305), .B(n_315), .C(n_322), .Y(n_302) );
AND2x2_ASAP7_75t_L g346 ( .A(n_304), .B(n_314), .Y(n_346) );
INVx2_ASAP7_75t_L g361 ( .A(n_304), .Y(n_361) );
OR2x2_ASAP7_75t_L g399 ( .A(n_304), .B(n_362), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_304), .B(n_442), .Y(n_441) );
AOI211xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_307), .B(n_309), .C(n_312), .Y(n_305) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_308), .B(n_346), .Y(n_345) );
OAI211xp5_ASAP7_75t_L g427 ( .A1(n_309), .A2(n_404), .B(n_428), .C(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_310), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g367 ( .A(n_311), .B(n_357), .Y(n_367) );
INVx1_ASAP7_75t_L g372 ( .A(n_311), .Y(n_372) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_316), .B(n_319), .Y(n_315) );
INVxp33_ASAP7_75t_L g423 ( .A(n_317), .Y(n_423) );
AND2x2_ASAP7_75t_L g402 ( .A(n_318), .B(n_381), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_323), .A2(n_385), .B(n_386), .Y(n_384) );
OAI322xp33_ASAP7_75t_L g403 ( .A1(n_325), .A2(n_404), .A3(n_405), .B1(n_406), .B2(n_407), .C1(n_409), .C2(n_413), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B1(n_335), .B2(n_339), .C(n_342), .Y(n_328) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g380 ( .A(n_333), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g424 ( .A(n_337), .Y(n_424) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_340), .B(n_360), .Y(n_426) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g389 ( .A(n_349), .B(n_357), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B1(n_355), .B2(n_357), .C(n_358), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_353), .A2(n_370), .B1(n_374), .B2(n_375), .C(n_376), .Y(n_369) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_357), .B(n_372), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B1(n_363), .B2(n_366), .Y(n_358) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx2_ASAP7_75t_SL g387 ( .A(n_362), .Y(n_387) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND5xp2_ASAP7_75t_L g368 ( .A(n_369), .B(n_390), .C(n_415), .D(n_425), .E(n_435), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_371), .B(n_373), .Y(n_370) );
NOR4xp25_ASAP7_75t_L g443 ( .A(n_372), .B(n_378), .C(n_444), .D(n_445), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_375), .A2(n_436), .B1(n_438), .B2(n_440), .C(n_443), .Y(n_435) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
OAI322xp33_ASAP7_75t_L g391 ( .A1(n_385), .A2(n_392), .A3(n_393), .B1(n_394), .B2(n_395), .C1(n_397), .C2(n_401), .Y(n_391) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_403), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g436 ( .A(n_411), .B(n_437), .Y(n_436) );
OAI22xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B1(n_423), .B2(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g747 ( .A(n_448), .Y(n_747) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_696), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_631), .Y(n_452) );
NAND4xp25_ASAP7_75t_SL g453 ( .A(n_454), .B(n_576), .C(n_600), .D(n_623), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_518), .B1(n_548), .B2(n_560), .C(n_563), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_491), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_457), .A2(n_477), .B1(n_519), .B2(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_457), .B(n_492), .Y(n_634) );
AND2x2_ASAP7_75t_L g653 ( .A(n_457), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_457), .B(n_637), .Y(n_723) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_477), .Y(n_457) );
AND2x2_ASAP7_75t_L g591 ( .A(n_458), .B(n_492), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_458), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g614 ( .A(n_458), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g619 ( .A(n_458), .B(n_478), .Y(n_619) );
INVx2_ASAP7_75t_L g651 ( .A(n_458), .Y(n_651) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_458), .Y(n_695) );
AND2x2_ASAP7_75t_L g712 ( .A(n_458), .B(n_589), .Y(n_712) );
INVx5_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g630 ( .A(n_459), .B(n_589), .Y(n_630) );
AND2x4_ASAP7_75t_L g644 ( .A(n_459), .B(n_477), .Y(n_644) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_459), .Y(n_648) );
AND2x2_ASAP7_75t_L g668 ( .A(n_459), .B(n_583), .Y(n_668) );
AND2x2_ASAP7_75t_L g718 ( .A(n_459), .B(n_493), .Y(n_718) );
AND2x2_ASAP7_75t_L g728 ( .A(n_459), .B(n_478), .Y(n_728) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_474), .Y(n_459) );
AOI21xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_465), .B(n_473), .Y(n_460) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx5_ASAP7_75t_L g483 ( .A(n_466), .Y(n_483) );
INVx2_ASAP7_75t_L g472 ( .A(n_470), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_472), .A2(n_499), .B(n_500), .C(n_501), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_472), .A2(n_501), .B(n_525), .C(n_526), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AND2x2_ASAP7_75t_L g584 ( .A(n_477), .B(n_492), .Y(n_584) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_477), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_477), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g674 ( .A(n_477), .Y(n_674) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g562 ( .A(n_478), .B(n_507), .Y(n_562) );
AND2x2_ASAP7_75t_L g589 ( .A(n_478), .B(n_508), .Y(n_589) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_490), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_483), .B(n_484), .C(n_489), .Y(n_481) );
INVx2_ASAP7_75t_L g497 ( .A(n_483), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_483), .A2(n_489), .B(n_534), .C(n_535), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g502 ( .A(n_489), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_491), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_505), .Y(n_491) );
OR2x2_ASAP7_75t_L g615 ( .A(n_492), .B(n_506), .Y(n_615) );
AND2x2_ASAP7_75t_L g652 ( .A(n_492), .B(n_562), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_492), .B(n_583), .Y(n_663) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_492), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_492), .B(n_619), .Y(n_736) );
INVx5_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
AND2x2_ASAP7_75t_L g570 ( .A(n_493), .B(n_506), .Y(n_570) );
AND2x2_ASAP7_75t_L g686 ( .A(n_493), .B(n_581), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_493), .B(n_619), .Y(n_708) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_506), .Y(n_654) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_507), .Y(n_606) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g583 ( .A(n_508), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_515), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_519), .B(n_596), .Y(n_715) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_520), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g567 ( .A(n_520), .B(n_568), .Y(n_567) );
INVx5_ASAP7_75t_SL g575 ( .A(n_520), .Y(n_575) );
OR2x2_ASAP7_75t_L g598 ( .A(n_520), .B(n_568), .Y(n_598) );
OR2x2_ASAP7_75t_L g608 ( .A(n_520), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g671 ( .A(n_520), .B(n_530), .Y(n_671) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_520), .B(n_529), .Y(n_709) );
NOR4xp25_ASAP7_75t_L g730 ( .A(n_520), .B(n_651), .C(n_731), .D(n_732), .Y(n_730) );
AND2x2_ASAP7_75t_L g740 ( .A(n_520), .B(n_572), .Y(n_740) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_527), .Y(n_520) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g565 ( .A(n_529), .B(n_561), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_529), .B(n_567), .Y(n_734) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_539), .Y(n_529) );
OR2x2_ASAP7_75t_L g574 ( .A(n_530), .B(n_575), .Y(n_574) );
INVx3_ASAP7_75t_L g581 ( .A(n_530), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_530), .B(n_550), .Y(n_593) );
INVxp67_ASAP7_75t_L g596 ( .A(n_530), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_530), .B(n_568), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_530), .B(n_540), .Y(n_662) );
AND2x2_ASAP7_75t_L g677 ( .A(n_530), .B(n_572), .Y(n_677) );
OR2x2_ASAP7_75t_L g706 ( .A(n_530), .B(n_540), .Y(n_706) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_538), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_539), .B(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_539), .B(n_575), .Y(n_714) );
OR2x2_ASAP7_75t_L g735 ( .A(n_539), .B(n_612), .Y(n_735) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g549 ( .A(n_540), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g572 ( .A(n_540), .B(n_568), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_540), .B(n_550), .Y(n_587) );
AND2x2_ASAP7_75t_L g657 ( .A(n_540), .B(n_581), .Y(n_657) );
AND2x2_ASAP7_75t_L g691 ( .A(n_540), .B(n_575), .Y(n_691) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_541), .B(n_575), .Y(n_594) );
AND2x2_ASAP7_75t_L g622 ( .A(n_541), .B(n_550), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_548), .B(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_549), .A2(n_637), .B1(n_673), .B2(n_690), .C(n_692), .Y(n_689) );
INVx5_ASAP7_75t_SL g568 ( .A(n_550), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B(n_554), .Y(n_551) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
OAI33xp33_ASAP7_75t_L g588 ( .A1(n_561), .A2(n_589), .A3(n_590), .B1(n_592), .B2(n_595), .B3(n_599), .Y(n_588) );
OR2x2_ASAP7_75t_L g604 ( .A(n_561), .B(n_605), .Y(n_604) );
AOI322xp5_ASAP7_75t_L g713 ( .A1(n_561), .A2(n_630), .A3(n_637), .B1(n_714), .B2(n_715), .C1(n_716), .C2(n_719), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_561), .B(n_589), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_SL g737 ( .A1(n_561), .A2(n_589), .B(n_738), .C(n_740), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_562), .A2(n_577), .B1(n_582), .B2(n_585), .C(n_588), .Y(n_576) );
INVx1_ASAP7_75t_L g669 ( .A(n_562), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_562), .B(n_718), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B1(n_569), .B2(n_571), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g646 ( .A(n_567), .B(n_581), .Y(n_646) );
AND2x2_ASAP7_75t_L g704 ( .A(n_567), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g612 ( .A(n_568), .B(n_575), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_568), .B(n_581), .Y(n_640) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_570), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_570), .B(n_648), .Y(n_702) );
OAI321xp33_ASAP7_75t_L g721 ( .A1(n_570), .A2(n_643), .A3(n_722), .B1(n_723), .B2(n_724), .C(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g688 ( .A(n_571), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_572), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g627 ( .A(n_572), .B(n_575), .Y(n_627) );
AOI321xp33_ASAP7_75t_L g685 ( .A1(n_572), .A2(n_589), .A3(n_686), .B1(n_687), .B2(n_688), .C(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g602 ( .A(n_574), .B(n_587), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_575), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_575), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_575), .B(n_661), .Y(n_698) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g621 ( .A(n_579), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g586 ( .A(n_580), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g694 ( .A(n_581), .Y(n_694) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_584), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g617 ( .A(n_589), .Y(n_617) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_591), .B(n_626), .Y(n_675) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OR2x2_ASAP7_75t_L g639 ( .A(n_594), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g684 ( .A(n_594), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_595), .A2(n_642), .B1(n_645), .B2(n_647), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g739 ( .A(n_598), .B(n_662), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B1(n_607), .B2(n_613), .C(n_616), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g637 ( .A(n_606), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_SL g683 ( .A(n_609), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_611), .B(n_661), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_611), .A2(n_679), .B(n_681), .Y(n_678) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g724 ( .A(n_612), .B(n_706), .Y(n_724) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_SL g626 ( .A(n_615), .Y(n_626) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_620), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g670 ( .A(n_622), .B(n_671), .Y(n_670) );
INVxp67_ASAP7_75t_L g732 ( .A(n_622), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_627), .B(n_628), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_626), .B(n_644), .Y(n_680) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g701 ( .A(n_630), .Y(n_701) );
NAND5xp2_ASAP7_75t_L g631 ( .A(n_632), .B(n_649), .C(n_658), .D(n_678), .E(n_685), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_638), .C(n_641), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g673 ( .A(n_637), .Y(n_673) );
CKINVDCx16_ASAP7_75t_R g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_645), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g687 ( .A(n_647), .Y(n_687) );
OAI21xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_653), .B(n_655), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_650), .A2(n_704), .B1(n_707), .B2(n_709), .C(n_710), .Y(n_703) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
AOI321xp33_ASAP7_75t_L g658 ( .A1(n_651), .A2(n_659), .A3(n_663), .B1(n_664), .B2(n_670), .C(n_672), .Y(n_658) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g729 ( .A(n_663), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_665), .B(n_669), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g681 ( .A(n_666), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NOR2xp67_ASAP7_75t_SL g693 ( .A(n_667), .B(n_674), .Y(n_693) );
AOI321xp33_ASAP7_75t_SL g725 ( .A1(n_670), .A2(n_726), .A3(n_727), .B1(n_728), .B2(n_729), .C(n_730), .Y(n_725) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B(n_675), .C(n_676), .Y(n_672) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_683), .B(n_691), .Y(n_720) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .C(n_695), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_721), .C(n_733), .Y(n_696) );
OAI211xp5_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_699), .B(n_703), .C(n_713), .Y(n_697) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_702), .A2(n_734), .B1(n_735), .B2(n_736), .C(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g722 ( .A(n_704), .Y(n_722) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g726 ( .A(n_724), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx3_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
BUFx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NOR3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_762), .C(n_765), .Y(n_756) );
INVx1_ASAP7_75t_L g764 ( .A(n_758), .Y(n_764) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
endmodule