module fake_jpeg_20085_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_56),
.B1(n_55),
.B2(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_3),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_71),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_88),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_45),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_52),
.C(n_48),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_4),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_46),
.B(n_43),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_93),
.B(n_97),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_42),
.C(n_5),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_98),
.Y(n_106)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_96),
.A2(n_99),
.B1(n_10),
.B2(n_13),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_6),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_9),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_33),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_105),
.C(n_15),
.Y(n_110)
);

AND2x4_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_14),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_105),
.A2(n_100),
.B1(n_101),
.B2(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_110),
.C(n_102),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_106),
.C(n_107),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_108),
.B(n_18),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_17),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_23),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_24),
.Y(n_118)
);


endmodule