module fake_jpeg_2919_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

CKINVDCx10_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_88),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_87),
.B1(n_88),
.B2(n_80),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_56),
.B1(n_53),
.B2(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_101),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_79),
.B1(n_71),
.B2(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_61),
.B1(n_75),
.B2(n_53),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_78),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_58),
.C(n_62),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_71),
.B1(n_55),
.B2(n_62),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_97),
.B1(n_74),
.B2(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_57),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_1),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_55),
.B1(n_56),
.B2(n_64),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_121),
.B1(n_61),
.B2(n_67),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_117),
.B1(n_77),
.B2(n_66),
.Y(n_124)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_94),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_112),
.B(n_52),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_2),
.Y(n_130)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_95),
.B(n_69),
.C(n_76),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_139),
.B1(n_9),
.B2(n_10),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_60),
.C(n_54),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_129),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_127),
.B(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_11),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_3),
.B(n_4),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_14),
.B(n_15),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_120),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

OR2x4_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_8),
.Y(n_141)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_9),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_28),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_10),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_163),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_170),
.B1(n_165),
.B2(n_127),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_162),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_31),
.C(n_49),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_161),
.C(n_19),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_29),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_27),
.B1(n_47),
.B2(n_45),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_168),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_16),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_17),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_122),
.B(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_18),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_174),
.B1(n_182),
.B2(n_155),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_122),
.B1(n_141),
.B2(n_146),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_33),
.B(n_44),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_161),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_40),
.C(n_43),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_160),
.C(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_188),
.A2(n_190),
.B1(n_177),
.B2(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_189),
.A2(n_176),
.B1(n_173),
.B2(n_174),
.Y(n_198)
);

NOR2x1p5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_147),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_179),
.B1(n_172),
.B2(n_171),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_178),
.B(n_157),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_193),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_SL g194 ( 
.A1(n_178),
.A2(n_167),
.A3(n_164),
.B1(n_169),
.B2(n_148),
.C1(n_41),
.C2(n_51),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_SL g195 ( 
.A(n_194),
.B(n_177),
.C(n_175),
.Y(n_195)
);

AOI31xp67_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_183),
.A3(n_185),
.B(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_182),
.B(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_202),
.A2(n_187),
.B1(n_197),
.B2(n_195),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_203),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_207),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_206),
.B(n_205),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_204),
.B(n_200),
.C(n_190),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_200),
.B(n_23),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_26),
.C(n_20),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);


endmodule