module real_jpeg_15737_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_0),
.Y(n_110)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_1),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_1),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_1),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_2),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_3),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_3),
.Y(n_297)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_4),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_4),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_4),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_4),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_4),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_5),
.A2(n_66),
.B1(n_71),
.B2(n_74),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_5),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_5),
.A2(n_74),
.B1(n_129),
.B2(n_132),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g238 ( 
.A1(n_5),
.A2(n_239),
.A3(n_242),
.B1(n_243),
.B2(n_248),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_5),
.B(n_31),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_5),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_5),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_5),
.B(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_6),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_6),
.A2(n_21),
.B1(n_275),
.B2(n_279),
.Y(n_274)
);

OAI22x1_ASAP7_75t_L g41 ( 
.A1(n_7),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_7),
.A2(n_45),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_7),
.A2(n_45),
.B1(n_204),
.B2(n_207),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_7),
.A2(n_45),
.B1(n_265),
.B2(n_268),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_8),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_11),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_232),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_231),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp67_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_167),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_16),
.B(n_167),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_97),
.C(n_123),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_17),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_58),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_18),
.B(n_59),
.C(n_89),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_40),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_20),
.B(n_49),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_21),
.A2(n_76),
.B(n_78),
.C(n_83),
.Y(n_75)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_26),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_30),
.Y(n_117)
);

NOR2x1p5_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_31),
.B(n_41),
.Y(n_229)
);

AO22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_36),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_50)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_49),
.Y(n_327)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_54),
.Y(n_326)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_88),
.B2(n_89),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_75),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_61),
.B(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_70),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_62),
.B(n_78),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_62),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_68),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_73),
.Y(n_143)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_73),
.Y(n_247)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_73),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_74),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_74),
.B(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_74),
.A2(n_196),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_74),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_75),
.B(n_263),
.Y(n_301)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_82),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_83),
.A2(n_174),
.B(n_180),
.Y(n_173)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_86),
.Y(n_262)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_90),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_90),
.B(n_212),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_90)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_97),
.A2(n_123),
.B1(n_124),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_97),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_118),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_98),
.A2(n_118),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_98),
.Y(n_330)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.A3(n_105),
.B1(n_111),
.B2(n_115),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_100),
.A2(n_183),
.B1(n_187),
.B2(n_196),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_103),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_115),
.B(n_324),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_118),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B(n_122),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g259 ( 
.A1(n_122),
.A2(n_260),
.B(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_148),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_128),
.A2(n_137),
.B(n_149),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_128),
.B(n_149),
.Y(n_257)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_136),
.Y(n_303)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_137),
.B(n_163),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_137),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_143),
.B1(n_144),
.B2(n_147),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_148),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_163),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_149),
.B(n_274),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B1(n_156),
.B2(n_160),
.Y(n_150)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_161),
.Y(n_241)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_199),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_180),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_224),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_210),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_221),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_218),
.B2(n_220),
.Y(n_212)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_229),
.B(n_320),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_334),
.B(n_339),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_311),
.B(n_333),
.Y(n_234)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_286),
.B(n_310),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_258),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_L g310 ( 
.A(n_237),
.B(n_258),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_255),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_238),
.B(n_255),
.Y(n_308)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_271),
.Y(n_258)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_264),
.Y(n_299)
);

INVx4_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_284),
.C(n_332),
.Y(n_331)
);

OAI21x1_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_305),
.B(n_309),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_300),
.B(n_304),
.Y(n_287)
);

NOR2x1_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_298),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_294),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_308),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_331),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_331),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_328),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_319),
.C(n_328),
.Y(n_338)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_338),
.Y(n_339)
);


endmodule