module fake_jpeg_13409_n_495 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_495);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_495;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_61),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_63),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_66),
.B(n_68),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_67),
.B(n_75),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_33),
.B(n_15),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_70),
.B(n_83),
.Y(n_187)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_72),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_79),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

CKINVDCx6p67_ASAP7_75t_R g183 ( 
.A(n_82),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_15),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_85),
.B(n_86),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_27),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_45),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_87),
.B(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_89),
.B(n_92),
.Y(n_173)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx2_ASAP7_75t_R g92 ( 
.A(n_22),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_96),
.B(n_98),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_97),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_99),
.Y(n_189)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_100),
.Y(n_184)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_103),
.B(n_107),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_13),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_104),
.B(n_119),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_46),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_114),
.Y(n_191)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_113),
.B(n_115),
.Y(n_175)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_118),
.Y(n_193)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_117),
.B(n_120),
.Y(n_157)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_19),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_42),
.Y(n_119)
);

BUFx16f_ASAP7_75t_L g120 ( 
.A(n_19),
.Y(n_120)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_25),
.B(n_35),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_46),
.B1(n_57),
.B2(n_36),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_122),
.A2(n_128),
.B1(n_144),
.B2(n_154),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_81),
.A2(n_32),
.B1(n_57),
.B2(n_44),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_124),
.A2(n_129),
.B1(n_139),
.B2(n_141),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_59),
.B1(n_55),
.B2(n_54),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_32),
.B1(n_25),
.B2(n_35),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_133),
.A2(n_146),
.B(n_183),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_135),
.A2(n_146),
.B1(n_184),
.B2(n_175),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_72),
.A2(n_25),
.B1(n_35),
.B2(n_54),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_90),
.A2(n_59),
.B1(n_55),
.B2(n_52),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_52),
.B1(n_50),
.B2(n_42),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_143),
.A2(n_161),
.B1(n_181),
.B2(n_131),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_61),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_153),
.A2(n_181),
.B1(n_161),
.B2(n_143),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_65),
.A2(n_11),
.B1(n_3),
.B2(n_5),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_155),
.A2(n_163),
.B1(n_172),
.B2(n_174),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_73),
.A2(n_80),
.B1(n_77),
.B2(n_112),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_93),
.A2(n_117),
.B1(n_121),
.B2(n_69),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_92),
.B(n_1),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_164),
.B(n_182),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_106),
.A2(n_74),
.B1(n_109),
.B2(n_101),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_165),
.A2(n_166),
.B1(n_177),
.B2(n_192),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_113),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_9),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_182),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_116),
.A2(n_9),
.B1(n_118),
.B2(n_87),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_100),
.A2(n_84),
.B1(n_82),
.B2(n_120),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_84),
.A2(n_22),
.B1(n_32),
.B2(n_57),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_97),
.A2(n_88),
.B1(n_99),
.B2(n_102),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_97),
.B(n_82),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_60),
.A2(n_61),
.B1(n_77),
.B2(n_80),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_186),
.A2(n_134),
.B1(n_138),
.B2(n_158),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_92),
.B(n_22),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_157),
.B(n_175),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_81),
.A2(n_22),
.B1(n_32),
.B2(n_57),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_195),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_196),
.B(n_200),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_201),
.A2(n_252),
.B1(n_233),
.B2(n_206),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_202),
.B(n_217),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_203),
.A2(n_148),
.B1(n_137),
.B2(n_162),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_145),
.B(n_187),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_205),
.B(n_210),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_146),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_206),
.Y(n_273)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_207),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_191),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_208),
.B(n_212),
.Y(n_260)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_153),
.B(n_136),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_213),
.A2(n_226),
.B(n_204),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_150),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_223),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_215),
.A2(n_221),
.B(n_226),
.C(n_218),
.Y(n_269)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_185),
.B(n_126),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_153),
.B(n_140),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_239),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_220),
.B(n_227),
.Y(n_303)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_156),
.Y(n_222)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_136),
.C(n_140),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_224),
.B(n_230),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_178),
.B(n_176),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_151),
.B(n_176),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_228),
.B(n_233),
.Y(n_278)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_127),
.Y(n_231)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_231),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_142),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_135),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_236),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_183),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_237),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_153),
.B(n_151),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_125),
.Y(n_240)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_130),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_241),
.B(n_242),
.Y(n_306)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_160),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_243),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_127),
.A2(n_194),
.B1(n_123),
.B2(n_147),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_245),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_132),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_160),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_247),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_130),
.B(n_131),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_255),
.Y(n_274)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_249),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_183),
.B(n_179),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_256),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_134),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_253),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_138),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_123),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_179),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_147),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_157),
.B(n_194),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_148),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_209),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_261),
.A2(n_268),
.B1(n_269),
.B2(n_246),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_162),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_267),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_212),
.A2(n_137),
.B1(n_219),
.B2(n_239),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_272),
.A2(n_282),
.B1(n_288),
.B2(n_249),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_231),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_201),
.A2(n_215),
.B1(n_204),
.B2(n_248),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_222),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_215),
.A2(n_224),
.B1(n_208),
.B2(n_197),
.Y(n_288)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_241),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_202),
.B(n_207),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_305),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_211),
.B(n_225),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_330),
.Y(n_353)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_264),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_311),
.B(n_314),
.Y(n_375)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_312),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_273),
.A2(n_215),
.B1(n_251),
.B2(n_231),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_313),
.A2(n_320),
.B(n_327),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_291),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_318),
.B(n_339),
.Y(n_371)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_290),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_323),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_273),
.A2(n_240),
.B(n_238),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_322),
.A2(n_296),
.B(n_286),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_277),
.B(n_216),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_282),
.A2(n_237),
.B1(n_198),
.B2(n_244),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_325),
.A2(n_326),
.B1(n_261),
.B2(n_267),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_280),
.A2(n_195),
.B(n_199),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_328),
.Y(n_372)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_331),
.Y(n_351)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_334),
.Y(n_355)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_336),
.Y(n_362)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_306),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_274),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_338),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_265),
.B(n_232),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_306),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_340),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_268),
.A2(n_234),
.B1(n_259),
.B2(n_242),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_341),
.A2(n_272),
.B1(n_270),
.B2(n_284),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_267),
.B(n_229),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_345),
.Y(n_374)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_343),
.A2(n_346),
.B(n_267),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_266),
.Y(n_344)
);

AOI221xp5_ASAP7_75t_L g364 ( 
.A1(n_344),
.A2(n_295),
.B1(n_271),
.B2(n_278),
.C(n_303),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_265),
.B(n_260),
.Y(n_345)
);

BUFx12_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_354),
.A2(n_357),
.B(n_368),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_356),
.A2(n_361),
.B1(n_369),
.B2(n_331),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_322),
.A2(n_305),
.B(n_296),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_359),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_337),
.A2(n_280),
.B(n_276),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_285),
.C(n_288),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_373),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_325),
.A2(n_269),
.B1(n_260),
.B2(n_293),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_364),
.B(n_320),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_365),
.A2(n_317),
.B1(n_338),
.B2(n_332),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_337),
.A2(n_283),
.B(n_297),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_317),
.A2(n_269),
.B1(n_299),
.B2(n_300),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_302),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_375),
.B(n_343),
.Y(n_377)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_386),
.C(n_387),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_378),
.B(n_393),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_339),
.Y(n_380)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_355),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_388),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_382),
.A2(n_384),
.B1(n_398),
.B2(n_399),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_309),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_383),
.B(n_390),
.C(n_368),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_361),
.A2(n_313),
.B1(n_345),
.B2(n_269),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_363),
.B(n_308),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_319),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_367),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_392),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_320),
.Y(n_390)
);

AOI221xp5_ASAP7_75t_L g391 ( 
.A1(n_359),
.A2(n_327),
.B1(n_342),
.B2(n_328),
.C(n_329),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_SL g415 ( 
.A(n_391),
.B(n_351),
.C(n_354),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_355),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_330),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_394),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_376),
.B(n_304),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_397),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_373),
.B(n_324),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_369),
.A2(n_341),
.B1(n_342),
.B2(n_335),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_356),
.A2(n_316),
.B1(n_270),
.B2(n_263),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_357),
.A2(n_301),
.B(n_312),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_400),
.A2(n_347),
.B(n_358),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_402),
.A2(n_365),
.B1(n_370),
.B2(n_362),
.Y(n_412)
);

O2A1O1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_404),
.A2(n_396),
.B(n_379),
.C(n_400),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_371),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_406),
.C(n_414),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_388),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_416),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_412),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_350),
.Y(n_413)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_374),
.C(n_347),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_415),
.B(n_389),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_396),
.A2(n_351),
.B(n_370),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_349),
.Y(n_417)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_417),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_384),
.A2(n_351),
.B1(n_362),
.B2(n_372),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_349),
.Y(n_423)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_423),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_390),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_374),
.C(n_394),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_427),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_414),
.B(n_406),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_416),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_430),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_408),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_432),
.B(n_433),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_378),
.Y(n_433)
);

AO21x1_ASAP7_75t_L g434 ( 
.A1(n_420),
.A2(n_396),
.B(n_379),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_434),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_422),
.A2(n_398),
.B1(n_399),
.B2(n_380),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_410),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_442),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_405),
.B(n_402),
.C(n_393),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_424),
.C(n_404),
.Y(n_454)
);

BUFx12_ASAP7_75t_L g439 ( 
.A(n_422),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_439),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_446),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_440),
.B(n_409),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_441),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_451),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_418),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_450),
.B(n_436),
.Y(n_460)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_431),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_403),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_452),
.A2(n_408),
.B(n_407),
.Y(n_463)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_430),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_453),
.B(n_454),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_454),
.B(n_442),
.Y(n_457)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_457),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_456),
.B(n_428),
.C(n_427),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_462),
.Y(n_470)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_460),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_455),
.A2(n_410),
.B1(n_426),
.B2(n_435),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_446),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_444),
.A2(n_415),
.B(n_426),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_464),
.A2(n_466),
.B(n_434),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_428),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_465),
.B(n_449),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_449),
.A2(n_425),
.B(n_452),
.Y(n_466)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_468),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_407),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_471),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_467),
.B(n_444),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_465),
.C(n_457),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_476),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_459),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_479),
.Y(n_487)
);

BUFx24_ASAP7_75t_SL g479 ( 
.A(n_474),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_472),
.A2(n_458),
.B(n_448),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_480),
.B(n_481),
.C(n_475),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_466),
.C(n_443),
.Y(n_481)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_484),
.Y(n_489)
);

AOI322xp5_ASAP7_75t_L g485 ( 
.A1(n_482),
.A2(n_468),
.A3(n_403),
.B1(n_439),
.B2(n_419),
.C1(n_469),
.C2(n_401),
.Y(n_485)
);

AOI322xp5_ASAP7_75t_L g491 ( 
.A1(n_485),
.A2(n_401),
.A3(n_438),
.B1(n_366),
.B2(n_421),
.C1(n_346),
.C2(n_348),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_445),
.C(n_430),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_486),
.A2(n_488),
.B(n_438),
.Y(n_490)
);

AOI31xp67_ASAP7_75t_SL g488 ( 
.A1(n_483),
.A2(n_419),
.A3(n_439),
.B(n_445),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_487),
.C(n_421),
.Y(n_493)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_491),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_489),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_492),
.Y(n_495)
);


endmodule