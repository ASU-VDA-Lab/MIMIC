module real_jpeg_2726_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_1),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_2),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_4),
.A2(n_30),
.B1(n_34),
.B2(n_63),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_63),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_5),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_80),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_30),
.B1(n_34),
.B2(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_6),
.A2(n_57),
.B1(n_58),
.B2(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_66),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_30),
.B1(n_34),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_70),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_70),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_70),
.Y(n_215)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_43),
.B1(n_57),
.B2(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_15),
.B(n_116),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_15),
.A2(n_24),
.B(n_54),
.C(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_15),
.B(n_56),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_104),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_15),
.B(n_41),
.C(n_83),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_104),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_15),
.B(n_46),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_15),
.B(n_87),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_20),
.B(n_107),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_92),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_21),
.B(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_22),
.B(n_51),
.C(n_67),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_23),
.A2(n_37),
.B1(n_38),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_23),
.Y(n_146)
);

AOI32xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.A3(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_24),
.B(n_54),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_36),
.Y(n_71)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_76)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_30),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_153),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_40),
.A2(n_41),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_41),
.B(n_211),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_44),
.A2(n_45),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_44),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_44),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_44),
.A2(n_45),
.B1(n_185),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_45),
.A2(n_153),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_45),
.B(n_172),
.Y(n_187)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_48),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_46),
.A2(n_171),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_67),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_61),
.B(n_64),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_52),
.A2(n_64),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_56),
.B1(n_62),
.B2(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_65),
.Y(n_121)
);

AO22x2_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_56)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_58),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_57),
.A2(n_60),
.B(n_104),
.Y(n_168)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_58),
.B(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B(n_72),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_75),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_77),
.A2(n_92),
.B1(n_93),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_88),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_86),
.B1(n_87),
.B2(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_81),
.A2(n_162),
.B(n_164),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_85),
.A2(n_97),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_85),
.A2(n_163),
.B1(n_181),
.B2(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_87),
.B(n_98),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_89),
.A2(n_104),
.B(n_187),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.C(n_101),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_101),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_124),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_122),
.B2(n_123),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B(n_121),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_121),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_154),
.B(n_232),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_138),
.B(n_141),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_147),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_147),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_152),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_175),
.B(n_231),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_173),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_157),
.B(n_173),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_166),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_161),
.B(n_166),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_193),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_169),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_226),
.B(n_230),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_195),
.B(n_225),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_188),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_183),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_184),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_192),
.C(n_194),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_207),
.B(n_224),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_218),
.B(n_223),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_213),
.B(n_217),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_216),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_221),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_229),
.Y(n_230)
);


endmodule