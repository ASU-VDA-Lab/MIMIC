module fake_netlist_6_373_n_1587 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1587);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1587;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_105),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_19),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_73),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_41),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_36),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_48),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_131),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_15),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_148),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_32),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_58),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_47),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_96),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_16),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_14),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_1),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_35),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_59),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_64),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_53),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_101),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_42),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_145),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_22),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_129),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_20),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_126),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_54),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_123),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_5),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_47),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_90),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_53),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_44),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_14),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_86),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_81),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_130),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_35),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_60),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_15),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_133),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_107),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_134),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_99),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_82),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_140),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_141),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_144),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_10),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_100),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_118),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_112),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_116),
.Y(n_228)
);

BUFx2_ASAP7_75t_SL g229 ( 
.A(n_154),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_72),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_76),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_48),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_13),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_92),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_34),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_25),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_8),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_150),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_74),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_50),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_113),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_0),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_49),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_52),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_70),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_80),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_17),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_68),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_57),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_16),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_89),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_33),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_142),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_152),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_138),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_117),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_43),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_61),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_77),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_137),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_102),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_29),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_65),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_46),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_52),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_143),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_50),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_127),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_7),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_159),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_18),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_88),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_12),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_54),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_43),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_7),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_84),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_66),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_45),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_11),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_155),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_4),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_20),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_58),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_111),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_45),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_24),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_38),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_56),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_25),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_30),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_139),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_4),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_115),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_91),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_12),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_151),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_1),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_103),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_42),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_37),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_97),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_87),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_136),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_36),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_38),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_56),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_69),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_158),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_275),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_207),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_245),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_207),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_290),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_249),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_207),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_207),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_287),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_292),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_165),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_207),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_164),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_244),
.B(n_2),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_207),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_210),
.B(n_3),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_207),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_287),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_256),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_207),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_173),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_192),
.Y(n_340)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_215),
.B(n_3),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_176),
.B(n_6),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_269),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_186),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_186),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_194),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_276),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_278),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_199),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_251),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_251),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_168),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_310),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_311),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_309),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_210),
.B(n_6),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_168),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_168),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_200),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_237),
.B(n_8),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_172),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_312),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_168),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_168),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_262),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_305),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_164),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_215),
.B(n_9),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_262),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_193),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_195),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_262),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_197),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_173),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_203),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_262),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_205),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_224),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_201),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_181),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_190),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_196),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_202),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_230),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_234),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_212),
.B(n_9),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_273),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_235),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_273),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_237),
.B(n_11),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_279),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_238),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_239),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_243),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_246),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_321),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_339),
.B(n_198),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_358),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_359),
.Y(n_405)
);

INVxp33_ASAP7_75t_SL g406 ( 
.A(n_318),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_336),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_160),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_367),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_198),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_160),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_225),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_324),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_320),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_371),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_225),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_331),
.Y(n_419)
);

NOR2x1_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_241),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_368),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_320),
.A2(n_325),
.B(n_322),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_337),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_372),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_375),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_378),
.B(n_161),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_333),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_322),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_325),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_329),
.B(n_206),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_381),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_338),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_391),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_391),
.B(n_163),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_323),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_341),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_369),
.B(n_204),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_393),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g447 ( 
.A(n_340),
.B(n_208),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_347),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_323),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_342),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_344),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_342),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_362),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_345),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_351),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_352),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_334),
.B(n_161),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_340),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g463 ( 
.A1(n_357),
.A2(n_279),
.B(n_248),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_346),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_328),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_361),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_332),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_356),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_407),
.B(n_453),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_433),
.Y(n_471)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_413),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_468),
.B(n_346),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_419),
.A2(n_328),
.B1(n_396),
.B2(n_395),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_349),
.Y(n_478)
);

BUFx4f_ASAP7_75t_L g479 ( 
.A(n_463),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_349),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_413),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_360),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_416),
.Y(n_483)
);

NOR2x1p5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_360),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_415),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_432),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_415),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_377),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_R g489 ( 
.A(n_410),
.B(n_348),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_R g491 ( 
.A(n_406),
.B(n_379),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_419),
.A2(n_397),
.B1(n_396),
.B2(n_395),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_407),
.B(n_379),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_423),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_453),
.B(n_380),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_432),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_380),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_456),
.B(n_319),
.Y(n_500)
);

INVx4_ASAP7_75t_SL g501 ( 
.A(n_443),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_467),
.B(n_411),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_453),
.B(n_386),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_467),
.B(n_386),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_425),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_455),
.A2(n_397),
.B1(n_394),
.B2(n_390),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_460),
.B(n_387),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_411),
.B(n_387),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_409),
.B(n_390),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_421),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_455),
.A2(n_282),
.B1(n_299),
.B2(n_294),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_455),
.B(n_394),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_443),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_411),
.B(n_241),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_413),
.B(n_170),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_455),
.B(n_191),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_413),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_418),
.B(n_177),
.Y(n_525)
);

AND2x2_ASAP7_75t_SL g526 ( 
.A(n_455),
.B(n_463),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_409),
.B(n_327),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_455),
.B(n_204),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_447),
.B(n_374),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_447),
.B(n_206),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_418),
.B(n_462),
.Y(n_531)
);

BUFx4f_ASAP7_75t_L g532 ( 
.A(n_463),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_462),
.A2(n_298),
.B1(n_271),
.B2(n_283),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_404),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_442),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_442),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g537 ( 
.A(n_417),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_421),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_457),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_446),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_401),
.B(n_252),
.C(n_247),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_422),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_415),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_415),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_420),
.B(n_204),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_449),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_464),
.A2(n_270),
.B1(n_268),
.B2(n_257),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_463),
.A2(n_277),
.B1(n_286),
.B2(n_233),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_401),
.B(n_293),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_435),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_401),
.B(n_264),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_461),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_435),
.Y(n_553)
);

NAND2x1p5_ASAP7_75t_L g554 ( 
.A(n_423),
.B(n_184),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_463),
.A2(n_288),
.B1(n_304),
.B2(n_229),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_449),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_443),
.B(n_204),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_452),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_452),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_465),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_458),
.B(n_272),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_428),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_438),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_438),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_438),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_422),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_434),
.B(n_209),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_417),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_399),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_464),
.B(n_211),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_451),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_399),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_399),
.Y(n_573)
);

NAND2x1p5_ASAP7_75t_L g574 ( 
.A(n_423),
.B(n_217),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_451),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_399),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_412),
.B(n_272),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_435),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_458),
.B(n_272),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_438),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_443),
.A2(n_214),
.B1(n_227),
.B2(n_231),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_403),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_427),
.B(n_441),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_427),
.B(n_350),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_443),
.B(n_214),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_435),
.Y(n_586)
);

CKINVDCx6p67_ASAP7_75t_R g587 ( 
.A(n_400),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_441),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_466),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_403),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_445),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_466),
.A2(n_363),
.B1(n_355),
.B2(n_354),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_426),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_443),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_443),
.A2(n_214),
.B1(n_267),
.B2(n_220),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_445),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_418),
.B(n_162),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_454),
.B(n_162),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_526),
.A2(n_443),
.B1(n_187),
.B2(n_240),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_512),
.B(n_499),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_526),
.A2(n_281),
.B1(n_314),
.B2(n_301),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_531),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_522),
.B(n_509),
.Y(n_604)
);

AND2x6_ASAP7_75t_SL g605 ( 
.A(n_476),
.B(n_242),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_500),
.B(n_436),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_481),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_503),
.B(n_454),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_479),
.A2(n_532),
.B(n_494),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_478),
.A2(n_218),
.B1(n_213),
.B2(n_317),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_569),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_527),
.B(n_454),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_471),
.B(n_405),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_472),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_469),
.B(n_459),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_L g616 ( 
.A(n_555),
.B(n_216),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_471),
.B(n_405),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_500),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_478),
.A2(n_260),
.B1(n_219),
.B2(n_221),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_481),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_569),
.Y(n_621)
);

BUFx8_ASAP7_75t_L g622 ( 
.A(n_568),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_473),
.B(n_408),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_572),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_572),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_573),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_518),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_542),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_472),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_523),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_479),
.A2(n_214),
.B1(n_263),
.B2(n_266),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_480),
.A2(n_259),
.B1(n_222),
.B2(n_223),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_498),
.B(n_445),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_511),
.B(n_445),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_539),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_482),
.B(n_445),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_482),
.B(n_166),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_532),
.A2(n_548),
.B1(n_510),
.B2(n_488),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_495),
.B(n_445),
.Y(n_639)
);

A2O1A1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_551),
.A2(n_440),
.B(n_300),
.C(n_303),
.Y(n_640)
);

AOI221xp5_ASAP7_75t_L g641 ( 
.A1(n_533),
.A2(n_178),
.B1(n_167),
.B2(n_169),
.C(n_175),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_504),
.B(n_166),
.Y(n_642)
);

INVx8_ASAP7_75t_L g643 ( 
.A(n_570),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_504),
.B(n_171),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_505),
.B(n_171),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_540),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_549),
.A2(n_295),
.B1(n_169),
.B2(n_175),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_513),
.B(n_459),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_514),
.B(n_450),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_538),
.B(n_450),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_516),
.A2(n_484),
.B1(n_570),
.B2(n_536),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_546),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_469),
.B(n_414),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_576),
.Y(n_654)
);

NAND3xp33_ASAP7_75t_L g655 ( 
.A(n_541),
.B(n_255),
.C(n_254),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_474),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_598),
.B(n_450),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_486),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_520),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_520),
.B(n_430),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_556),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_535),
.B(n_536),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_525),
.B(n_430),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_525),
.B(n_431),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_558),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_559),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_309),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_542),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_584),
.A2(n_583),
.B1(n_508),
.B2(n_470),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_566),
.B(n_439),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_580),
.B(n_431),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_529),
.B(n_174),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_492),
.B(n_174),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_563),
.B(n_444),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_566),
.B(n_424),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_477),
.B(n_179),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_582),
.Y(n_678)
);

BUFx8_ASAP7_75t_L g679 ( 
.A(n_568),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_570),
.B(n_179),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_564),
.B(n_565),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_590),
.B(n_226),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_570),
.B(n_185),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_519),
.B(n_228),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_474),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_515),
.A2(n_214),
.B1(n_178),
.B2(n_183),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_588),
.B(n_429),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_486),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_554),
.A2(n_236),
.B(n_261),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_561),
.B(n_232),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_561),
.B(n_250),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_490),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_475),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_579),
.B(n_253),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_588),
.B(n_448),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_577),
.B(n_188),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_530),
.B(n_189),
.Y(n_697)
);

INVx8_ASAP7_75t_L g698 ( 
.A(n_567),
.Y(n_698)
);

NOR3xp33_ASAP7_75t_L g699 ( 
.A(n_597),
.B(n_316),
.C(n_189),
.Y(n_699)
);

BUFx8_ASAP7_75t_L g700 ( 
.A(n_589),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_575),
.B(n_291),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_547),
.B(n_316),
.C(n_274),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_521),
.B(n_258),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_521),
.B(n_265),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_567),
.A2(n_274),
.B1(n_284),
.B2(n_285),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_524),
.B(n_543),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_554),
.A2(n_315),
.B1(n_313),
.B2(n_308),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_524),
.B(n_285),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g709 ( 
.A1(n_554),
.A2(n_289),
.B(n_307),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_497),
.Y(n_710)
);

AND2x6_ASAP7_75t_SL g711 ( 
.A(n_567),
.B(n_315),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_567),
.B(n_13),
.Y(n_712)
);

INVx8_ASAP7_75t_L g713 ( 
.A(n_483),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_524),
.B(n_289),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_545),
.A2(n_307),
.B1(n_308),
.B2(n_313),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_537),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_490),
.Y(n_717)
);

NOR3xp33_ASAP7_75t_L g718 ( 
.A(n_493),
.B(n_306),
.C(n_297),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_L g719 ( 
.A(n_537),
.B(n_306),
.C(n_297),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_545),
.A2(n_296),
.B1(n_295),
.B2(n_291),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_496),
.A2(n_296),
.B(n_280),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_506),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_496),
.A2(n_280),
.B(n_183),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_543),
.B(n_182),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_543),
.B(n_180),
.Y(n_725)
);

NOR2x1p5_ASAP7_75t_L g726 ( 
.A(n_587),
.B(n_19),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_553),
.B(n_62),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_574),
.B(n_21),
.Y(n_728)
);

INVxp33_ASAP7_75t_L g729 ( 
.A(n_489),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_491),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_553),
.B(n_153),
.Y(n_731)
);

O2A1O1Ixp5_ASAP7_75t_L g732 ( 
.A1(n_594),
.A2(n_21),
.B(n_23),
.C(n_26),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_553),
.B(n_132),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_636),
.A2(n_639),
.B(n_609),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_601),
.A2(n_604),
.B1(n_638),
.B2(n_670),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_671),
.B(n_571),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_612),
.B(n_574),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_614),
.A2(n_594),
.B(n_517),
.Y(n_738)
);

NOR2x1p5_ASAP7_75t_L g739 ( 
.A(n_660),
.B(n_483),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_730),
.B(n_507),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_599),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_620),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_614),
.A2(n_550),
.B(n_502),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_620),
.Y(n_744)
);

OA22x2_ASAP7_75t_L g745 ( 
.A1(n_712),
.A2(n_592),
.B1(n_507),
.B2(n_571),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_631),
.A2(n_595),
.B1(n_581),
.B2(n_562),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_651),
.B(n_560),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_608),
.B(n_657),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_668),
.B(n_571),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_730),
.B(n_560),
.Y(n_750)
);

INVx11_ASAP7_75t_L g751 ( 
.A(n_622),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_713),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_685),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_709),
.A2(n_557),
.B(n_585),
.C(n_534),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_628),
.B(n_560),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_656),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_678),
.B(n_528),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_659),
.B(n_552),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_693),
.Y(n_759)
);

AO21x1_ASAP7_75t_L g760 ( 
.A1(n_689),
.A2(n_596),
.B(n_586),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_690),
.B(n_544),
.Y(n_761)
);

OAI21xp33_ASAP7_75t_L g762 ( 
.A1(n_602),
.A2(n_552),
.B(n_593),
.Y(n_762)
);

AOI21x1_ASAP7_75t_L g763 ( 
.A1(n_706),
.A2(n_485),
.B(n_578),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_703),
.A2(n_487),
.B(n_544),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_620),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_603),
.B(n_501),
.Y(n_766)
);

AO21x1_ASAP7_75t_L g767 ( 
.A1(n_637),
.A2(n_23),
.B(n_26),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_647),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_691),
.B(n_487),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_704),
.A2(n_487),
.B(n_591),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_694),
.B(n_635),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_627),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_661),
.A2(n_591),
.B(n_75),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_628),
.B(n_552),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_732),
.A2(n_591),
.B(n_67),
.Y(n_775)
);

AO22x1_ASAP7_75t_L g776 ( 
.A1(n_718),
.A2(n_593),
.B1(n_28),
.B2(n_30),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_664),
.A2(n_78),
.B(n_125),
.Y(n_777)
);

AO21x1_ASAP7_75t_L g778 ( 
.A1(n_642),
.A2(n_27),
.B(n_31),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_665),
.A2(n_63),
.B(n_122),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_646),
.B(n_121),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_681),
.A2(n_98),
.B(n_119),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_669),
.B(n_593),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_676),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_696),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_652),
.B(n_37),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_647),
.A2(n_644),
.B(n_640),
.C(n_645),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_600),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_649),
.A2(n_106),
.B(n_104),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_627),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_627),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_650),
.A2(n_95),
.B(n_94),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_684),
.A2(n_93),
.B(n_85),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_708),
.A2(n_83),
.B(n_40),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_600),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_662),
.B(n_49),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_659),
.Y(n_796)
);

BUFx4f_ASAP7_75t_L g797 ( 
.A(n_713),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_714),
.A2(n_648),
.B(n_633),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_616),
.A2(n_51),
.B(n_55),
.C(n_57),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_673),
.A2(n_51),
.B(n_683),
.C(n_680),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_666),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_713),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_669),
.B(n_729),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_602),
.A2(n_707),
.B1(n_712),
.B2(n_641),
.Y(n_804)
);

BUFx8_ASAP7_75t_L g805 ( 
.A(n_606),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_643),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_634),
.A2(n_675),
.B(n_672),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_667),
.B(n_607),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_682),
.A2(n_724),
.B(n_725),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_663),
.B(n_673),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_674),
.B(n_677),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_630),
.B(n_613),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_680),
.B(n_683),
.Y(n_813)
);

BUFx4f_ASAP7_75t_L g814 ( 
.A(n_687),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_617),
.B(n_623),
.Y(n_815)
);

NAND2x1_ASAP7_75t_L g816 ( 
.A(n_710),
.B(n_722),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_611),
.A2(n_654),
.B(n_626),
.Y(n_817)
);

CKINVDCx8_ASAP7_75t_R g818 ( 
.A(n_605),
.Y(n_818)
);

OAI21xp33_ASAP7_75t_L g819 ( 
.A1(n_707),
.A2(n_641),
.B(n_686),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_621),
.A2(n_625),
.B(n_624),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_727),
.A2(n_733),
.B(n_731),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_658),
.A2(n_717),
.B(n_692),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_615),
.B(n_716),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_643),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_699),
.B(n_610),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_688),
.B(n_619),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_712),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_701),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_687),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_632),
.B(n_723),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_705),
.A2(n_698),
.B1(n_715),
.B2(n_720),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_697),
.A2(n_655),
.B(n_721),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_698),
.A2(n_702),
.B1(n_686),
.B2(n_718),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_653),
.B(n_687),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_721),
.A2(n_723),
.B(n_719),
.C(n_653),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_719),
.B(n_698),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_653),
.A2(n_695),
.B(n_726),
.C(n_711),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_695),
.B(n_622),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_679),
.A2(n_604),
.B(n_601),
.C(n_499),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_695),
.A2(n_631),
.B1(n_600),
.B2(n_602),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_700),
.B(n_679),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_700),
.B(n_631),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_604),
.A2(n_601),
.B(n_499),
.C(n_509),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_636),
.A2(n_532),
.B(n_479),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_604),
.B(n_612),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_636),
.A2(n_532),
.B(n_479),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_609),
.A2(n_532),
.B(n_479),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_599),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_599),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_599),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_618),
.B(n_456),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_622),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_620),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_599),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_631),
.A2(n_600),
.B1(n_602),
.B2(n_670),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_601),
.A2(n_728),
.B1(n_638),
.B2(n_604),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_599),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_599),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_670),
.B(n_500),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_631),
.A2(n_600),
.B1(n_602),
.B2(n_670),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_601),
.B(n_456),
.C(n_584),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_601),
.A2(n_604),
.B1(n_638),
.B2(n_670),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_609),
.A2(n_532),
.B(n_479),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_601),
.A2(n_638),
.B(n_604),
.C(n_709),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_601),
.B(n_456),
.C(n_584),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_604),
.B(n_612),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_604),
.B(n_612),
.Y(n_867)
);

NAND2x1p5_ASAP7_75t_L g868 ( 
.A(n_614),
.B(n_629),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_601),
.A2(n_604),
.B1(n_638),
.B2(n_670),
.Y(n_869)
);

NOR2x1_ASAP7_75t_R g870 ( 
.A(n_660),
.B(n_483),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_601),
.B(n_456),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_L g872 ( 
.A(n_601),
.B(n_456),
.C(n_584),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_801),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_845),
.B(n_866),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_855),
.A2(n_860),
.B(n_819),
.C(n_867),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_742),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_847),
.A2(n_863),
.B(n_844),
.Y(n_877)
);

AO31x2_ASAP7_75t_L g878 ( 
.A1(n_760),
.A2(n_855),
.A3(n_860),
.B(n_737),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_847),
.A2(n_863),
.B(n_846),
.Y(n_879)
);

AND3x1_ASAP7_75t_L g880 ( 
.A(n_861),
.B(n_865),
.C(n_872),
.Y(n_880)
);

OAI21x1_ASAP7_75t_SL g881 ( 
.A1(n_767),
.A2(n_778),
.B(n_787),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_742),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_763),
.A2(n_770),
.B(n_764),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_766),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_851),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_734),
.A2(n_769),
.B(n_761),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_815),
.A2(n_821),
.B(n_807),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_735),
.B(n_862),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_813),
.A2(n_864),
.B(n_840),
.C(n_804),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_869),
.A2(n_843),
.B(n_856),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_736),
.B(n_749),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_748),
.B(n_859),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_804),
.B(n_871),
.Y(n_893)
);

AND3x2_ASAP7_75t_L g894 ( 
.A(n_755),
.B(n_774),
.C(n_782),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_840),
.B(n_810),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_811),
.A2(n_825),
.B1(n_833),
.B2(n_842),
.Y(n_896)
);

AO21x1_ASAP7_75t_L g897 ( 
.A1(n_787),
.A2(n_794),
.B(n_775),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_754),
.A2(n_798),
.B(n_809),
.Y(n_898)
);

NAND3xp33_ASAP7_75t_SL g899 ( 
.A(n_762),
.B(n_800),
.C(n_783),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_756),
.Y(n_900)
);

OAI222xp33_ASAP7_75t_L g901 ( 
.A1(n_794),
.A2(n_745),
.B1(n_768),
.B2(n_799),
.C1(n_831),
.C2(n_783),
.Y(n_901)
);

OAI22x1_ASAP7_75t_L g902 ( 
.A1(n_827),
.A2(n_740),
.B1(n_829),
.B2(n_750),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_771),
.B(n_812),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_823),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_830),
.B(n_780),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_803),
.B(n_828),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_752),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_742),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_808),
.B(n_741),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_868),
.A2(n_738),
.B(n_743),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_848),
.B(n_849),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_753),
.Y(n_912)
);

AOI21x1_ASAP7_75t_SL g913 ( 
.A1(n_757),
.A2(n_826),
.B(n_785),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_786),
.A2(n_784),
.B(n_835),
.C(n_839),
.Y(n_914)
);

AO31x2_ASAP7_75t_L g915 ( 
.A1(n_746),
.A2(n_832),
.A3(n_793),
.B(n_773),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_802),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_817),
.A2(n_820),
.B(n_816),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_780),
.A2(n_854),
.B(n_850),
.C(n_858),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_857),
.B(n_759),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_824),
.Y(n_920)
);

AOI21x1_ASAP7_75t_SL g921 ( 
.A1(n_795),
.A2(n_792),
.B(n_776),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_824),
.Y(n_922)
);

AOI221xp5_ASAP7_75t_L g923 ( 
.A1(n_837),
.A2(n_827),
.B1(n_834),
.B2(n_795),
.C(n_747),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_796),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_836),
.B(n_758),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_796),
.B(n_765),
.Y(n_926)
);

AOI21x1_ASAP7_75t_L g927 ( 
.A1(n_781),
.A2(n_779),
.B(n_777),
.Y(n_927)
);

OAI21xp33_ASAP7_75t_L g928 ( 
.A1(n_838),
.A2(n_841),
.B(n_824),
.Y(n_928)
);

BUFx12f_ASAP7_75t_L g929 ( 
.A(n_852),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_805),
.Y(n_930)
);

INVx5_ASAP7_75t_L g931 ( 
.A(n_744),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_772),
.A2(n_789),
.B(n_744),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_788),
.A2(n_791),
.B(n_739),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_797),
.A2(n_806),
.B(n_814),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_765),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_790),
.A2(n_853),
.B1(n_806),
.B2(n_797),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_790),
.A2(n_853),
.B(n_870),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_818),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_751),
.Y(n_939)
);

AOI21xp33_ASAP7_75t_L g940 ( 
.A1(n_813),
.A2(n_840),
.B(n_855),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_851),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_855),
.A2(n_860),
.B(n_819),
.C(n_845),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_855),
.A2(n_860),
.B(n_819),
.C(n_845),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_845),
.B(n_866),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_806),
.B(n_824),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_845),
.B(n_866),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_763),
.A2(n_770),
.B(n_764),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_752),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_742),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_763),
.A2(n_770),
.B(n_764),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_763),
.A2(n_770),
.B(n_764),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_763),
.A2(n_770),
.B(n_764),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_851),
.Y(n_953)
);

OAI21x1_ASAP7_75t_L g954 ( 
.A1(n_763),
.A2(n_770),
.B(n_764),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_736),
.B(n_851),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_813),
.B(n_601),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_822),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_855),
.B(n_860),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_845),
.B(n_866),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_752),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_845),
.B(n_866),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_855),
.A2(n_860),
.B1(n_866),
.B2(n_845),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_845),
.B(n_866),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_851),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_763),
.A2(n_770),
.B(n_764),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_845),
.B(n_866),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_855),
.A2(n_860),
.B(n_819),
.C(n_845),
.Y(n_967)
);

AO31x2_ASAP7_75t_L g968 ( 
.A1(n_760),
.A2(n_860),
.A3(n_855),
.B(n_737),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_783),
.B(n_456),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_855),
.A2(n_860),
.B(n_819),
.C(n_845),
.Y(n_970)
);

AND3x4_ASAP7_75t_L g971 ( 
.A(n_861),
.B(n_719),
.C(n_865),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_766),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_845),
.B(n_866),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_845),
.B(n_866),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_736),
.B(n_851),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_766),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_855),
.A2(n_860),
.B(n_819),
.C(n_845),
.Y(n_977)
);

AOI21xp33_ASAP7_75t_L g978 ( 
.A1(n_813),
.A2(n_840),
.B(n_855),
.Y(n_978)
);

NAND3x1_ASAP7_75t_L g979 ( 
.A(n_838),
.B(n_834),
.C(n_813),
.Y(n_979)
);

NAND2x1_ASAP7_75t_SL g980 ( 
.A(n_749),
.B(n_716),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_742),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_855),
.B(n_860),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_845),
.B(n_866),
.Y(n_983)
);

AO21x1_ASAP7_75t_L g984 ( 
.A1(n_855),
.A2(n_860),
.B(n_864),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_855),
.A2(n_860),
.B1(n_866),
.B2(n_845),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_845),
.B(n_866),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_874),
.B(n_944),
.Y(n_987)
);

AO32x1_ASAP7_75t_L g988 ( 
.A1(n_962),
.A2(n_985),
.A3(n_957),
.B1(n_913),
.B2(n_897),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_956),
.B(n_893),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_929),
.Y(n_990)
);

CKINVDCx8_ASAP7_75t_R g991 ( 
.A(n_930),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_893),
.A2(n_986),
.B1(n_946),
.B2(n_983),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_896),
.A2(n_895),
.B1(n_956),
.B2(n_971),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_959),
.B(n_961),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_884),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_963),
.B(n_966),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_973),
.B(n_974),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_885),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_887),
.A2(n_888),
.B(n_886),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_L g1000 ( 
.A(n_889),
.B(n_880),
.C(n_895),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_903),
.B(n_892),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_875),
.B(n_942),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_884),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_955),
.B(n_975),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_907),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_904),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_971),
.A2(n_906),
.B1(n_891),
.B2(n_899),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_SL g1008 ( 
.A1(n_905),
.A2(n_890),
.B(n_977),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_875),
.A2(n_970),
.B1(n_967),
.B2(n_943),
.Y(n_1009)
);

AO21x1_ASAP7_75t_L g1010 ( 
.A1(n_958),
.A2(n_982),
.B(n_905),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_906),
.B(n_964),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_942),
.B(n_943),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_967),
.B(n_970),
.Y(n_1013)
);

INVx3_ASAP7_75t_R g1014 ( 
.A(n_938),
.Y(n_1014)
);

INVxp67_ASAP7_75t_SL g1015 ( 
.A(n_941),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_977),
.A2(n_958),
.B1(n_982),
.B2(n_909),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_953),
.B(n_941),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_876),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_929),
.Y(n_1019)
);

NOR2xp67_ASAP7_75t_SL g1020 ( 
.A(n_969),
.B(n_931),
.Y(n_1020)
);

INVx3_ASAP7_75t_SL g1021 ( 
.A(n_916),
.Y(n_1021)
);

AND2x2_ASAP7_75t_SL g1022 ( 
.A(n_925),
.B(n_923),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_984),
.B(n_914),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_972),
.Y(n_1024)
);

BUFx4_ASAP7_75t_SL g1025 ( 
.A(n_907),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_SL g1026 ( 
.A(n_931),
.B(n_936),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_877),
.A2(n_879),
.B(n_910),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_948),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_919),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_911),
.B(n_918),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_914),
.B(n_878),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_878),
.B(n_968),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_934),
.B(n_945),
.Y(n_1033)
);

CKINVDCx8_ASAP7_75t_R g1034 ( 
.A(n_945),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_912),
.B(n_900),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_938),
.B(n_900),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_976),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_957),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_881),
.A2(n_902),
.B1(n_928),
.B2(n_924),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_976),
.B(n_945),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_935),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_L g1042 ( 
.A1(n_894),
.A2(n_939),
.B1(n_920),
.B2(n_922),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_878),
.B(n_968),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_980),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_878),
.B(n_968),
.Y(n_1045)
);

INVx6_ASAP7_75t_SL g1046 ( 
.A(n_948),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_876),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_968),
.B(n_935),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_979),
.A2(n_931),
.B1(n_926),
.B2(n_922),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_931),
.Y(n_1050)
);

AOI21xp33_ASAP7_75t_SL g1051 ( 
.A1(n_937),
.A2(n_979),
.B(n_933),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_920),
.B(n_960),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_960),
.A2(n_882),
.B1(n_949),
.B2(n_981),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_908),
.B(n_981),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_882),
.A2(n_949),
.B1(n_981),
.B2(n_908),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_908),
.Y(n_1056)
);

CKINVDCx8_ASAP7_75t_R g1057 ( 
.A(n_981),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_SL g1058 ( 
.A1(n_932),
.A2(n_913),
.B(n_921),
.C(n_901),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_915),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_SL g1060 ( 
.A(n_927),
.B(n_917),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_883),
.B(n_947),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_950),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_951),
.Y(n_1063)
);

AOI221x1_ASAP7_75t_L g1064 ( 
.A1(n_965),
.A2(n_860),
.B1(n_855),
.B2(n_978),
.C(n_940),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_952),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_954),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_884),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_945),
.B(n_806),
.Y(n_1068)
);

NAND2x1p5_ASAP7_75t_L g1069 ( 
.A(n_931),
.B(n_945),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_874),
.B(n_944),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_969),
.B(n_736),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_904),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_907),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_934),
.B(n_713),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_873),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_969),
.Y(n_1076)
);

INVxp67_ASAP7_75t_SL g1077 ( 
.A(n_941),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_893),
.A2(n_840),
.B1(n_804),
.B2(n_855),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_969),
.B(n_953),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_887),
.A2(n_888),
.B(n_886),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_969),
.Y(n_1081)
);

BUFx12f_ASAP7_75t_L g1082 ( 
.A(n_929),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_969),
.B(n_736),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_874),
.B(n_944),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_969),
.Y(n_1085)
);

CKINVDCx6p67_ASAP7_75t_R g1086 ( 
.A(n_929),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_929),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_874),
.B(n_944),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_945),
.B(n_806),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_873),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_907),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_907),
.Y(n_1092)
);

INVxp67_ASAP7_75t_SL g1093 ( 
.A(n_941),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_955),
.B(n_975),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_884),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_884),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_893),
.B(n_813),
.C(n_601),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_874),
.B(n_944),
.Y(n_1098)
);

INVx3_ASAP7_75t_SL g1099 ( 
.A(n_969),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_893),
.A2(n_860),
.B1(n_855),
.B2(n_874),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_893),
.A2(n_860),
.B1(n_855),
.B2(n_874),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_969),
.B(n_736),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_956),
.B(n_601),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_887),
.A2(n_888),
.B(n_898),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_969),
.B(n_953),
.Y(n_1105)
);

INVx6_ASAP7_75t_L g1106 ( 
.A(n_1018),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_1033),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_1018),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1035),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_998),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_993),
.B(n_989),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1075),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_SL g1113 ( 
.A1(n_1010),
.A2(n_1048),
.B(n_1051),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_987),
.A2(n_996),
.B1(n_1084),
.B2(n_1098),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1090),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1000),
.A2(n_1078),
.B1(n_1022),
.B2(n_1097),
.Y(n_1116)
);

INVx6_ASAP7_75t_L g1117 ( 
.A(n_1018),
.Y(n_1117)
);

OAI22xp33_ASAP7_75t_SL g1118 ( 
.A1(n_1001),
.A2(n_1007),
.B1(n_992),
.B2(n_1070),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1100),
.A2(n_1101),
.B1(n_1103),
.B2(n_1009),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_SL g1120 ( 
.A1(n_1009),
.A2(n_1101),
.B1(n_1100),
.B2(n_1016),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1018),
.Y(n_1121)
);

BUFx8_ASAP7_75t_L g1122 ( 
.A(n_990),
.Y(n_1122)
);

CKINVDCx11_ASAP7_75t_R g1123 ( 
.A(n_1019),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_1047),
.Y(n_1124)
);

BUFx2_ASAP7_75t_SL g1125 ( 
.A(n_1005),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1033),
.B(n_1068),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1050),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1033),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1079),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1105),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_SL g1131 ( 
.A1(n_987),
.A2(n_1088),
.B1(n_1070),
.B2(n_1084),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1047),
.Y(n_1132)
);

CKINVDCx6p67_ASAP7_75t_R g1133 ( 
.A(n_1021),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_1016),
.A2(n_992),
.B1(n_1012),
.B2(n_1002),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1001),
.B(n_994),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1099),
.A2(n_1004),
.B1(n_1094),
.B2(n_1012),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1047),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_1011),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_1047),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1041),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1029),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_994),
.A2(n_1088),
.B1(n_1098),
.B2(n_997),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1071),
.A2(n_1083),
.B1(n_1102),
.B2(n_997),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1036),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1006),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_1082),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_996),
.B(n_1076),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1015),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1077),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_999),
.A2(n_1080),
.B(n_1027),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1050),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1069),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1061),
.A2(n_1065),
.B(n_1104),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1013),
.B(n_1023),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1063),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1093),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1023),
.A2(n_1059),
.B1(n_1085),
.B2(n_1081),
.Y(n_1157)
);

BUFx10_ASAP7_75t_L g1158 ( 
.A(n_1028),
.Y(n_1158)
);

BUFx2_ASAP7_75t_R g1159 ( 
.A(n_991),
.Y(n_1159)
);

INVx6_ASAP7_75t_L g1160 ( 
.A(n_1089),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_1086),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1064),
.A2(n_1045),
.B(n_1032),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1048),
.Y(n_1163)
);

OAI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1074),
.A2(n_1072),
.B1(n_1044),
.B2(n_1034),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1089),
.B(n_1040),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1030),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1062),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1017),
.B(n_1052),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1054),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1008),
.B(n_1074),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1066),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1042),
.A2(n_1039),
.B1(n_1031),
.B2(n_1053),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1031),
.B(n_1073),
.Y(n_1173)
);

BUFx2_ASAP7_75t_SL g1174 ( 
.A(n_1091),
.Y(n_1174)
);

BUFx4f_ASAP7_75t_L g1175 ( 
.A(n_1069),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_1020),
.B(n_1096),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_1092),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1025),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1049),
.A2(n_1087),
.B1(n_995),
.B2(n_1003),
.Y(n_1179)
);

NOR2x1_ASAP7_75t_R g1180 ( 
.A(n_1056),
.B(n_1014),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1056),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1032),
.A2(n_1045),
.B(n_1043),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1024),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1026),
.A2(n_1096),
.B1(n_1037),
.B2(n_1095),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1057),
.A2(n_1067),
.B1(n_1037),
.B2(n_1055),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_R g1186 ( 
.A(n_1058),
.B(n_988),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_988),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_988),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1046),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1060),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1046),
.A2(n_989),
.B1(n_813),
.B2(n_987),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1018),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_989),
.B(n_987),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_989),
.A2(n_893),
.B1(n_813),
.B2(n_840),
.Y(n_1194)
);

CKINVDCx11_ASAP7_75t_R g1195 ( 
.A(n_1019),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1035),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1038),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1025),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_989),
.A2(n_813),
.B1(n_994),
.B2(n_987),
.Y(n_1199)
);

INVxp33_ASAP7_75t_L g1200 ( 
.A(n_1004),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1035),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1035),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1025),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1050),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1035),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1008),
.B(n_1033),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_998),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1035),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1050),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1035),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1038),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1135),
.B(n_1193),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1135),
.B(n_1154),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1148),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1129),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1199),
.B(n_1114),
.Y(n_1216)
);

OR2x6_ASAP7_75t_L g1217 ( 
.A(n_1206),
.B(n_1170),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1149),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1182),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1154),
.B(n_1120),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1155),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1130),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1163),
.B(n_1111),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1182),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1200),
.B(n_1191),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1162),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1156),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1162),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1162),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1187),
.A2(n_1188),
.A3(n_1166),
.B(n_1155),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1206),
.Y(n_1231)
);

BUFx2_ASAP7_75t_R g1232 ( 
.A(n_1198),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1113),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1113),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1110),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1142),
.B(n_1147),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1194),
.A2(n_1119),
.B(n_1116),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1107),
.B(n_1128),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1131),
.B(n_1143),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1206),
.B(n_1134),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1206),
.B(n_1173),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1153),
.Y(n_1242)
);

OR2x6_ASAP7_75t_L g1243 ( 
.A(n_1170),
.B(n_1150),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1170),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1207),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1167),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1171),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1145),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1170),
.B(n_1144),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1200),
.B(n_1126),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1190),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1172),
.B(n_1176),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1133),
.A2(n_1179),
.B1(n_1138),
.B2(n_1164),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1118),
.A2(n_1175),
.B(n_1141),
.Y(n_1254)
);

CKINVDCx12_ASAP7_75t_R g1255 ( 
.A(n_1180),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1145),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1186),
.A2(n_1211),
.B(n_1197),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1112),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1176),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1115),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1186),
.A2(n_1169),
.B(n_1183),
.Y(n_1261)
);

INVx5_ASAP7_75t_L g1262 ( 
.A(n_1106),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1140),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1109),
.Y(n_1264)
);

NAND2x1_ASAP7_75t_L g1265 ( 
.A(n_1106),
.B(n_1117),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1168),
.B(n_1133),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1196),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1201),
.Y(n_1268)
);

BUFx12f_ASAP7_75t_L g1269 ( 
.A(n_1123),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1202),
.B(n_1210),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1205),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1208),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1136),
.A2(n_1185),
.B(n_1184),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1226),
.B(n_1157),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1243),
.B(n_1152),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1242),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1244),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1228),
.B(n_1165),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1221),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1247),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1236),
.B(n_1152),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_L g1282 ( 
.A(n_1259),
.B(n_1192),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1239),
.B(n_1160),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1229),
.B(n_1165),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1216),
.B(n_1181),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1257),
.B(n_1165),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1257),
.B(n_1177),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1223),
.B(n_1209),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1257),
.B(n_1230),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1237),
.A2(n_1195),
.B1(n_1123),
.B2(n_1146),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1252),
.A2(n_1175),
.B1(n_1160),
.B2(n_1203),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1225),
.A2(n_1195),
.B1(n_1146),
.B2(n_1160),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1219),
.B(n_1174),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1253),
.B(n_1160),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1213),
.B(n_1209),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1213),
.B(n_1151),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1241),
.B(n_1224),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1224),
.B(n_1125),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1244),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1243),
.B(n_1204),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1247),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1223),
.B(n_1127),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1266),
.B(n_1159),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1246),
.B(n_1127),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1273),
.B(n_1254),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1261),
.B(n_1108),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1281),
.B(n_1215),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1294),
.A2(n_1240),
.B1(n_1252),
.B2(n_1231),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1281),
.B(n_1222),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1305),
.B(n_1259),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1294),
.A2(n_1240),
.B1(n_1252),
.B2(n_1231),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1290),
.A2(n_1220),
.B1(n_1252),
.B2(n_1212),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1297),
.B(n_1238),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1283),
.B(n_1269),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1279),
.Y(n_1315)
);

OAI21xp33_ASAP7_75t_L g1316 ( 
.A1(n_1290),
.A2(n_1220),
.B(n_1252),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1291),
.B(n_1259),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1288),
.B(n_1235),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1283),
.B(n_1269),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1291),
.B(n_1262),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1302),
.B(n_1245),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1292),
.B(n_1251),
.C(n_1248),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1286),
.B(n_1249),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1295),
.B(n_1263),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1292),
.B(n_1262),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1286),
.B(n_1249),
.Y(n_1326)
);

OAI221xp5_ASAP7_75t_L g1327 ( 
.A1(n_1285),
.A2(n_1265),
.B1(n_1256),
.B2(n_1217),
.C(n_1234),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1274),
.A2(n_1231),
.B1(n_1217),
.B2(n_1250),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_L g1329 ( 
.A(n_1285),
.B(n_1251),
.C(n_1270),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1303),
.A2(n_1217),
.B1(n_1175),
.B2(n_1231),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_R g1331 ( 
.A(n_1274),
.B(n_1198),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1293),
.B(n_1258),
.C(n_1260),
.Y(n_1332)
);

OAI221xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1274),
.A2(n_1217),
.B1(n_1250),
.B2(n_1234),
.C(n_1233),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1278),
.B(n_1217),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1296),
.B(n_1280),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1284),
.B(n_1261),
.Y(n_1336)
);

NAND3xp33_ASAP7_75t_L g1337 ( 
.A(n_1293),
.B(n_1298),
.C(n_1260),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1282),
.B(n_1262),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1293),
.B(n_1298),
.C(n_1258),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1296),
.B(n_1271),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1282),
.B(n_1262),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1280),
.A2(n_1227),
.B1(n_1214),
.B2(n_1218),
.Y(n_1342)
);

NAND3xp33_ASAP7_75t_L g1343 ( 
.A(n_1298),
.B(n_1268),
.C(n_1264),
.Y(n_1343)
);

OAI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1299),
.A2(n_1265),
.B1(n_1233),
.B2(n_1189),
.C(n_1267),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_L g1345 ( 
.A(n_1304),
.B(n_1214),
.C(n_1218),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1301),
.B(n_1272),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1336),
.B(n_1289),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1337),
.B(n_1289),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1315),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1315),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1344),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1337),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1323),
.B(n_1326),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1339),
.B(n_1346),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1339),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1326),
.B(n_1287),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1334),
.B(n_1276),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1310),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1307),
.B(n_1309),
.Y(n_1359)
);

NOR2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1322),
.B(n_1244),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1327),
.B(n_1272),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1332),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1332),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1343),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1313),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1329),
.B(n_1301),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1343),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1335),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1340),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1342),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1329),
.B(n_1277),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1349),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1349),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1356),
.B(n_1300),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1356),
.B(n_1300),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1349),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1358),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1361),
.A2(n_1316),
.B1(n_1320),
.B2(n_1312),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1356),
.B(n_1300),
.Y(n_1379)
);

NAND2xp67_ASAP7_75t_L g1380 ( 
.A(n_1366),
.B(n_1122),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1371),
.B(n_1338),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1358),
.B(n_1318),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1350),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1350),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1352),
.B(n_1322),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1357),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1350),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1360),
.B(n_1341),
.Y(n_1388)
);

INVxp67_ASAP7_75t_SL g1389 ( 
.A(n_1371),
.Y(n_1389)
);

NOR3x1_ASAP7_75t_L g1390 ( 
.A(n_1352),
.B(n_1325),
.C(n_1317),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1350),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1351),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1360),
.B(n_1345),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1348),
.B(n_1324),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1356),
.B(n_1275),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1359),
.B(n_1314),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1360),
.B(n_1345),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1353),
.B(n_1275),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1348),
.B(n_1321),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1370),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1348),
.B(n_1306),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1357),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1365),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1370),
.B(n_1306),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1365),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1370),
.B(n_1306),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1353),
.B(n_1275),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1400),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1383),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1404),
.B(n_1352),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1385),
.B(n_1351),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1372),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1383),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1404),
.B(n_1355),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1392),
.B(n_1377),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1396),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1372),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1380),
.B(n_1319),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1381),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1382),
.B(n_1351),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1378),
.B(n_1351),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1373),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1390),
.B(n_1361),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1390),
.B(n_1355),
.Y(n_1424)
);

NOR2x1_ASAP7_75t_L g1425 ( 
.A(n_1393),
.B(n_1362),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1406),
.B(n_1355),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1398),
.B(n_1353),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1373),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1388),
.Y(n_1429)
);

OAI31xp33_ASAP7_75t_L g1430 ( 
.A1(n_1393),
.A2(n_1316),
.A3(n_1362),
.B(n_1363),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1407),
.B(n_1353),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1393),
.B(n_1368),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1397),
.B(n_1368),
.Y(n_1433)
);

AOI32xp33_ASAP7_75t_L g1434 ( 
.A1(n_1397),
.A2(n_1362),
.A3(n_1363),
.B1(n_1364),
.B2(n_1367),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1395),
.B(n_1347),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1381),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1395),
.B(n_1374),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1386),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1388),
.Y(n_1439)
);

NOR3xp33_ASAP7_75t_L g1440 ( 
.A(n_1389),
.B(n_1312),
.C(n_1363),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1397),
.B(n_1369),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1376),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1384),
.A2(n_1367),
.B(n_1364),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1388),
.B(n_1386),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1376),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1374),
.B(n_1347),
.Y(n_1446)
);

NAND2x1_ASAP7_75t_L g1447 ( 
.A(n_1402),
.B(n_1365),
.Y(n_1447)
);

AOI21xp33_ASAP7_75t_L g1448 ( 
.A1(n_1406),
.A2(n_1367),
.B(n_1364),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1399),
.B(n_1354),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1443),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1423),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1449),
.B(n_1399),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1443),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1434),
.B(n_1375),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1425),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_1411),
.Y(n_1456)
);

NOR2x1p5_ASAP7_75t_L g1457 ( 
.A(n_1436),
.B(n_1203),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1429),
.B(n_1381),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1421),
.A2(n_1440),
.B1(n_1424),
.B2(n_1420),
.Y(n_1459)
);

AND2x4_ASAP7_75t_SL g1460 ( 
.A(n_1444),
.B(n_1403),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1439),
.B(n_1444),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1408),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1430),
.B(n_1375),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1415),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1448),
.B(n_1441),
.Y(n_1465)
);

AND2x4_ASAP7_75t_SL g1466 ( 
.A(n_1444),
.B(n_1403),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1446),
.B(n_1379),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1432),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1412),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1418),
.B(n_1122),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1443),
.A2(n_1391),
.B(n_1384),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1419),
.Y(n_1472)
);

NOR2x1_ASAP7_75t_L g1473 ( 
.A(n_1419),
.B(n_1401),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1433),
.B(n_1379),
.Y(n_1474)
);

OR2x6_ASAP7_75t_L g1475 ( 
.A(n_1447),
.B(n_1380),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1412),
.Y(n_1476)
);

AND3x2_ASAP7_75t_L g1477 ( 
.A(n_1417),
.B(n_1178),
.C(n_1189),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1447),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1449),
.B(n_1122),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1427),
.B(n_1354),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1410),
.B(n_1161),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1446),
.B(n_1402),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1427),
.B(n_1405),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1438),
.A2(n_1311),
.B1(n_1308),
.B2(n_1330),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1409),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1469),
.Y(n_1486)
);

OAI21xp33_ASAP7_75t_L g1487 ( 
.A1(n_1459),
.A2(n_1414),
.B(n_1410),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1455),
.B(n_1438),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1471),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1455),
.Y(n_1490)
);

OAI322xp33_ASAP7_75t_L g1491 ( 
.A1(n_1459),
.A2(n_1414),
.A3(n_1426),
.B1(n_1354),
.B2(n_1401),
.C1(n_1366),
.C2(n_1428),
.Y(n_1491)
);

AOI21xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1479),
.A2(n_1426),
.B(n_1232),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1469),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1456),
.B(n_1431),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1476),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1456),
.B(n_1431),
.Y(n_1496)
);

OAI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1463),
.A2(n_1331),
.B(n_1333),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1461),
.B(n_1437),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1476),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1461),
.B(n_1437),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1462),
.Y(n_1501)
);

AOI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1451),
.A2(n_1422),
.B(n_1417),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1464),
.B(n_1481),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1462),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1485),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1485),
.Y(n_1506)
);

NAND2xp33_ASAP7_75t_SL g1507 ( 
.A(n_1457),
.B(n_1161),
.Y(n_1507)
);

INVxp67_ASAP7_75t_SL g1508 ( 
.A(n_1457),
.Y(n_1508)
);

INVxp67_ASAP7_75t_L g1509 ( 
.A(n_1472),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1484),
.A2(n_1394),
.B1(n_1435),
.B2(n_1365),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1464),
.B(n_1435),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1509),
.B(n_1468),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1507),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1490),
.B(n_1472),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1499),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1488),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1511),
.B(n_1465),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1499),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1492),
.A2(n_1454),
.B(n_1470),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1510),
.A2(n_1465),
.B1(n_1475),
.B2(n_1473),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1505),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1498),
.B(n_1458),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1494),
.B(n_1452),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1506),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1498),
.B(n_1458),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1486),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1488),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1507),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1508),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1493),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1500),
.B(n_1477),
.Y(n_1531)
);

AO21x1_ASAP7_75t_L g1532 ( 
.A1(n_1520),
.A2(n_1489),
.B(n_1453),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1513),
.A2(n_1491),
.B1(n_1487),
.B2(n_1502),
.C(n_1501),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1516),
.Y(n_1534)
);

NOR2x1_ASAP7_75t_L g1535 ( 
.A(n_1514),
.B(n_1504),
.Y(n_1535)
);

AND3x1_ASAP7_75t_L g1536 ( 
.A(n_1519),
.B(n_1503),
.C(n_1497),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1529),
.A2(n_1473),
.B(n_1488),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1528),
.A2(n_1513),
.B1(n_1525),
.B2(n_1531),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1522),
.A2(n_1496),
.B1(n_1475),
.B2(n_1500),
.Y(n_1539)
);

NAND3xp33_ASAP7_75t_SL g1540 ( 
.A(n_1512),
.B(n_1452),
.C(n_1450),
.Y(n_1540)
);

OAI322xp33_ASAP7_75t_L g1541 ( 
.A1(n_1517),
.A2(n_1495),
.A3(n_1453),
.B1(n_1450),
.B2(n_1489),
.C1(n_1485),
.C2(n_1478),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_SL g1542 ( 
.A1(n_1527),
.A2(n_1478),
.B(n_1453),
.C(n_1450),
.Y(n_1542)
);

AOI211x1_ASAP7_75t_SL g1543 ( 
.A1(n_1517),
.A2(n_1474),
.B(n_1480),
.C(n_1409),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1538),
.B(n_1525),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_L g1545 ( 
.A(n_1540),
.B(n_1541),
.Y(n_1545)
);

NOR2xp67_ASAP7_75t_L g1546 ( 
.A(n_1534),
.B(n_1537),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1535),
.Y(n_1547)
);

AO22x2_ASAP7_75t_L g1548 ( 
.A1(n_1539),
.A2(n_1526),
.B1(n_1518),
.B2(n_1515),
.Y(n_1548)
);

NAND3xp33_ASAP7_75t_L g1549 ( 
.A(n_1533),
.B(n_1530),
.C(n_1524),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1532),
.B(n_1523),
.Y(n_1550)
);

NAND4xp75_ASAP7_75t_L g1551 ( 
.A(n_1536),
.B(n_1526),
.C(n_1521),
.D(n_1482),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1542),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1543),
.Y(n_1553)
);

OAI211xp5_ASAP7_75t_L g1554 ( 
.A1(n_1533),
.A2(n_1523),
.B(n_1482),
.C(n_1467),
.Y(n_1554)
);

NAND4xp75_ASAP7_75t_L g1555 ( 
.A(n_1532),
.B(n_1467),
.C(n_1483),
.D(n_1255),
.Y(n_1555)
);

NAND2x1p5_ASAP7_75t_L g1556 ( 
.A(n_1547),
.B(n_1255),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1545),
.A2(n_1475),
.B1(n_1460),
.B2(n_1466),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1546),
.B(n_1475),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1544),
.B(n_1475),
.Y(n_1559)
);

NAND3xp33_ASAP7_75t_SL g1560 ( 
.A(n_1550),
.B(n_1483),
.C(n_1158),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_SL g1561 ( 
.A(n_1549),
.B(n_1554),
.C(n_1552),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1557),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1561),
.B(n_1553),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1558),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1559),
.B(n_1551),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1556),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1560),
.Y(n_1567)
);

NAND4xp75_ASAP7_75t_L g1568 ( 
.A(n_1563),
.B(n_1555),
.C(n_1548),
.D(n_1442),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1564),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1566),
.B(n_1460),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1562),
.B(n_1548),
.Y(n_1571)
);

NAND3x1_ASAP7_75t_L g1572 ( 
.A(n_1563),
.B(n_1158),
.C(n_1422),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1569),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1568),
.Y(n_1574)
);

NAND5xp2_ASAP7_75t_L g1575 ( 
.A(n_1570),
.B(n_1565),
.C(n_1567),
.D(n_1158),
.E(n_1328),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1573),
.B(n_1571),
.Y(n_1576)
);

NAND4xp25_ASAP7_75t_SL g1577 ( 
.A(n_1576),
.B(n_1574),
.C(n_1575),
.D(n_1572),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1577),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1577),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1578),
.A2(n_1471),
.B(n_1466),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1579),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1580),
.A2(n_1413),
.B(n_1428),
.Y(n_1582)
);

AOI31xp33_ASAP7_75t_L g1583 ( 
.A1(n_1581),
.A2(n_1108),
.A3(n_1139),
.B(n_1124),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1582),
.A2(n_1471),
.B(n_1466),
.Y(n_1584)
);

AOI222xp33_ASAP7_75t_L g1585 ( 
.A1(n_1584),
.A2(n_1583),
.B1(n_1460),
.B2(n_1445),
.C1(n_1442),
.C2(n_1413),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_R g1586 ( 
.A1(n_1585),
.A2(n_1445),
.B1(n_1405),
.B2(n_1394),
.C(n_1387),
.Y(n_1586)
);

AOI211xp5_ASAP7_75t_L g1587 ( 
.A1(n_1586),
.A2(n_1137),
.B(n_1121),
.C(n_1132),
.Y(n_1587)
);


endmodule