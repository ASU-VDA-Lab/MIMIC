module fake_jpeg_11185_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_0),
.B(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_11),
.B(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_6),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_16),
.B1(n_17),
.B2(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_10),
.B2(n_17),
.Y(n_31)
);

OR2x4_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_28),
.B1(n_30),
.B2(n_26),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_24),
.B(n_37),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_34),
.Y(n_48)
);

NOR2xp67_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_45),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_33),
.C(n_39),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_32),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_32),
.Y(n_53)
);


endmodule