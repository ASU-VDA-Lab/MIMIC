module fake_jpeg_15293_n_254 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_27),
.Y(n_54)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_21),
.B1(n_32),
.B2(n_19),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_59),
.B1(n_64),
.B2(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_29),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_54),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_21),
.B1(n_27),
.B2(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_29),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_65),
.C(n_29),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_19),
.B1(n_26),
.B2(n_18),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_32),
.B1(n_18),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_23),
.B1(n_17),
.B2(n_22),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_17),
.B1(n_26),
.B2(n_31),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_0),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_31),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_29),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_73),
.B(n_64),
.Y(n_105)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_75),
.A2(n_79),
.B1(n_82),
.B2(n_46),
.Y(n_111)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_39),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_41),
.B1(n_40),
.B2(n_42),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_39),
.B(n_40),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_99),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_105),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_39),
.B(n_38),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_63),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_1),
.Y(n_139)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_52),
.A3(n_66),
.B1(n_65),
.B2(n_57),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

AO21x1_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_81),
.B(n_38),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_46),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_87),
.B1(n_91),
.B2(n_80),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_88),
.B1(n_86),
.B2(n_84),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_118),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_116),
.B1(n_95),
.B2(n_106),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_83),
.B1(n_52),
.B2(n_70),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_45),
.B1(n_72),
.B2(n_97),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_125),
.B1(n_137),
.B2(n_114),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_69),
.B1(n_77),
.B2(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_51),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_51),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_39),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_73),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_135),
.C(n_60),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_140),
.B(n_102),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_101),
.C(n_112),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_92),
.Y(n_149)
);

AO21x2_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_60),
.B(n_42),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_103),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_38),
.B(n_72),
.C(n_76),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_150),
.B1(n_160),
.B2(n_137),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_129),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_SL g145 ( 
.A1(n_139),
.A2(n_105),
.A3(n_111),
.B1(n_116),
.B2(n_95),
.C1(n_96),
.C2(n_7),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_15),
.C(n_14),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_96),
.B(n_102),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_29),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_60),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_107),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_156),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_107),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_161),
.C(n_133),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_120),
.B(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_125),
.B(n_20),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_1),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_2),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_2),
.B(n_3),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_173),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_171),
.B1(n_185),
.B2(n_137),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_180),
.C(n_184),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_182),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_134),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_183),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_137),
.C(n_119),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_124),
.B1(n_137),
.B2(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_170),
.A2(n_141),
.B1(n_150),
.B2(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_147),
.C(n_152),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_148),
.B1(n_137),
.B2(n_159),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_194),
.B1(n_121),
.B2(n_136),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_164),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_156),
.C(n_154),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_195),
.C(n_200),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_148),
.B1(n_142),
.B2(n_151),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_142),
.C(n_162),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_163),
.C(n_143),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_145),
.B(n_157),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_201),
.B(n_192),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_118),
.C(n_117),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_185),
.C(n_3),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_177),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_209),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_208),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_211),
.Y(n_220)
);

AOI31xp67_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_179),
.A3(n_176),
.B(n_178),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_179),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_215),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_200),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_2),
.C(n_3),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_202),
.B(n_193),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_223),
.B(n_205),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_187),
.B(n_198),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_4),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_190),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_228),
.C(n_4),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_195),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_227),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_216),
.B1(n_207),
.B2(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_231),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_220),
.B(n_4),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_235),
.C(n_232),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_6),
.C(n_7),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_219),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_6),
.B(n_9),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_9),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_234),
.A2(n_226),
.B1(n_222),
.B2(n_218),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_9),
.Y(n_247)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_241),
.B(n_219),
.C(n_239),
.D(n_10),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_245),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_6),
.C(n_7),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_10),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_12),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_12),
.B(n_13),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_252),
.B(n_249),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_45),
.Y(n_254)
);


endmodule