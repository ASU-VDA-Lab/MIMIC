module fake_jpeg_1143_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_SL g6 ( 
.A(n_5),
.Y(n_6)
);

INVx11_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_0),
.A2(n_4),
.B1(n_5),
.B2(n_3),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_6),
.B1(n_12),
.B2(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_13),
.Y(n_19)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_2),
.B(n_13),
.C(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_16),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_28),
.B(n_15),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_20),
.B(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_6),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_21),
.B(n_23),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_32),
.Y(n_35)
);

FAx1_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_24),
.CI(n_20),
.CON(n_31),
.SN(n_31)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_25),
.B(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.C(n_26),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_8),
.B(n_7),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_10),
.B(n_7),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_8),
.Y(n_38)
);

OA21x2_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_10),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_10),
.Y(n_41)
);


endmodule