module fake_jpeg_533_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_58),
.Y(n_64)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_55),
.Y(n_60)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_1),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_50),
.B1(n_43),
.B2(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_46),
.B1(n_43),
.B2(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_67),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_41),
.B1(n_45),
.B2(n_49),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_69),
.B1(n_54),
.B2(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_57),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_48),
.B1(n_47),
.B2(n_49),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_49),
.B(n_39),
.C(n_4),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_76),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_60),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_59),
.B1(n_4),
.B2(n_5),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_83),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_56),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_61),
.B(n_59),
.C(n_21),
.Y(n_84)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_71),
.B(n_76),
.C(n_8),
.D(n_9),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_88),
.B1(n_7),
.B2(n_8),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_29),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_9),
.Y(n_104)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_84),
.B(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_108),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_23),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_109),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_27),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_110),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_28),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_10),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_10),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_113),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_14),
.Y(n_114)
);

BUFx4f_ASAP7_75t_SL g116 ( 
.A(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_119),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_15),
.C(n_16),
.Y(n_122)
);

OA21x2_ASAP7_75t_SL g131 ( 
.A1(n_122),
.A2(n_127),
.B(n_22),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_103),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_106),
.B1(n_96),
.B2(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_133),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_117),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_36),
.B(n_31),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_125),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_35),
.B1(n_116),
.B2(n_120),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_115),
.C(n_124),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_137),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_138),
.B1(n_128),
.B2(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_140),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_144),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_134),
.Y(n_146)
);


endmodule