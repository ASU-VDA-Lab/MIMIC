module fake_jpeg_30279_n_542 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_542);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_11),
.B(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_58),
.Y(n_107)
);

HAxp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_1),
.CON(n_57),
.SN(n_57)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_57),
.B(n_70),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_28),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_77),
.Y(n_111)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_9),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_99),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_26),
.Y(n_99)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_51),
.Y(n_138)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_33),
.B1(n_30),
.B2(n_48),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_105),
.A2(n_159),
.B1(n_75),
.B2(n_81),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_109),
.B(n_114),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_29),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_124),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_29),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_61),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_132),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_61),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_37),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_147),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_40),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_144),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_74),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_51),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_50),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_153),
.B(n_155),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_59),
.B(n_50),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_55),
.A2(n_30),
.B1(n_33),
.B2(n_37),
.Y(n_159)
);

BUFx16f_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

BUFx12_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_88),
.B1(n_43),
.B2(n_102),
.Y(n_167)
);

AO22x2_ASAP7_75t_L g261 ( 
.A1(n_167),
.A2(n_210),
.B1(n_98),
.B2(n_97),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_45),
.B1(n_99),
.B2(n_94),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_168),
.A2(n_222),
.B1(n_45),
.B2(n_121),
.Y(n_237)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_171),
.Y(n_252)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_174),
.Y(n_236)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_177),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_178),
.Y(n_265)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_181),
.Y(n_278)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_182),
.Y(n_238)
);

CKINVDCx6p67_ASAP7_75t_R g183 ( 
.A(n_116),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_48),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_185),
.B(n_191),
.Y(n_275)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_111),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_202),
.Y(n_232)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_189),
.Y(n_269)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_190),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_107),
.B(n_21),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_22),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_193),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_21),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_194),
.B(n_197),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_40),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_214),
.Y(n_231)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_145),
.B(n_46),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_199),
.Y(n_279)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_133),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_166),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_203),
.B(n_205),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_123),
.A2(n_126),
.B1(n_156),
.B2(n_62),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_226),
.B1(n_125),
.B2(n_118),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_146),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_46),
.Y(n_206)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_143),
.Y(n_207)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_207),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

AO22x1_ASAP7_75t_SL g210 ( 
.A1(n_150),
.A2(n_63),
.B1(n_68),
.B2(n_69),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_210),
.A2(n_224),
.B1(n_118),
.B2(n_157),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_131),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_141),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_213),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_112),
.B(n_41),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_41),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_217),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_108),
.B(n_47),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_137),
.A2(n_45),
.B(n_22),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_218),
.A2(n_28),
.B(n_2),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_112),
.B(n_47),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_221),
.Y(n_259)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_220),
.A2(n_223),
.B1(n_225),
.B2(n_125),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_136),
.B(n_34),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_122),
.B(n_44),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_131),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_108),
.A2(n_90),
.B1(n_92),
.B2(n_95),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_122),
.B(n_54),
.C(n_78),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_45),
.C(n_136),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_229),
.B(n_237),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_170),
.A2(n_121),
.B1(n_110),
.B2(n_157),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_251),
.B1(n_276),
.B2(n_226),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g298 ( 
.A1(n_242),
.A2(n_253),
.B1(n_261),
.B2(n_225),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_94),
.Y(n_243)
);

NAND2x1_ASAP7_75t_L g322 ( 
.A(n_243),
.B(n_184),
.Y(n_322)
);

OAI22x1_ASAP7_75t_L g253 ( 
.A1(n_167),
.A2(n_160),
.B1(n_44),
.B2(n_96),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_175),
.B(n_9),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_SL g316 ( 
.A(n_257),
.B(n_14),
.C(n_15),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_115),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_260),
.B(n_266),
.C(n_270),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_177),
.A2(n_128),
.B1(n_127),
.B2(n_84),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_218),
.A2(n_152),
.B1(n_162),
.B2(n_150),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_264),
.A2(n_168),
.B1(n_213),
.B2(n_190),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_174),
.B(n_100),
.C(n_89),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_167),
.A2(n_30),
.B1(n_33),
.B2(n_93),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_272),
.B(n_229),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_195),
.B(n_162),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_199),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_216),
.B(n_11),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_227),
.A2(n_152),
.B1(n_91),
.B2(n_25),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_253),
.A2(n_210),
.B1(n_171),
.B2(n_204),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_281),
.A2(n_286),
.B1(n_316),
.B2(n_263),
.Y(n_333)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_228),
.Y(n_282)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_284),
.A2(n_292),
.B1(n_298),
.B2(n_328),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_208),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_285),
.B(n_287),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_180),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_169),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_288),
.B(n_294),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_289),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_172),
.B1(n_220),
.B2(n_193),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_290),
.A2(n_242),
.B1(n_271),
.B2(n_261),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_212),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_300),
.Y(n_340)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_293),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_231),
.B(n_207),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_188),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_306),
.Y(n_330)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_182),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_250),
.A2(n_181),
.B1(n_223),
.B2(n_183),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_246),
.B(n_178),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

AND2x6_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_184),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_308),
.A2(n_325),
.B(n_291),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_236),
.A2(n_223),
.B1(n_183),
.B2(n_200),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_309),
.A2(n_321),
.B1(n_323),
.B2(n_327),
.Y(n_360)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

BUFx12f_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_312),
.Y(n_348)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_196),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_319),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_259),
.B(n_178),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_318),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_255),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_231),
.B(n_201),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_320),
.B(n_325),
.Y(n_367)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

NAND2x1_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_243),
.Y(n_334)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_248),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_176),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_326),
.B(n_176),
.Y(n_368)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_333),
.B(n_338),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_SL g391 ( 
.A1(n_334),
.A2(n_289),
.B(n_305),
.Y(n_391)
);

XOR2x2_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_260),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_316),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_324),
.A2(n_263),
.B1(n_276),
.B2(n_243),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_283),
.A2(n_272),
.B(n_267),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_349),
.A2(n_350),
.B(n_335),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_292),
.A2(n_325),
.B(n_283),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_353),
.A2(n_356),
.B1(n_358),
.B2(n_370),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_284),
.A2(n_261),
.B1(n_243),
.B2(n_277),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_315),
.A2(n_261),
.B1(n_279),
.B2(n_189),
.Y(n_358)
);

OAI32xp33_ASAP7_75t_L g359 ( 
.A1(n_300),
.A2(n_257),
.A3(n_273),
.B1(n_233),
.B2(n_240),
.Y(n_359)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_290),
.A2(n_173),
.B1(n_280),
.B2(n_244),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_362),
.A2(n_364),
.B1(n_365),
.B2(n_304),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_363),
.B(n_367),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_298),
.A2(n_244),
.B1(n_238),
.B2(n_245),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_298),
.A2(n_238),
.B1(n_278),
.B2(n_241),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_324),
.A2(n_278),
.B1(n_10),
.B2(n_12),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_366),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_368),
.B(n_293),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_298),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_371),
.A2(n_394),
.B1(n_401),
.B2(n_366),
.Y(n_421)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

MAJx2_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_314),
.C(n_308),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_381),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_289),
.Y(n_375)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_332),
.Y(n_376)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_369),
.Y(n_377)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_299),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_380),
.B(n_384),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_367),
.B(n_286),
.C(n_322),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_382),
.B(n_334),
.C(n_359),
.Y(n_420)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_383),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_296),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_344),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_385),
.Y(n_406)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_387),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_388),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_355),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_389),
.B(n_397),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_391),
.A2(n_393),
.B1(n_395),
.B2(n_399),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_333),
.A2(n_328),
.B1(n_311),
.B2(n_327),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_339),
.A2(n_312),
.B1(n_303),
.B2(n_289),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_338),
.A2(n_356),
.B1(n_363),
.B2(n_358),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_330),
.B(n_312),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_398),
.A2(n_349),
.B(n_368),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_335),
.A2(n_323),
.B1(n_321),
.B2(n_310),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_370),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_337),
.B(n_1),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_404),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_332),
.B(n_1),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_403),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_331),
.B(n_1),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_3),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_348),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_407),
.B(n_417),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_415),
.A2(n_430),
.B(n_431),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_345),
.Y(n_419)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_419),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_427),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_421),
.A2(n_346),
.B1(n_4),
.B2(n_6),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_334),
.C(n_347),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_435),
.C(n_424),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_381),
.B(n_351),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_426),
.B(n_354),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_390),
.B(n_351),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_375),
.A2(n_344),
.B(n_360),
.Y(n_428)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_428),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_396),
.A2(n_353),
.B1(n_357),
.B2(n_347),
.Y(n_429)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_429),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_387),
.A2(n_398),
.B(n_392),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_385),
.B(n_341),
.Y(n_433)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_433),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_396),
.A2(n_372),
.B1(n_382),
.B2(n_395),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_372),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_376),
.B(n_329),
.C(n_352),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_440),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_441),
.A2(n_462),
.B1(n_425),
.B2(n_411),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_436),
.A2(n_379),
.B1(n_392),
.B2(n_393),
.Y(n_445)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_445),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_422),
.B(n_392),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_447),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_420),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_448),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_SL g449 ( 
.A(n_413),
.B(n_379),
.C(n_403),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_449),
.B(n_451),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_399),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_454),
.C(n_455),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_430),
.A2(n_377),
.B(n_388),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_452),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_436),
.A2(n_386),
.B1(n_383),
.B2(n_357),
.Y(n_453)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_329),
.C(n_352),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_401),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_409),
.Y(n_456)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_456),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_SL g457 ( 
.A(n_415),
.B(n_421),
.C(n_406),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_R g464 ( 
.A(n_457),
.B(n_458),
.Y(n_464)
);

XOR2x2_ASAP7_75t_L g458 ( 
.A(n_411),
.B(n_341),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_459),
.B(n_425),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_406),
.B(n_354),
.Y(n_460)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_460),
.Y(n_474)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_473),
.A2(n_470),
.B1(n_442),
.B2(n_474),
.Y(n_489)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_460),
.Y(n_475)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_475),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_445),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_462),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_438),
.B(n_412),
.C(n_423),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_478),
.B(n_454),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_461),
.Y(n_479)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_479),
.Y(n_498)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_437),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_481),
.Y(n_500)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_443),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_451),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_482),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_423),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_484),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_440),
.B(n_432),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_490),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_465),
.B(n_446),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_489),
.Y(n_507)
);

OAI322xp33_ASAP7_75t_L g488 ( 
.A1(n_484),
.A2(n_449),
.A3(n_418),
.B1(n_447),
.B2(n_441),
.C1(n_444),
.C2(n_439),
.Y(n_488)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_488),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_463),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_464),
.A2(n_458),
.B(n_455),
.C(n_450),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_494),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_467),
.B(n_476),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_483),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_444),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_473),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_469),
.B(n_410),
.Y(n_499)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_499),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_478),
.B(n_418),
.Y(n_501)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_501),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_467),
.C(n_476),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_503),
.B(n_504),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_477),
.C(n_470),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_487),
.B(n_477),
.C(n_471),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_509),
.C(n_515),
.Y(n_516)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_500),
.Y(n_511)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_511),
.Y(n_517)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_485),
.Y(n_512)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_512),
.Y(n_521)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_495),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_514),
.B(n_432),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_489),
.C(n_491),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_518),
.B(n_519),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_506),
.B(n_494),
.C(n_498),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_522),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_497),
.C(n_471),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_510),
.A2(n_464),
.B(n_492),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_524),
.A2(n_525),
.B(n_497),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_468),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_502),
.C(n_509),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_527),
.A2(n_528),
.B(n_516),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_525),
.A2(n_466),
.B(n_510),
.Y(n_528)
);

AOI322xp5_ASAP7_75t_L g532 ( 
.A1(n_529),
.A2(n_531),
.A3(n_519),
.B1(n_492),
.B2(n_521),
.C1(n_507),
.C2(n_414),
.Y(n_532)
);

AOI321xp33_ASAP7_75t_L g531 ( 
.A1(n_517),
.A2(n_492),
.A3(n_507),
.B1(n_412),
.B2(n_414),
.C(n_416),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_532),
.A2(n_533),
.B(n_534),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_526),
.B(n_472),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_533),
.A2(n_530),
.B(n_409),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_535),
.B(n_416),
.Y(n_537)
);

OAI311xp33_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_536),
.A3(n_456),
.B1(n_6),
.C1(n_7),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_3),
.C(n_4),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_4),
.B(n_6),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_6),
.Y(n_541)
);

AO21x1_ASAP7_75t_L g542 ( 
.A1(n_541),
.A2(n_7),
.B(n_8),
.Y(n_542)
);


endmodule