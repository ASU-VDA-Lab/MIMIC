module fake_jpeg_7853_n_38 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g19 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_2),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_11),
.C(n_6),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_17),
.B1(n_3),
.B2(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_29),
.Y(n_33)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_7),
.B1(n_9),
.B2(n_12),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_31),
.Y(n_37)
);

A2O1A1O1Ixp25_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_30),
.B(n_33),
.C(n_25),
.D(n_13),
.Y(n_38)
);


endmodule