module fake_netlist_1_7545_n_858 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_858);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_858;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_462;
wire n_232;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_522;
wire n_264;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_695;
wire n_650;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g107 ( .A(n_99), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_17), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_105), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_102), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_61), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_65), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_70), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_20), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_26), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_51), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_85), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_103), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_94), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_22), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g124 ( .A(n_59), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_27), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_28), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_23), .Y(n_127) );
BUFx10_ASAP7_75t_L g128 ( .A(n_64), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_24), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_26), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_101), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_100), .Y(n_132) );
INVx1_ASAP7_75t_SL g133 ( .A(n_5), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_15), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_62), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_13), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_93), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_15), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_21), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_9), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_86), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
INVx2_ASAP7_75t_SL g143 ( .A(n_48), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_4), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_37), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_57), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_1), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_97), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_74), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_104), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_120), .B(n_108), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_120), .B(n_0), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_143), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_107), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_143), .B(n_0), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_128), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_107), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_108), .B(n_1), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_126), .B(n_2), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_126), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_109), .B(n_2), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_124), .B(n_3), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_146), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_107), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_139), .B(n_3), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_128), .Y(n_166) );
BUFx12f_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_109), .B(n_4), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_107), .Y(n_169) );
BUFx12f_ASAP7_75t_L g170 ( .A(n_128), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_112), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_112), .B(n_5), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_113), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_162), .A2(n_136), .B1(n_123), .B2(n_125), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_164), .Y(n_175) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_152), .A2(n_139), .B1(n_144), .B2(n_129), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_168), .Y(n_177) );
OAI22xp33_ASAP7_75t_R g178 ( .A1(n_161), .A2(n_133), .B1(n_148), .B2(n_150), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_168), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_168), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_156), .B(n_150), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_151), .A2(n_130), .B1(n_127), .B2(n_147), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_151), .B(n_114), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_151), .B(n_115), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
AO22x2_ASAP7_75t_L g187 ( .A1(n_168), .A2(n_113), .B1(n_118), .B2(n_121), .Y(n_187) );
OA22x2_ASAP7_75t_L g188 ( .A1(n_160), .A2(n_140), .B1(n_138), .B2(n_145), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_168), .Y(n_189) );
INVxp67_ASAP7_75t_SL g190 ( .A(n_152), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_167), .Y(n_191) );
OAI22xp33_ASAP7_75t_L g192 ( .A1(n_152), .A2(n_134), .B1(n_148), .B2(n_142), .Y(n_192) );
OAI22xp33_ASAP7_75t_SL g193 ( .A1(n_166), .A2(n_142), .B1(n_141), .B2(n_118), .Y(n_193) );
AO22x2_ASAP7_75t_L g194 ( .A1(n_168), .A2(n_121), .B1(n_135), .B2(n_141), .Y(n_194) );
AO22x2_ASAP7_75t_L g195 ( .A1(n_168), .A2(n_135), .B1(n_7), .B2(n_8), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_160), .B(n_110), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_162), .A2(n_119), .B1(n_137), .B2(n_132), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_167), .B(n_107), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_160), .B(n_111), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_167), .B(n_116), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_167), .A2(n_149), .B1(n_131), .B2(n_122), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_167), .A2(n_117), .B1(n_107), .B2(n_8), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_170), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_170), .A2(n_6), .B1(n_10), .B2(n_11), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_170), .B(n_10), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_170), .B(n_11), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_170), .B(n_12), .Y(n_209) );
INVx1_ASAP7_75t_SL g210 ( .A(n_162), .Y(n_210) );
OR2x6_ASAP7_75t_L g211 ( .A(n_162), .B(n_12), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_168), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_173), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_156), .B(n_13), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_156), .B(n_14), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g216 ( .A1(n_158), .A2(n_14), .B1(n_16), .B2(n_17), .Y(n_216) );
AO22x2_ASAP7_75t_L g217 ( .A1(n_156), .A2(n_16), .B1(n_18), .B2(n_19), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_158), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_166), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_156), .B(n_24), .Y(n_220) );
INVxp33_ASAP7_75t_L g221 ( .A(n_196), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_213), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_213), .Y(n_223) );
OR2x2_ASAP7_75t_L g224 ( .A(n_210), .B(n_163), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_177), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_177), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_179), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_190), .B(n_158), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_175), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_179), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_180), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_184), .B(n_159), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
INVxp67_ASAP7_75t_SL g235 ( .A(n_189), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_196), .B(n_155), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_189), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_184), .B(n_159), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g239 ( .A(n_212), .B(n_173), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_183), .Y(n_240) );
XNOR2xp5_ASAP7_75t_L g241 ( .A(n_211), .B(n_163), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_212), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_183), .Y(n_243) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_187), .A2(n_173), .B(n_171), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_185), .B(n_159), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_211), .B(n_165), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_187), .Y(n_247) );
XOR2xp5_ASAP7_75t_L g248 ( .A(n_174), .B(n_165), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_211), .B(n_165), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_187), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_187), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_194), .Y(n_252) );
XNOR2x2_ASAP7_75t_L g253 ( .A(n_217), .B(n_161), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_194), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_200), .B(n_155), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_200), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_185), .B(n_155), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_194), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_198), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_194), .A2(n_173), .B(n_171), .Y(n_260) );
AND2x2_ASAP7_75t_SL g261 ( .A(n_214), .B(n_171), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_214), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_191), .B(n_161), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_214), .Y(n_264) );
XOR2xp5_ASAP7_75t_L g265 ( .A(n_174), .B(n_25), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_181), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_181), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_197), .B(n_153), .Y(n_268) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_207), .B(n_172), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_181), .Y(n_270) );
INVxp33_ASAP7_75t_L g271 ( .A(n_188), .Y(n_271) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_207), .B(n_172), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_195), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_211), .B(n_153), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_191), .B(n_172), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_186), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_197), .Y(n_277) );
AND2x6_ASAP7_75t_L g278 ( .A(n_208), .B(n_153), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_195), .Y(n_279) );
XOR2xp5_ASAP7_75t_L g280 ( .A(n_188), .B(n_25), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_186), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_195), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_244), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_222), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_222), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_228), .B(n_208), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_228), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_225), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_229), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_226), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_249), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_229), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_233), .B(n_209), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_233), .B(n_192), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_238), .B(n_209), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_246), .B(n_220), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_261), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_230), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_226), .Y(n_303) );
INVx3_ASAP7_75t_SL g304 ( .A(n_249), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_238), .B(n_195), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_245), .B(n_198), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_261), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_230), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_256), .B(n_182), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_245), .B(n_193), .Y(n_310) );
BUFx4f_ASAP7_75t_L g311 ( .A(n_261), .Y(n_311) );
INVx8_ASAP7_75t_L g312 ( .A(n_249), .Y(n_312) );
BUFx5_ASAP7_75t_L g313 ( .A(n_269), .Y(n_313) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_246), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_256), .B(n_176), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_249), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_260), .A2(n_220), .B(n_215), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_230), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_249), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_246), .B(n_198), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_246), .B(n_198), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_257), .B(n_201), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_240), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_247), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_227), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_269), .B(n_201), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_269), .B(n_272), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_241), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_272), .B(n_217), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_244), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_227), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_272), .B(n_188), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_274), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_290), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_312), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_312), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_288), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g338 ( .A(n_311), .B(n_247), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_314), .B(n_274), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_288), .Y(n_340) );
CKINVDCx6p67_ASAP7_75t_R g341 ( .A(n_304), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_291), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_313), .B(n_235), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_327), .B(n_224), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_313), .B(n_235), .Y(n_345) );
INVx8_ASAP7_75t_L g346 ( .A(n_312), .Y(n_346) );
OR2x6_ASAP7_75t_L g347 ( .A(n_312), .B(n_250), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_291), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_312), .B(n_250), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_236), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_290), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_290), .Y(n_353) );
INVx6_ASAP7_75t_L g354 ( .A(n_333), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_333), .Y(n_355) );
NOR2xp33_ASAP7_75t_SL g356 ( .A(n_311), .B(n_251), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_292), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_291), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_294), .B(n_274), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_313), .B(n_255), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_328), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_292), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_294), .B(n_333), .Y(n_364) );
AND2x6_ASAP7_75t_L g365 ( .A(n_301), .B(n_251), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g366 ( .A(n_352), .B(n_294), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_352), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_342), .Y(n_368) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_352), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_344), .B(n_248), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_335), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_342), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_359), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVxp67_ASAP7_75t_L g375 ( .A(n_359), .Y(n_375) );
BUFx4f_ASAP7_75t_SL g376 ( .A(n_341), .Y(n_376) );
CKINVDCx6p67_ASAP7_75t_R g377 ( .A(n_341), .Y(n_377) );
BUFx8_ASAP7_75t_L g378 ( .A(n_359), .Y(n_378) );
INVx4_ASAP7_75t_L g379 ( .A(n_346), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_346), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g382 ( .A(n_339), .B(n_294), .Y(n_382) );
INVx5_ASAP7_75t_SL g383 ( .A(n_341), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_339), .B(n_294), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_334), .B(n_286), .Y(n_385) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_346), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_346), .Y(n_389) );
BUFx12f_ASAP7_75t_L g390 ( .A(n_335), .Y(n_390) );
BUFx2_ASAP7_75t_R g391 ( .A(n_344), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_346), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_346), .Y(n_393) );
BUFx3_ASAP7_75t_L g394 ( .A(n_346), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_379), .B(n_335), .Y(n_395) );
INVx6_ASAP7_75t_L g396 ( .A(n_386), .Y(n_396) );
BUFx10_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_378), .A2(n_329), .B1(n_312), .B2(n_294), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_370), .A2(n_313), .B1(n_311), .B2(n_301), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_368), .Y(n_400) );
BUFx10_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_370), .A2(n_313), .B1(n_311), .B2(n_301), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_372), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_378), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_369), .A2(n_311), .B1(n_319), .B2(n_301), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_369), .A2(n_241), .B1(n_178), .B2(n_248), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_386), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_386), .Y(n_408) );
INVx8_ASAP7_75t_L g409 ( .A(n_386), .Y(n_409) );
CKINVDCx6p67_ASAP7_75t_R g410 ( .A(n_377), .Y(n_410) );
INVx4_ASAP7_75t_L g411 ( .A(n_377), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_369), .A2(n_311), .B1(n_319), .B2(n_301), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_376), .Y(n_413) );
INVx6_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
BUFx10_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_369), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_390), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_378), .A2(n_313), .B1(n_311), .B2(n_329), .Y(n_421) );
BUFx12f_ASAP7_75t_L g422 ( .A(n_378), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_373), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_371), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_379), .A2(n_313), .B1(n_329), .B2(n_178), .Y(n_426) );
INVx6_ASAP7_75t_L g427 ( .A(n_379), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_379), .A2(n_313), .B1(n_329), .B2(n_280), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_373), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_376), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_379), .A2(n_304), .B1(n_312), .B2(n_307), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_377), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_387), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_387), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_391), .A2(n_304), .B1(n_339), .B2(n_294), .Y(n_435) );
BUFx10_ASAP7_75t_L g436 ( .A(n_380), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_387), .A2(n_313), .B1(n_280), .B2(n_326), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_387), .A2(n_313), .B1(n_326), .B2(n_312), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_406), .B(n_219), .C(n_205), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_426), .A2(n_313), .B1(n_393), .B2(n_392), .Y(n_441) );
INVx5_ASAP7_75t_SL g442 ( .A(n_410), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_404), .A2(n_265), .B(n_305), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_400), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_422), .A2(n_313), .B1(n_393), .B2(n_392), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g446 ( .A1(n_422), .A2(n_393), .B1(n_392), .B2(n_389), .Y(n_446) );
INVxp33_ASAP7_75t_SL g447 ( .A(n_432), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_403), .B(n_305), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_413), .A2(n_328), .B1(n_265), .B2(n_362), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_423), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_437), .A2(n_313), .B1(n_393), .B2(n_392), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_403), .B(n_367), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_410), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_413), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_428), .A2(n_313), .B1(n_389), .B2(n_394), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_404), .A2(n_313), .B1(n_389), .B2(n_394), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_427), .A2(n_383), .B1(n_389), .B2(n_394), .Y(n_457) );
INVx2_ASAP7_75t_SL g458 ( .A(n_397), .Y(n_458) );
INVx5_ASAP7_75t_L g459 ( .A(n_409), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_399), .A2(n_313), .B1(n_394), .B2(n_312), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_418), .B(n_362), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_402), .A2(n_381), .B1(n_305), .B2(n_327), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_398), .A2(n_391), .B1(n_434), .B2(n_432), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_425), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_407), .Y(n_465) );
BUFx12f_ASAP7_75t_L g466 ( .A(n_411), .Y(n_466) );
OAI21xp33_ASAP7_75t_L g467 ( .A1(n_419), .A2(n_271), .B(n_217), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_427), .A2(n_383), .B1(n_366), .B2(n_253), .Y(n_468) );
OR2x2_ASAP7_75t_SL g469 ( .A(n_396), .B(n_371), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_427), .A2(n_383), .B1(n_366), .B2(n_253), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g471 ( .A1(n_434), .A2(n_366), .B1(n_380), .B2(n_382), .Y(n_471) );
OAI22xp33_ASAP7_75t_L g472 ( .A1(n_411), .A2(n_366), .B1(n_380), .B2(n_382), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_396), .A2(n_304), .B1(n_383), .B2(n_384), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_435), .A2(n_310), .B1(n_326), .B2(n_305), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_397), .Y(n_475) );
BUFx12f_ASAP7_75t_L g476 ( .A(n_411), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g477 ( .A1(n_424), .A2(n_217), .B(n_204), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_397), .Y(n_478) );
INVx4_ASAP7_75t_R g479 ( .A(n_433), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_409), .A2(n_381), .B1(n_327), .B2(n_365), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_401), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_409), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_409), .A2(n_381), .B1(n_365), .B2(n_339), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_396), .A2(n_304), .B1(n_383), .B2(n_384), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_396), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_401), .Y(n_486) );
CKINVDCx6p67_ASAP7_75t_R g487 ( .A(n_430), .Y(n_487) );
CKINVDCx11_ASAP7_75t_R g488 ( .A(n_430), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_401), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_421), .A2(n_365), .B1(n_339), .B2(n_335), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_416), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_407), .B(n_337), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_414), .A2(n_383), .B1(n_384), .B2(n_382), .Y(n_493) );
AOI222xp33_ASAP7_75t_L g494 ( .A1(n_417), .A2(n_310), .B1(n_332), .B2(n_326), .C1(n_277), .C2(n_268), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_407), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_438), .A2(n_365), .B1(n_336), .B2(n_335), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_427), .A2(n_414), .B1(n_350), .B2(n_361), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_405), .A2(n_365), .B1(n_336), .B2(n_335), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_424), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_414), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_412), .A2(n_365), .B1(n_336), .B2(n_364), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_429), .B(n_367), .Y(n_502) );
OAI222xp33_ASAP7_75t_L g503 ( .A1(n_395), .A2(n_375), .B1(n_384), .B2(n_382), .C1(n_347), .C2(n_349), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_414), .A2(n_383), .B1(n_365), .B2(n_356), .Y(n_504) );
OAI222xp33_ASAP7_75t_L g505 ( .A1(n_395), .A2(n_375), .B1(n_349), .B2(n_347), .C1(n_315), .C2(n_337), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_408), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_433), .A2(n_365), .B1(n_336), .B2(n_364), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_431), .A2(n_365), .B1(n_336), .B2(n_364), .Y(n_508) );
CKINVDCx11_ASAP7_75t_R g509 ( .A(n_408), .Y(n_509) );
INVx4_ASAP7_75t_SL g510 ( .A(n_408), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_395), .A2(n_349), .B1(n_347), .B2(n_307), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_463), .A2(n_365), .B1(n_364), .B2(n_336), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_443), .A2(n_340), .B1(n_365), .B2(n_343), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_494), .A2(n_364), .B1(n_336), .B2(n_360), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_440), .A2(n_364), .B1(n_336), .B2(n_360), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_468), .A2(n_360), .B1(n_349), .B2(n_347), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_470), .A2(n_360), .B1(n_349), .B2(n_347), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_499), .B(n_429), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_477), .A2(n_216), .B1(n_218), .B2(n_332), .C(n_221), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_499), .B(n_416), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_441), .A2(n_360), .B1(n_349), .B2(n_347), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_459), .A2(n_420), .B1(n_415), .B2(n_408), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_459), .A2(n_457), .B1(n_497), .B2(n_483), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_465), .B(n_415), .C(n_408), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_459), .A2(n_420), .B1(n_415), .B2(n_349), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_474), .A2(n_340), .B1(n_345), .B2(n_343), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_455), .A2(n_360), .B1(n_347), .B2(n_415), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_466), .A2(n_416), .B1(n_420), .B2(n_415), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_467), .A2(n_420), .B1(n_316), .B2(n_344), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_466), .A2(n_420), .B1(n_436), .B2(n_356), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_449), .A2(n_332), .B1(n_273), .B2(n_282), .C1(n_279), .C2(n_350), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_451), .A2(n_462), .B1(n_460), .B2(n_501), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_458), .B(n_436), .Y(n_533) );
OAI211xp5_ASAP7_75t_SL g534 ( .A1(n_488), .A2(n_224), .B(n_315), .C(n_309), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_490), .A2(n_316), .B1(n_273), .B2(n_282), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_493), .A2(n_315), .B1(n_274), .B2(n_436), .Y(n_536) );
OAI222xp33_ASAP7_75t_L g537 ( .A1(n_500), .A2(n_315), .B1(n_279), .B2(n_338), .C1(n_385), .C2(n_309), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_459), .A2(n_338), .B1(n_374), .B2(n_371), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_481), .B(n_157), .C(n_154), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_511), .A2(n_374), .B1(n_371), .B2(n_350), .Y(n_540) );
OAI222xp33_ASAP7_75t_L g541 ( .A1(n_500), .A2(n_338), .B1(n_309), .B2(n_260), .C1(n_343), .C2(n_345), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_476), .A2(n_374), .B1(n_371), .B2(n_345), .Y(n_542) );
OA21x2_ASAP7_75t_L g543 ( .A1(n_505), .A2(n_351), .B(n_334), .Y(n_543) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_476), .A2(n_374), .B1(n_371), .B2(n_354), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_452), .B(n_371), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_482), .A2(n_374), .B1(n_354), .B2(n_338), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_456), .A2(n_508), .B1(n_480), .B2(n_471), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_445), .A2(n_374), .B1(n_361), .B2(n_354), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_495), .A2(n_374), .B1(n_361), .B2(n_354), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_495), .A2(n_354), .B1(n_357), .B2(n_363), .Y(n_550) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_482), .A2(n_354), .B1(n_355), .B2(n_298), .Y(n_551) );
OAI22xp33_ASAP7_75t_L g552 ( .A1(n_453), .A2(n_363), .B1(n_353), .B2(n_357), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_446), .A2(n_286), .B1(n_297), .B2(n_298), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_450), .B(n_342), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_442), .A2(n_354), .B1(n_355), .B2(n_296), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g556 ( .A1(n_461), .A2(n_297), .B1(n_322), .B2(n_203), .C(n_153), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_485), .A2(n_353), .B1(n_278), .B2(n_355), .Y(n_557) );
NAND3xp33_ASAP7_75t_SL g558 ( .A(n_453), .B(n_297), .C(n_202), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_486), .B(n_154), .C(n_169), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_485), .A2(n_278), .B1(n_355), .B2(n_299), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_442), .A2(n_355), .B1(n_298), .B2(n_296), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_439), .B(n_348), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_464), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_504), .A2(n_278), .B1(n_299), .B2(n_320), .Y(n_564) );
AOI222xp33_ASAP7_75t_L g565 ( .A1(n_503), .A2(n_296), .B1(n_298), .B2(n_153), .C1(n_322), .C2(n_286), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_498), .A2(n_278), .B1(n_299), .B2(n_321), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_444), .B(n_348), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_496), .A2(n_278), .B1(n_299), .B2(n_321), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_447), .A2(n_286), .B1(n_299), .B2(n_321), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_442), .A2(n_358), .B1(n_348), .B2(n_286), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_479), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_502), .B(n_348), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_507), .A2(n_358), .B1(n_286), .B2(n_333), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_447), .A2(n_278), .B1(n_299), .B2(n_320), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_472), .A2(n_278), .B1(n_299), .B2(n_320), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_502), .B(n_358), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_487), .A2(n_278), .B1(n_321), .B2(n_320), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_473), .A2(n_286), .B1(n_296), .B2(n_358), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_487), .A2(n_333), .B1(n_254), .B2(n_252), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_492), .A2(n_333), .B1(n_254), .B2(n_252), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_489), .B(n_154), .C(n_157), .Y(n_581) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_509), .A2(n_333), .B(n_322), .C(n_306), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_484), .A2(n_258), .B1(n_285), .B2(n_284), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_458), .A2(n_306), .B1(n_258), .B2(n_239), .C(n_317), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_464), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_452), .B(n_154), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_469), .A2(n_287), .B1(n_284), .B2(n_285), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_491), .A2(n_331), .B1(n_292), .B2(n_325), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_448), .A2(n_331), .B1(n_293), .B2(n_325), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_469), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_509), .A2(n_331), .B1(n_293), .B2(n_325), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_475), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_478), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_478), .B(n_506), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_478), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_510), .B(n_291), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_488), .A2(n_293), .B1(n_303), .B2(n_285), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_454), .A2(n_284), .B1(n_287), .B2(n_289), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_454), .A2(n_303), .B1(n_289), .B2(n_287), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_510), .A2(n_303), .B1(n_289), .B2(n_324), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_510), .B(n_154), .Y(n_601) );
OA21x2_ASAP7_75t_L g602 ( .A1(n_510), .A2(n_317), .B(n_262), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_463), .A2(n_324), .B1(n_306), .B2(n_317), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_439), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_443), .A2(n_306), .B(n_300), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_443), .A2(n_324), .B1(n_295), .B2(n_323), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_443), .A2(n_291), .B1(n_295), .B2(n_323), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_463), .A2(n_324), .B1(n_263), .B2(n_275), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_518), .B(n_27), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_545), .B(n_154), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_513), .A2(n_275), .B(n_263), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_518), .B(n_28), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_571), .B(n_29), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_590), .B(n_154), .C(n_157), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_604), .B(n_29), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_604), .B(n_30), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_520), .B(n_30), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_520), .B(n_586), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_586), .B(n_31), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_590), .B(n_154), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_513), .A2(n_154), .B(n_157), .C(n_169), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_582), .A2(n_295), .B(n_300), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_514), .A2(n_239), .B1(n_157), .B2(n_169), .C(n_154), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_592), .B(n_32), .Y(n_624) );
NOR3xp33_ASAP7_75t_SL g625 ( .A(n_534), .B(n_33), .C(n_34), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_524), .B(n_283), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_544), .B(n_283), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_592), .B(n_33), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_565), .A2(n_324), .B1(n_157), .B2(n_169), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_594), .B(n_34), .Y(n_630) );
AOI211xp5_ASAP7_75t_SL g631 ( .A1(n_522), .A2(n_283), .B(n_330), .C(n_318), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_594), .B(n_585), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_572), .B(n_35), .Y(n_633) );
OAI221xp5_ASAP7_75t_SL g634 ( .A1(n_603), .A2(n_264), .B1(n_262), .B2(n_300), .C(n_295), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g635 ( .A1(n_571), .A2(n_528), .B(n_542), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_523), .A2(n_157), .B1(n_169), .B2(n_330), .Y(n_636) );
OAI221xp5_ASAP7_75t_SL g637 ( .A1(n_515), .A2(n_608), .B1(n_547), .B2(n_512), .C(n_517), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_593), .B(n_551), .C(n_546), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_576), .B(n_35), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_606), .A2(n_157), .B1(n_169), .B2(n_330), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_516), .B(n_36), .C(n_37), .D(n_38), .Y(n_641) );
OA21x2_ASAP7_75t_L g642 ( .A1(n_593), .A2(n_264), .B(n_323), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_554), .B(n_36), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_555), .B(n_157), .C(n_169), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_563), .B(n_157), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_561), .B(n_169), .C(n_323), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_533), .B(n_169), .C(n_323), .Y(n_647) );
AOI21xp33_ASAP7_75t_SL g648 ( .A1(n_525), .A2(n_39), .B(n_40), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_587), .A2(n_330), .B1(n_283), .B2(n_308), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_602), .B(n_169), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_526), .B(n_562), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_602), .B(n_169), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_529), .A2(n_300), .B1(n_318), .B2(n_308), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_526), .B(n_40), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_567), .B(n_41), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_595), .B(n_283), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_595), .B(n_283), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_540), .B(n_41), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_549), .B(n_295), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_558), .B(n_42), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_602), .B(n_543), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_595), .B(n_330), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_578), .A2(n_318), .B1(n_308), .B2(n_302), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_578), .A2(n_530), .B1(n_591), .B2(n_607), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_533), .B(n_330), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_543), .B(n_43), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_532), .A2(n_330), .B1(n_283), .B2(n_308), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_552), .B(n_318), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_543), .B(n_44), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_536), .B(n_308), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_598), .B(n_45), .Y(n_671) );
AOI21xp5_ASAP7_75t_SL g672 ( .A1(n_570), .A2(n_259), .B(n_300), .Y(n_672) );
AND2x2_ASAP7_75t_SL g673 ( .A(n_550), .B(n_302), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_597), .A2(n_302), .B1(n_259), .B2(n_266), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g675 ( .A1(n_553), .A2(n_302), .B1(n_259), .B2(n_267), .C(n_266), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_531), .A2(n_46), .B(n_47), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_521), .A2(n_231), .B1(n_237), .B2(n_232), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_539), .B(n_199), .C(n_206), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_589), .B(n_199), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_559), .B(n_206), .C(n_231), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_556), .A2(n_242), .B1(n_234), .B2(n_237), .C(n_232), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_527), .A2(n_234), .B1(n_242), .B2(n_270), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_564), .A2(n_270), .B1(n_267), .B2(n_281), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_583), .B(n_49), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_601), .B(n_50), .Y(n_685) );
OAI221xp5_ASAP7_75t_SL g686 ( .A1(n_569), .A2(n_52), .B1(n_53), .B2(n_54), .C(n_55), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_575), .A2(n_281), .B1(n_276), .B2(n_243), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_548), .A2(n_281), .B1(n_276), .B2(n_243), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_601), .B(n_56), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g690 ( .A1(n_581), .A2(n_276), .B(n_243), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_538), .B(n_58), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_519), .B(n_240), .C(n_63), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_569), .A2(n_240), .B1(n_66), .B2(n_67), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_599), .B(n_60), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_596), .B(n_605), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_596), .B(n_68), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_600), .B(n_69), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_584), .A2(n_71), .B1(n_72), .B2(n_75), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_535), .B(n_77), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_588), .B(n_79), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_573), .B(n_80), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_541), .A2(n_81), .B1(n_82), .B2(n_83), .C(n_84), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_580), .B(n_87), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_557), .B(n_88), .C(n_89), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_641), .B(n_537), .C(n_577), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_635), .B(n_579), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_632), .B(n_566), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_664), .A2(n_568), .B1(n_560), .B2(n_574), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_660), .B(n_90), .C(n_91), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_613), .B(n_92), .C(n_95), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_618), .B(n_96), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_648), .B(n_106), .C(n_654), .Y(n_712) );
NAND4xp75_ASAP7_75t_L g713 ( .A(n_673), .B(n_661), .C(n_695), .D(n_627), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_651), .B(n_610), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_676), .B(n_658), .C(n_615), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_637), .B(n_630), .Y(n_716) );
NAND3xp33_ASAP7_75t_L g717 ( .A(n_636), .B(n_638), .C(n_702), .Y(n_717) );
NOR3xp33_ASAP7_75t_SL g718 ( .A(n_611), .B(n_675), .C(n_686), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_661), .B(n_695), .Y(n_719) );
NOR4xp25_ASAP7_75t_SL g720 ( .A(n_627), .B(n_665), .C(n_626), .D(n_697), .Y(n_720) );
NAND3xp33_ASAP7_75t_SL g721 ( .A(n_621), .B(n_631), .C(n_666), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_609), .B(n_612), .Y(n_722) );
OA211x2_ASAP7_75t_L g723 ( .A1(n_626), .A2(n_665), .B(n_697), .C(n_656), .Y(n_723) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_672), .B(n_647), .Y(n_724) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_616), .B(n_643), .C(n_655), .Y(n_725) );
NOR2xp33_ASAP7_75t_SL g726 ( .A(n_673), .B(n_634), .Y(n_726) );
INVx4_ASAP7_75t_SL g727 ( .A(n_666), .Y(n_727) );
AO21x2_ASAP7_75t_L g728 ( .A1(n_650), .A2(n_652), .B(n_614), .Y(n_728) );
NAND3xp33_ASAP7_75t_L g729 ( .A(n_625), .B(n_669), .C(n_692), .Y(n_729) );
AND2x4_ASAP7_75t_L g730 ( .A(n_656), .B(n_662), .Y(n_730) );
NOR3xp33_ASAP7_75t_L g731 ( .A(n_617), .B(n_628), .C(n_624), .Y(n_731) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_642), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_669), .B(n_644), .C(n_657), .Y(n_733) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_633), .B(n_639), .C(n_619), .Y(n_734) );
OAI21xp5_ASAP7_75t_L g735 ( .A1(n_646), .A2(n_680), .B(n_671), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_685), .B(n_689), .Y(n_736) );
NAND4xp75_ASAP7_75t_L g737 ( .A(n_691), .B(n_701), .C(n_689), .D(n_685), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_694), .B(n_699), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_645), .B(n_696), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_699), .B(n_684), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_667), .B(n_698), .C(n_649), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g742 ( .A(n_623), .B(n_693), .C(n_700), .Y(n_742) );
AO21x2_ASAP7_75t_L g743 ( .A1(n_690), .A2(n_659), .B(n_701), .Y(n_743) );
NAND4xp75_ASAP7_75t_L g744 ( .A(n_622), .B(n_670), .C(n_668), .D(n_703), .Y(n_744) );
AO21x2_ASAP7_75t_L g745 ( .A1(n_678), .A2(n_704), .B(n_679), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_663), .B(n_653), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_682), .B(n_677), .Y(n_747) );
NAND4xp75_ASAP7_75t_L g748 ( .A(n_681), .B(n_640), .C(n_629), .D(n_688), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_674), .Y(n_749) );
AOI22x1_ASAP7_75t_L g750 ( .A1(n_683), .A2(n_453), .B1(n_476), .B2(n_466), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_687), .B(n_632), .Y(n_751) );
NAND3xp33_ASAP7_75t_SL g752 ( .A(n_635), .B(n_648), .C(n_500), .Y(n_752) );
NOR3xp33_ASAP7_75t_L g753 ( .A(n_641), .B(n_660), .C(n_613), .Y(n_753) );
NAND4xp75_ASAP7_75t_L g754 ( .A(n_613), .B(n_571), .C(n_673), .D(n_513), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_632), .B(n_618), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g756 ( .A(n_635), .B(n_660), .C(n_636), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_632), .B(n_651), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_641), .B(n_660), .C(n_613), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_632), .B(n_594), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_635), .B(n_487), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_632), .B(n_651), .Y(n_761) );
OAI211xp5_ASAP7_75t_SL g762 ( .A1(n_625), .A2(n_443), .B(n_635), .C(n_406), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_641), .A2(n_534), .B1(n_664), .B2(n_514), .Y(n_763) );
NOR3xp33_ASAP7_75t_L g764 ( .A(n_641), .B(n_660), .C(n_613), .Y(n_764) );
AO21x2_ASAP7_75t_L g765 ( .A1(n_620), .A2(n_652), .B(n_650), .Y(n_765) );
NAND4xp75_ASAP7_75t_SL g766 ( .A(n_760), .B(n_706), .C(n_716), .D(n_752), .Y(n_766) );
XOR2x2_ASAP7_75t_L g767 ( .A(n_737), .B(n_752), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_719), .B(n_759), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_732), .Y(n_769) );
INVxp67_ASAP7_75t_L g770 ( .A(n_716), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_732), .Y(n_771) );
INVx2_ASAP7_75t_SL g772 ( .A(n_765), .Y(n_772) );
XNOR2xp5_ASAP7_75t_L g773 ( .A(n_754), .B(n_750), .Y(n_773) );
XNOR2xp5_ASAP7_75t_L g774 ( .A(n_755), .B(n_714), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_762), .B(n_757), .Y(n_775) );
NAND4xp75_ASAP7_75t_SL g776 ( .A(n_740), .B(n_762), .C(n_738), .D(n_720), .Y(n_776) );
XNOR2xp5_ASAP7_75t_L g777 ( .A(n_756), .B(n_761), .Y(n_777) );
NAND4xp75_ASAP7_75t_L g778 ( .A(n_723), .B(n_724), .C(n_718), .D(n_708), .Y(n_778) );
NAND4xp75_ASAP7_75t_SL g779 ( .A(n_718), .B(n_763), .C(n_713), .D(n_727), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_727), .B(n_765), .Y(n_780) );
NAND4xp75_ASAP7_75t_L g781 ( .A(n_735), .B(n_722), .C(n_751), .D(n_711), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_753), .A2(n_764), .B1(n_758), .B2(n_726), .Y(n_782) );
NOR4xp25_ASAP7_75t_L g783 ( .A(n_763), .B(n_717), .C(n_721), .D(n_729), .Y(n_783) );
XNOR2xp5_ASAP7_75t_L g784 ( .A(n_736), .B(n_707), .Y(n_784) );
INVx3_ASAP7_75t_L g785 ( .A(n_728), .Y(n_785) );
INVx6_ASAP7_75t_L g786 ( .A(n_730), .Y(n_786) );
XNOR2xp5_ASAP7_75t_L g787 ( .A(n_753), .B(n_764), .Y(n_787) );
XOR2x2_ASAP7_75t_L g788 ( .A(n_758), .B(n_710), .Y(n_788) );
NAND4xp75_ASAP7_75t_L g789 ( .A(n_749), .B(n_739), .C(n_721), .D(n_705), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_733), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_743), .B(n_746), .Y(n_791) );
NAND4xp75_ASAP7_75t_L g792 ( .A(n_705), .B(n_743), .C(n_744), .D(n_734), .Y(n_792) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_731), .Y(n_793) );
AO22x2_ASAP7_75t_L g794 ( .A1(n_789), .A2(n_725), .B1(n_731), .B2(n_734), .Y(n_794) );
INVxp67_ASAP7_75t_L g795 ( .A(n_793), .Y(n_795) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_769), .Y(n_796) );
INVxp67_ASAP7_75t_L g797 ( .A(n_793), .Y(n_797) );
INVx1_ASAP7_75t_SL g798 ( .A(n_786), .Y(n_798) );
OA22x2_ASAP7_75t_L g799 ( .A1(n_782), .A2(n_725), .B1(n_715), .B2(n_712), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_771), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_772), .Y(n_801) );
XOR2x2_ASAP7_75t_L g802 ( .A(n_767), .B(n_709), .Y(n_802) );
XNOR2xp5_ASAP7_75t_L g803 ( .A(n_767), .B(n_715), .Y(n_803) );
XNOR2x1_ASAP7_75t_L g804 ( .A(n_787), .B(n_747), .Y(n_804) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_772), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_768), .B(n_745), .Y(n_806) );
XOR2x2_ASAP7_75t_L g807 ( .A(n_766), .B(n_748), .Y(n_807) );
XOR2x2_ASAP7_75t_L g808 ( .A(n_779), .B(n_741), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_768), .B(n_745), .Y(n_809) );
XOR2x2_ASAP7_75t_L g810 ( .A(n_787), .B(n_742), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_786), .Y(n_811) );
XOR2xp5_ASAP7_75t_L g812 ( .A(n_804), .B(n_773), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_794), .A2(n_778), .B1(n_788), .B2(n_783), .Y(n_813) );
OA22x2_ASAP7_75t_L g814 ( .A1(n_803), .A2(n_770), .B1(n_777), .B2(n_780), .Y(n_814) );
XNOR2x1_ASAP7_75t_L g815 ( .A(n_810), .B(n_788), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_807), .Y(n_816) );
XNOR2x1_ASAP7_75t_L g817 ( .A(n_807), .B(n_776), .Y(n_817) );
AOI22x1_ASAP7_75t_L g818 ( .A1(n_794), .A2(n_791), .B1(n_780), .B2(n_790), .Y(n_818) );
XNOR2x1_ASAP7_75t_L g819 ( .A(n_808), .B(n_781), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_796), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g821 ( .A(n_799), .B(n_780), .Y(n_821) );
AOI22x1_ASAP7_75t_L g822 ( .A1(n_794), .A2(n_791), .B1(n_785), .B2(n_792), .Y(n_822) );
XNOR2xp5_ASAP7_75t_L g823 ( .A(n_808), .B(n_784), .Y(n_823) );
BUFx2_ASAP7_75t_L g824 ( .A(n_794), .Y(n_824) );
XNOR2x1_ASAP7_75t_L g825 ( .A(n_802), .B(n_774), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_800), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_820), .Y(n_827) );
INVxp67_ASAP7_75t_SL g828 ( .A(n_815), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_826), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_826), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_824), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_821), .Y(n_832) );
INVxp67_ASAP7_75t_L g833 ( .A(n_812), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_821), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_828), .A2(n_813), .B1(n_814), .B2(n_799), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_833), .A2(n_814), .B1(n_799), .B2(n_803), .Y(n_836) );
AO22x2_ASAP7_75t_L g837 ( .A1(n_831), .A2(n_815), .B1(n_825), .B2(n_819), .Y(n_837) );
NAND4xp75_ASAP7_75t_L g838 ( .A(n_834), .B(n_817), .C(n_816), .D(n_822), .Y(n_838) );
INVxp67_ASAP7_75t_L g839 ( .A(n_834), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g840 ( .A1(n_836), .A2(n_816), .B1(n_802), .B2(n_810), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_837), .A2(n_818), .B1(n_832), .B2(n_804), .Y(n_841) );
NOR4xp25_ASAP7_75t_L g842 ( .A(n_839), .B(n_827), .C(n_795), .D(n_797), .Y(n_842) );
NOR4xp25_ASAP7_75t_L g843 ( .A(n_841), .B(n_838), .C(n_835), .D(n_827), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_840), .B(n_823), .Y(n_844) );
INVxp67_ASAP7_75t_SL g845 ( .A(n_844), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_843), .Y(n_846) );
AND2x4_ASAP7_75t_L g847 ( .A(n_845), .B(n_811), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_846), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_847), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_847), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_849), .Y(n_851) );
BUFx8_ASAP7_75t_L g852 ( .A(n_851), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_852), .A2(n_846), .B1(n_850), .B2(n_848), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_853), .Y(n_854) );
OAI22xp33_ASAP7_75t_L g855 ( .A1(n_854), .A2(n_842), .B1(n_798), .B2(n_829), .Y(n_855) );
OR2x2_ASAP7_75t_L g856 ( .A(n_855), .B(n_830), .Y(n_856) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_856), .A2(n_775), .B1(n_805), .B2(n_801), .C(n_809), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_857), .A2(n_775), .B1(n_806), .B2(n_809), .Y(n_858) );
endmodule