module fake_jpeg_32122_n_106 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_36),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_59),
.Y(n_60)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_37),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_31),
.Y(n_69)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_51),
.A3(n_32),
.B1(n_40),
.B2(n_11),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_6),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_71),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_7),
.C(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_12),
.Y(n_82)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_15),
.Y(n_93)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_80),
.B1(n_60),
.B2(n_16),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_80),
.Y(n_95)
);

NOR2xp67_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_13),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_89),
.B(n_93),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_90),
.C(n_91),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_92),
.C(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_94),
.C(n_86),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_102),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_88),
.B(n_22),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_19),
.B(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_24),
.Y(n_106)
);


endmodule