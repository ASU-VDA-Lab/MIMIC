module fake_jpeg_17674_n_123 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_123);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_31),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_0),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_6),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_37),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_7),
.B1(n_24),
.B2(n_17),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_23),
.B1(n_30),
.B2(n_36),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_7),
.C(n_24),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_18),
.B(n_26),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_20),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_42),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

OA21x2_ASAP7_75t_L g62 ( 
.A1(n_29),
.A2(n_23),
.B(n_20),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_28),
.A2(n_23),
.B1(n_26),
.B2(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_37),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_34),
.A2(n_18),
.B(n_28),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_59),
.B(n_61),
.Y(n_75)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_54),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_81),
.C(n_62),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_62),
.B1(n_55),
.B2(n_47),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_85),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_75),
.C(n_73),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_96),
.B1(n_70),
.B2(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_52),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_89),
.C(n_93),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_79),
.B(n_81),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_79),
.B1(n_69),
.B2(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_111),
.B(n_112),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_99),
.C(n_100),
.Y(n_113)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_109),
.B(n_101),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_108),
.A2(n_101),
.B(n_102),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_107),
.C(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_117),
.B(n_118),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_115),
.C(n_120),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_122),
.B(n_83),
.Y(n_123)
);


endmodule