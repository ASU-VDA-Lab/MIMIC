module fake_jpeg_31552_n_386 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_57),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_67),
.Y(n_99)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_30),
.Y(n_91)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_15),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_69),
.A2(n_22),
.B1(n_39),
.B2(n_23),
.Y(n_119)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_33),
.B(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_76),
.Y(n_113)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_74),
.Y(n_109)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_20),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_37),
.B(n_14),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_79),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_20),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_25),
.B1(n_29),
.B2(n_41),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_84),
.A2(n_97),
.B1(n_119),
.B2(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_104),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_23),
.B1(n_19),
.B2(n_38),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_94),
.A2(n_103),
.B1(n_115),
.B2(n_122),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_96),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_43),
.B1(n_19),
.B2(n_38),
.Y(n_97)
);

BUFx16f_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_118),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_30),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_23),
.B1(n_34),
.B2(n_40),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_45),
.B(n_29),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_28),
.B1(n_41),
.B2(n_40),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_45),
.B(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_121),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_58),
.A2(n_23),
.B1(n_22),
.B2(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_42),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_60),
.B(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_50),
.B(n_14),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_39),
.B1(n_13),
.B2(n_12),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_65),
.A2(n_39),
.B1(n_13),
.B2(n_4),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_51),
.B(n_0),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_52),
.B1(n_66),
.B2(n_73),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_130),
.A2(n_133),
.B1(n_145),
.B2(n_150),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_75),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_131),
.B(n_163),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_74),
.B1(n_70),
.B2(n_72),
.Y(n_133)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_136),
.B(n_156),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_141),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_158),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_68),
.C(n_79),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_171),
.C(n_88),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_39),
.B1(n_1),
.B2(n_4),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_148),
.A2(n_152),
.B(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_155),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_95),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_101),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_5),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_8),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_86),
.B(n_9),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_125),
.B(n_9),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_9),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_106),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_106),
.A2(n_111),
.B1(n_95),
.B2(n_93),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_168),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_83),
.A2(n_10),
.B1(n_108),
.B2(n_93),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_169),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_82),
.B(n_10),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_96),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_109),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_83),
.B(n_108),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_106),
.A2(n_111),
.B1(n_102),
.B2(n_88),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_111),
.B(n_117),
.C(n_116),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_112),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_92),
.C(n_102),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_124),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_176),
.B(n_178),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_140),
.B(n_90),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_90),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_179),
.B(n_183),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_131),
.B(n_112),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_109),
.B(n_81),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_159),
.B(n_157),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_132),
.A2(n_129),
.B(n_87),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_187),
.A2(n_212),
.B(n_161),
.Y(n_248)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_81),
.C(n_87),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_156),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_134),
.B(n_109),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_192),
.B(n_202),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_195),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_92),
.C(n_128),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_167),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_201),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_134),
.B(n_128),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_213),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_147),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_117),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_SL g208 ( 
.A(n_162),
.B(n_116),
.C(n_146),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_208),
.B(n_141),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_155),
.A2(n_132),
.B(n_139),
.C(n_170),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_156),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_164),
.B(n_147),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_173),
.B1(n_145),
.B2(n_139),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_217),
.A2(n_219),
.B1(n_223),
.B2(n_247),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_243),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_133),
.B1(n_130),
.B2(n_143),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_222),
.A2(n_248),
.B(n_185),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_192),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_225),
.B(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_137),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_177),
.C(n_193),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_187),
.B(n_205),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_205),
.B1(n_178),
.B2(n_183),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_233),
.A2(n_246),
.B1(n_191),
.B2(n_211),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_163),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_238),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_137),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_236),
.B(n_244),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_175),
.B(n_146),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_168),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_177),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_174),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_184),
.B(n_169),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_181),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_205),
.A2(n_172),
.B1(n_153),
.B2(n_149),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_190),
.A2(n_152),
.B1(n_160),
.B2(n_135),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_249),
.B(n_251),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_260),
.B(n_276),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_214),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_264),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_211),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_270),
.C(n_275),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_195),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_231),
.A2(n_197),
.B(n_212),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_226),
.B(n_217),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_233),
.A2(n_190),
.B1(n_204),
.B2(n_179),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_274),
.B1(n_224),
.B2(n_221),
.Y(n_279)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_268),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_215),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_223),
.A2(n_185),
.B1(n_208),
.B2(n_204),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_226),
.B1(n_220),
.B2(n_245),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_224),
.B(n_189),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_273),
.B(n_237),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_215),
.B(n_230),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_189),
.B(n_181),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_182),
.C(n_194),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_229),
.C(n_244),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_138),
.C(n_199),
.Y(n_278)
);

NOR3xp33_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_220),
.C(n_243),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_279),
.B(n_298),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_281),
.B(n_282),
.C(n_284),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_285),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_234),
.C(n_240),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_266),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_290),
.Y(n_303)
);

XOR2x2_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_237),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_271),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_294),
.B1(n_250),
.B2(n_261),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_SL g289 ( 
.A(n_258),
.B(n_238),
.C(n_241),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_SL g306 ( 
.A(n_289),
.B(n_255),
.C(n_262),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_293),
.A2(n_257),
.B(n_254),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_261),
.A2(n_246),
.B1(n_219),
.B2(n_235),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_269),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_296),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_302),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_253),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_273),
.B(n_255),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_239),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_247),
.B1(n_227),
.B2(n_232),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_263),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_304),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_300),
.C(n_282),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_272),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_307),
.A2(n_321),
.B(n_286),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_276),
.B(n_262),
.C(n_264),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_308),
.B(n_316),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_285),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_317),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_249),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_318),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_289),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_296),
.B(n_277),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_291),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_287),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_252),
.C(n_259),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_291),
.C(n_284),
.Y(n_326)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_303),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_325),
.B(n_328),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_334),
.C(n_335),
.Y(n_345)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_309),
.B(n_303),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_314),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_312),
.B(n_301),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_299),
.C(n_279),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_299),
.C(n_293),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_294),
.C(n_302),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_338),
.C(n_335),
.Y(n_348)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_315),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_288),
.C(n_301),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_349),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_SL g341 ( 
.A1(n_339),
.A2(n_304),
.B(n_307),
.C(n_305),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_352),
.B(n_292),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_334),
.B(n_315),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_343),
.B(n_346),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g359 ( 
.A1(n_344),
.A2(n_292),
.B(n_268),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_333),
.B(n_306),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_348),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_304),
.C(n_307),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_332),
.A2(n_313),
.B(n_305),
.Y(n_350)
);

OAI221xp5_ASAP7_75t_L g353 ( 
.A1(n_350),
.A2(n_323),
.B1(n_331),
.B2(n_308),
.C(n_339),
.Y(n_353)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

FAx1_ASAP7_75t_SL g354 ( 
.A(n_349),
.B(n_319),
.CI(n_330),
.CON(n_354),
.SN(n_354)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_357),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_351),
.B(n_336),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_326),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_358),
.A2(n_362),
.B1(n_363),
.B2(n_142),
.Y(n_366)
);

AOI21x1_ASAP7_75t_L g371 ( 
.A1(n_359),
.A2(n_154),
.B(n_362),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_360),
.A2(n_186),
.B(n_209),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_341),
.A2(n_292),
.B1(n_329),
.B2(n_199),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_341),
.A2(n_348),
.B1(n_345),
.B2(n_329),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_361),
.A2(n_341),
.B1(n_345),
.B2(n_194),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_364),
.B(n_366),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_360),
.A2(n_209),
.B1(n_186),
.B2(n_161),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_355),
.A2(n_154),
.B(n_135),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g374 ( 
.A1(n_370),
.A2(n_354),
.B(n_356),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_371),
.A2(n_372),
.B(n_367),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_363),
.C(n_354),
.Y(n_372)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_376),
.Y(n_379)
);

AOI21x1_ASAP7_75t_L g376 ( 
.A1(n_365),
.A2(n_369),
.B(n_370),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_377),
.B(n_372),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_382),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_368),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_381),
.A2(n_378),
.B(n_379),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_383),
.B(n_379),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_384),
.Y(n_386)
);


endmodule