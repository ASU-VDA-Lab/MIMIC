module fake_aes_11019_n_671 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_671);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_671;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_40), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_47), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_10), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_81), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_70), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_25), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_4), .Y(n_91) );
BUFx3_ASAP7_75t_L g92 ( .A(n_0), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_27), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_2), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_66), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_71), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_19), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_32), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_68), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_26), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_44), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_17), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_65), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_62), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_43), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_50), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_83), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_67), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_56), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_72), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_22), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_37), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_84), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_21), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_63), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_12), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_60), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_10), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_14), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_61), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_9), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_31), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_91), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_99), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_120), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_86), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_99), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_92), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_92), .B(n_1), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_90), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_113), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
OAI21x1_ASAP7_75t_L g138 ( .A1(n_89), .A2(n_39), .B(n_80), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_113), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_123), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_123), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_93), .A2(n_38), .B(n_79), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_95), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_95), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_117), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_97), .B(n_5), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_98), .Y(n_150) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_98), .A2(n_41), .B(n_78), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_91), .B(n_6), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_94), .B(n_7), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_100), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_130), .B(n_85), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_145), .B(n_94), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_132), .Y(n_158) );
XOR2xp5_ASAP7_75t_L g159 ( .A(n_148), .B(n_96), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_129), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_144), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_129), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_125), .B(n_102), .Y(n_164) );
INVx8_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_129), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
BUFx10_ASAP7_75t_L g168 ( .A(n_132), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_148), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_125), .B(n_121), .Y(n_171) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_152), .B(n_100), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_127), .A2(n_119), .B1(n_102), .B2(n_104), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_128), .B(n_85), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_128), .B(n_106), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_133), .B(n_106), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_133), .B(n_115), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_137), .B(n_110), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_137), .B(n_119), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_126), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_152), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_142), .B(n_104), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_142), .B(n_115), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_146), .B(n_109), .Y(n_187) );
BUFx8_ASAP7_75t_SL g188 ( .A(n_152), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_153), .A2(n_87), .B1(n_122), .B2(n_101), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_146), .B(n_108), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_182), .B(n_153), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_158), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_177), .B(n_154), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_173), .A2(n_153), .B1(n_154), .B2(n_147), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_173), .A2(n_153), .B1(n_149), .B2(n_127), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_186), .B(n_147), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_171), .B(n_147), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_182), .B(n_124), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_156), .B(n_147), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_158), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_158), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_173), .A2(n_124), .B1(n_150), .B2(n_144), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g206 ( .A1(n_170), .A2(n_126), .B1(n_138), .B2(n_143), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_175), .B(n_126), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_169), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_164), .B(n_126), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_165), .A2(n_150), .B1(n_140), .B2(n_131), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_174), .A2(n_131), .B(n_134), .C(n_136), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_176), .B(n_107), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_188), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_169), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_164), .B(n_131), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_184), .B(n_114), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_184), .B(n_111), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_180), .B(n_140), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_180), .B(n_134), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_169), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_185), .B(n_134), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_185), .B(n_141), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
NAND2xp33_ASAP7_75t_L g228 ( .A(n_165), .B(n_150), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_178), .B(n_136), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_172), .B(n_151), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_165), .B(n_136), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_172), .A2(n_150), .B1(n_141), .B2(n_140), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_184), .B(n_105), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_157), .B(n_141), .Y(n_234) );
INVxp67_ASAP7_75t_L g235 ( .A(n_157), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_172), .B(n_103), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_189), .B(n_101), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g238 ( .A(n_168), .B(n_118), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_179), .B(n_118), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_168), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_168), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_192), .A2(n_150), .B1(n_112), .B2(n_116), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_235), .A2(n_187), .B(n_181), .C(n_191), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_197), .B(n_168), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_194), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_215), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_221), .B(n_159), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_217), .Y(n_248) );
CKINVDCx14_ASAP7_75t_R g249 ( .A(n_198), .Y(n_249) );
BUFx2_ASAP7_75t_SL g250 ( .A(n_196), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_201), .B(n_159), .Y(n_252) );
NAND2x1p5_ASAP7_75t_L g253 ( .A(n_196), .B(n_150), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_208), .A2(n_143), .B(n_151), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_208), .A2(n_191), .B(n_155), .Y(n_257) );
O2A1O1Ixp5_ASAP7_75t_L g258 ( .A1(n_193), .A2(n_160), .B(n_163), .C(n_190), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_225), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_195), .A2(n_129), .B1(n_135), .B2(n_139), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_196), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_210), .A2(n_181), .B(n_151), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_238), .A2(n_135), .B1(n_139), .B2(n_143), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_221), .B(n_7), .Y(n_264) );
OR2x6_ASAP7_75t_SL g265 ( .A(n_237), .B(n_8), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_194), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_212), .A2(n_161), .B(n_183), .C(n_155), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_225), .B(n_8), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g269 ( .A1(n_236), .A2(n_135), .B1(n_139), .B2(n_143), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_234), .B(n_9), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_209), .A2(n_161), .B(n_183), .C(n_162), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_226), .B(n_151), .Y(n_272) );
AOI21xp33_ASAP7_75t_L g273 ( .A1(n_228), .A2(n_205), .B(n_207), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_226), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_203), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_203), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_222), .Y(n_277) );
NOR2xp67_ASAP7_75t_L g278 ( .A(n_242), .B(n_11), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_222), .B(n_135), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_222), .B(n_11), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_210), .A2(n_162), .B(n_167), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_200), .B(n_139), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_231), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_214), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_214), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_204), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_239), .A2(n_199), .B(n_219), .C(n_220), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_240), .B(n_139), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_242), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_213), .B(n_12), .Y(n_290) );
AOI21xp33_ASAP7_75t_L g291 ( .A1(n_228), .A2(n_139), .B(n_135), .Y(n_291) );
AO32x2_ASAP7_75t_L g292 ( .A1(n_260), .A2(n_206), .A3(n_230), .B1(n_135), .B2(n_232), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_254), .Y(n_293) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_272), .A2(n_218), .B(n_204), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_272), .A2(n_218), .B(n_240), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_248), .B(n_202), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_289), .A2(n_229), .B1(n_211), .B2(n_241), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_270), .A2(n_241), .B(n_233), .C(n_216), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_245), .Y(n_300) );
BUFx8_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_268), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_256), .B(n_230), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_266), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_249), .B(n_224), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_259), .A2(n_230), .B1(n_224), .B2(n_216), .Y(n_306) );
OAI22x1_ASAP7_75t_L g307 ( .A1(n_264), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_276), .Y(n_308) );
O2A1O1Ixp5_ASAP7_75t_SL g309 ( .A1(n_260), .A2(n_291), .B(n_282), .C(n_279), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_274), .B(n_227), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_247), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_SL g312 ( .A1(n_267), .A2(n_167), .B(n_166), .C(n_190), .Y(n_312) );
AO32x2_ASAP7_75t_L g313 ( .A1(n_269), .A2(n_167), .A3(n_166), .B1(n_163), .B2(n_17), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_275), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_254), .Y(n_315) );
NOR2xp67_ASAP7_75t_R g316 ( .A(n_254), .B(n_227), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_286), .Y(n_317) );
OAI22xp33_ASAP7_75t_L g318 ( .A1(n_265), .A2(n_166), .B1(n_15), .B2(n_16), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_255), .A2(n_49), .B(n_77), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_262), .A2(n_48), .B(n_76), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_247), .B(n_13), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_246), .Y(n_322) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_290), .B(n_16), .C(n_18), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_277), .A2(n_20), .B1(n_23), .B2(n_24), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_252), .A2(n_28), .B1(n_29), .B2(n_30), .C(n_33), .Y(n_325) );
CKINVDCx6p67_ASAP7_75t_R g326 ( .A(n_247), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_282), .A2(n_34), .B(n_35), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_317), .Y(n_328) );
AO21x2_ASAP7_75t_L g329 ( .A1(n_312), .A2(n_263), .B(n_278), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_314), .B(n_244), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_315), .B(n_251), .Y(n_331) );
AO21x2_ASAP7_75t_L g332 ( .A1(n_312), .A2(n_291), .B(n_288), .Y(n_332) );
OA21x2_ASAP7_75t_L g333 ( .A1(n_320), .A2(n_258), .B(n_288), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_315), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_302), .A2(n_287), .B(n_243), .C(n_244), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_318), .A2(n_283), .B1(n_250), .B2(n_261), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_301), .Y(n_338) );
OA21x2_ASAP7_75t_L g339 ( .A1(n_299), .A2(n_273), .B(n_281), .Y(n_339) );
CKINVDCx8_ASAP7_75t_R g340 ( .A(n_315), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_296), .B(n_253), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_298), .B(n_273), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_308), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_294), .B(n_271), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_303), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_310), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_311), .A2(n_253), .B1(n_257), .B2(n_284), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_301), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_295), .B(n_285), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_299), .A2(n_319), .B(n_327), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_306), .A2(n_257), .B(n_285), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_293), .B(n_285), .Y(n_354) );
OA21x2_ASAP7_75t_L g355 ( .A1(n_327), .A2(n_284), .B(n_42), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_347), .B(n_321), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_337), .A2(n_318), .B1(n_326), .B2(n_305), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_337), .A2(n_305), .B1(n_307), .B2(n_325), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_334), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_328), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_347), .B(n_293), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_346), .Y(n_363) );
AO21x2_ASAP7_75t_L g364 ( .A1(n_352), .A2(n_323), .B(n_292), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_334), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_343), .B(n_297), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_346), .B(n_306), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_335), .B(n_292), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_335), .B(n_292), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_341), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_352), .A2(n_325), .B(n_292), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g374 ( .A1(n_336), .A2(n_324), .B1(n_309), .B2(n_284), .C(n_313), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_334), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_334), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_343), .B(n_322), .C(n_316), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_353), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_341), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_344), .B(n_313), .Y(n_381) );
OA211x2_ASAP7_75t_L g382 ( .A1(n_348), .A2(n_313), .B(n_45), .C(n_46), .Y(n_382) );
NAND2x1_ASAP7_75t_L g383 ( .A(n_355), .B(n_313), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_379), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_376), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_356), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_356), .B(n_344), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_361), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_361), .B(n_330), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_367), .B(n_330), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_369), .B(n_339), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_376), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_370), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_369), .B(n_353), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_363), .B(n_345), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_371), .B(n_353), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_372), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_371), .B(n_339), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_357), .B(n_345), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_381), .B(n_339), .Y(n_400) );
BUFx12f_ASAP7_75t_L g401 ( .A(n_357), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_379), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_379), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_377), .Y(n_405) );
INVxp67_ASAP7_75t_SL g406 ( .A(n_383), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_365), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_380), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_363), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_368), .B(n_342), .Y(n_411) );
AO22x1_ASAP7_75t_L g412 ( .A1(n_358), .A2(n_349), .B1(n_338), .B2(n_331), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_370), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_359), .A2(n_342), .B1(n_338), .B2(n_349), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_368), .B(n_350), .Y(n_415) );
OA21x2_ASAP7_75t_L g416 ( .A1(n_374), .A2(n_350), .B(n_351), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_378), .A2(n_331), .B1(n_354), .B2(n_329), .C(n_332), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_381), .Y(n_418) );
AO21x2_ASAP7_75t_L g419 ( .A1(n_364), .A2(n_332), .B(n_329), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_362), .B(n_331), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_365), .B(n_354), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_365), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_386), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_418), .B(n_364), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_418), .B(n_364), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_385), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_401), .A2(n_382), .B1(n_370), .B2(n_373), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_384), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_400), .B(n_373), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_385), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_400), .B(n_373), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_392), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_415), .B(n_362), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_400), .B(n_373), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_410), .B(n_377), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_410), .B(n_383), .Y(n_439) );
BUFx2_ASAP7_75t_L g440 ( .A(n_392), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_415), .B(n_375), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_401), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_386), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_391), .B(n_375), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_395), .B(n_375), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_404), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_388), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_388), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_391), .B(n_366), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_403), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_391), .B(n_366), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_398), .B(n_366), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_398), .B(n_360), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_360), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_421), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_401), .B(n_340), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_403), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_394), .B(n_360), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_397), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_404), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_397), .Y(n_461) );
INVx6_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_394), .B(n_360), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_411), .B(n_339), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_387), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_407), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_396), .B(n_360), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_396), .B(n_360), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_402), .B(n_339), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_402), .B(n_351), .Y(n_470) );
OR2x6_ASAP7_75t_L g471 ( .A(n_412), .B(n_355), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_407), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_408), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_408), .B(n_351), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_393), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_411), .B(n_399), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_405), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_423), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_431), .B(n_433), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_465), .B(n_399), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_476), .B(n_387), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_443), .Y(n_483) );
INVxp33_ASAP7_75t_L g484 ( .A(n_460), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_466), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_476), .B(n_409), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_443), .B(n_409), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_431), .B(n_416), .Y(n_488) );
OR2x6_ASAP7_75t_L g489 ( .A(n_471), .B(n_412), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_446), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_447), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_435), .B(n_420), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_447), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_448), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_466), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_433), .B(n_416), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_448), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_436), .B(n_453), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_459), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_444), .B(n_405), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_466), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_436), .B(n_416), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_459), .B(n_395), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_461), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_435), .B(n_420), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_461), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_446), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_453), .B(n_416), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_473), .Y(n_509) );
BUFx2_ASAP7_75t_L g510 ( .A(n_442), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_416), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_441), .B(n_405), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_473), .B(n_390), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_438), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_454), .B(n_406), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_442), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_472), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_438), .Y(n_518) );
OR2x6_ASAP7_75t_L g519 ( .A(n_471), .B(n_393), .Y(n_519) );
INVx3_ASAP7_75t_SL g520 ( .A(n_456), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_444), .B(n_390), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_441), .B(n_389), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_428), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_445), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_445), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_449), .B(n_406), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_449), .B(n_389), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_451), .B(n_422), .Y(n_528) );
OR4x1_ASAP7_75t_L g529 ( .A(n_471), .B(n_382), .C(n_414), .D(n_413), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_451), .B(n_422), .Y(n_530) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_471), .B(n_393), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_452), .B(n_407), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_455), .B(n_413), .Y(n_533) );
NAND2x1_ASAP7_75t_L g534 ( .A(n_428), .B(n_421), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_452), .B(n_422), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_458), .B(n_419), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_424), .B(n_413), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_434), .B(n_417), .C(n_429), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_524), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_525), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
NOR2x1_ASAP7_75t_L g542 ( .A(n_510), .B(n_471), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_521), .B(n_479), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_516), .B(n_486), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_514), .B(n_424), .Y(n_545) );
INVxp67_ASAP7_75t_L g546 ( .A(n_523), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_522), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_518), .B(n_426), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_479), .B(n_440), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_478), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_498), .B(n_462), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_489), .A2(n_475), .B(n_417), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_498), .B(n_462), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_490), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_488), .B(n_426), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_527), .B(n_440), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_538), .B(n_477), .C(n_439), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_481), .B(n_432), .Y(n_558) );
INVxp33_ASAP7_75t_L g559 ( .A(n_512), .Y(n_559) );
AO22x1_ASAP7_75t_L g560 ( .A1(n_531), .A2(n_475), .B1(n_432), .B2(n_439), .Y(n_560) );
OAI21xp33_ASAP7_75t_L g561 ( .A1(n_484), .A2(n_469), .B(n_464), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_500), .B(n_462), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_480), .B(n_464), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_520), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_492), .B(n_463), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_482), .Y(n_566) );
NAND2x1_ASAP7_75t_SL g567 ( .A(n_520), .B(n_474), .Y(n_567) );
INVxp67_ASAP7_75t_SL g568 ( .A(n_507), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_515), .B(n_462), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_488), .B(n_469), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_505), .B(n_458), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_496), .B(n_470), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_515), .B(n_462), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_496), .B(n_474), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_526), .B(n_455), .Y(n_575) );
NOR2xp67_ASAP7_75t_SL g576 ( .A(n_523), .B(n_340), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_526), .B(n_455), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_528), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_489), .A2(n_437), .B1(n_425), .B2(n_427), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_507), .Y(n_580) );
OAI32xp33_ASAP7_75t_L g581 ( .A1(n_484), .A2(n_430), .A3(n_425), .B1(n_427), .B2(n_437), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_489), .A2(n_519), .B1(n_534), .B2(n_537), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_483), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_530), .B(n_463), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_491), .Y(n_585) );
AOI211x1_ASAP7_75t_L g586 ( .A1(n_502), .A2(n_470), .B(n_467), .C(n_468), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_485), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_493), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_539), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_540), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_564), .Y(n_591) );
OAI31xp33_ASAP7_75t_L g592 ( .A1(n_582), .A2(n_502), .A3(n_508), .B(n_511), .Y(n_592) );
INVxp33_ASAP7_75t_L g593 ( .A(n_567), .Y(n_593) );
AOI32xp33_ASAP7_75t_L g594 ( .A1(n_582), .A2(n_511), .A3(n_508), .B1(n_536), .B2(n_535), .Y(n_594) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_561), .A2(n_536), .B(n_519), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_550), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_544), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_551), .B(n_519), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_547), .B(n_535), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_586), .A2(n_513), .B1(n_529), .B2(n_503), .C(n_494), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_580), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_559), .B(n_509), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_566), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_548), .B(n_528), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_583), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_585), .Y(n_606) );
INVxp67_ASAP7_75t_L g607 ( .A(n_541), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_578), .B(n_532), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_588), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_556), .Y(n_610) );
AOI221xp5_ASAP7_75t_SL g611 ( .A1(n_552), .A2(n_497), .B1(n_506), .B2(n_504), .C(n_499), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_548), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g613 ( .A(n_576), .B(n_533), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_553), .B(n_533), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_587), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_552), .A2(n_487), .B1(n_529), .B2(n_455), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_546), .A2(n_517), .B(n_501), .C(n_495), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_569), .B(n_533), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_549), .A2(n_455), .B1(n_501), .B2(n_495), .Y(n_619) );
NOR2x1_ASAP7_75t_L g620 ( .A(n_557), .B(n_517), .Y(n_620) );
BUFx3_ASAP7_75t_L g621 ( .A(n_554), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_592), .A2(n_579), .B1(n_542), .B2(n_546), .C(n_568), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_616), .B(n_579), .Y(n_623) );
O2A1O1Ixp5_ASAP7_75t_L g624 ( .A1(n_616), .A2(n_560), .B(n_568), .C(n_581), .Y(n_624) );
AOI211xp5_ASAP7_75t_SL g625 ( .A1(n_591), .A2(n_558), .B(n_543), .C(n_574), .Y(n_625) );
NOR2xp67_ASAP7_75t_L g626 ( .A(n_595), .B(n_572), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_594), .A2(n_600), .B1(n_611), .B2(n_597), .C(n_602), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_598), .B(n_614), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_593), .A2(n_572), .B(n_574), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_620), .A2(n_555), .B(n_570), .C(n_545), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_612), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_602), .A2(n_555), .B1(n_545), .B2(n_570), .C(n_563), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_610), .A2(n_573), .B1(n_562), .B2(n_575), .C(n_577), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_593), .A2(n_584), .B1(n_571), .B2(n_565), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_618), .B(n_455), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_596), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_617), .A2(n_485), .B(n_425), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_613), .A2(n_450), .B1(n_457), .B2(n_427), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_589), .B(n_468), .Y(n_639) );
NAND4xp25_ASAP7_75t_L g640 ( .A(n_621), .B(n_467), .C(n_421), .D(n_472), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_613), .A2(n_472), .B1(n_457), .B2(n_450), .C(n_437), .Y(n_641) );
NAND4xp75_ASAP7_75t_L g642 ( .A(n_624), .B(n_599), .C(n_608), .D(n_590), .Y(n_642) );
OA211x2_ASAP7_75t_L g643 ( .A1(n_627), .A2(n_607), .B(n_604), .C(n_619), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_625), .A2(n_621), .B(n_608), .C(n_609), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_622), .A2(n_619), .B1(n_603), .B2(n_606), .C(n_605), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_623), .A2(n_601), .B(n_615), .C(n_355), .Y(n_646) );
OAI211xp5_ASAP7_75t_SL g647 ( .A1(n_625), .A2(n_601), .B(n_615), .C(n_457), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_626), .A2(n_419), .B1(n_430), .B2(n_450), .Y(n_648) );
AOI31xp33_ASAP7_75t_L g649 ( .A1(n_638), .A2(n_331), .A3(n_430), .B(n_354), .Y(n_649) );
OAI21xp33_ASAP7_75t_L g650 ( .A1(n_629), .A2(n_354), .B(n_419), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_630), .A2(n_419), .B1(n_329), .B2(n_332), .C(n_355), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_640), .A2(n_355), .B(n_351), .C(n_329), .Y(n_652) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_644), .A2(n_632), .B1(n_634), .B2(n_641), .C(n_633), .Y(n_653) );
NAND4xp25_ASAP7_75t_SL g654 ( .A(n_645), .B(n_628), .C(n_639), .D(n_631), .Y(n_654) );
NAND4xp25_ASAP7_75t_SL g655 ( .A(n_646), .B(n_643), .C(n_648), .D(n_642), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_651), .B(n_636), .C(n_637), .D(n_635), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_647), .A2(n_351), .B(n_332), .C(n_333), .Y(n_657) );
NAND4xp25_ASAP7_75t_SL g658 ( .A(n_652), .B(n_36), .C(n_51), .D(n_52), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_656), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_657), .B(n_650), .Y(n_660) );
NOR3xp33_ASAP7_75t_SL g661 ( .A(n_655), .B(n_649), .C(n_54), .Y(n_661) );
INVxp33_ASAP7_75t_SL g662 ( .A(n_654), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_660), .Y(n_663) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_662), .Y(n_664) );
OAI22xp5_ASAP7_75t_SL g665 ( .A1(n_664), .A2(n_662), .B1(n_659), .B2(n_661), .Y(n_665) );
OAI22xp5_ASAP7_75t_SL g666 ( .A1(n_663), .A2(n_653), .B1(n_658), .B2(n_333), .Y(n_666) );
AOI22x1_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_53), .B1(n_55), .B2(n_57), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_667), .A2(n_665), .B1(n_333), .B2(n_64), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_58), .B1(n_59), .B2(n_69), .C(n_73), .Y(n_669) );
AO21x2_ASAP7_75t_L g670 ( .A1(n_669), .A2(n_74), .B(n_75), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_82), .B1(n_333), .B2(n_662), .Y(n_671) );
endmodule