module fake_jpeg_21107_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_6),
.B(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_18),
.A2(n_17),
.B1(n_13),
.B2(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_12),
.B(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_1),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_26),
.Y(n_45)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_24),
.B1(n_17),
.B2(n_13),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_39),
.B1(n_42),
.B2(n_41),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_24),
.B1(n_13),
.B2(n_16),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_26),
.C(n_19),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_19),
.C(n_20),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_26),
.B1(n_20),
.B2(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_15),
.B1(n_14),
.B2(n_10),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_30),
.B1(n_28),
.B2(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_36),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_25),
.C(n_11),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_46),
.B(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_60),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_54),
.B1(n_47),
.B2(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_51),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_56),
.C(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_66),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_43),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_2),
.B(n_4),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_6),
.C(n_7),
.Y(n_71)
);

NOR2xp67_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_65),
.Y(n_70)
);

AOI31xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.A3(n_7),
.B(n_9),
.Y(n_72)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_72),
.Y(n_73)
);


endmodule