module fake_netlist_5_1655_n_973 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_973);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_973;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_523;
wire n_268;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_640;
wire n_275;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_947;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_448;
wire n_259;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_579;
wire n_250;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_964;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_795;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_432;
wire n_553;
wire n_727;
wire n_395;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_328;
wire n_214;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_928;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_477;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_891;
wire n_466;
wire n_239;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_966;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_679;
wire n_425;
wire n_513;
wire n_237;
wire n_647;
wire n_527;
wire n_707;
wire n_407;
wire n_710;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_404;
wire n_233;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_960;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_80),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_103),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_3),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_65),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_106),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_46),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_167),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_101),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_66),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_177),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_186),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_96),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_56),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_71),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_133),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_182),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_78),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_99),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_55),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_27),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_4),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_150),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_51),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_113),
.Y(n_231)
);

BUFx2_ASAP7_75t_SL g232 ( 
.A(n_180),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_87),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_84),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_154),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_155),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_193),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_173),
.Y(n_239)
);

BUFx8_ASAP7_75t_SL g240 ( 
.A(n_164),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_21),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_57),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_49),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_44),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_23),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_104),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_142),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_21),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_157),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_132),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_123),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_199),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_9),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_172),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_110),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_61),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_36),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_159),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_69),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_174),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_13),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_22),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_12),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_168),
.Y(n_264)
);

BUFx2_ASAP7_75t_SL g265 ( 
.A(n_93),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_83),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_75),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_187),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_72),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_112),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_102),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_25),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_45),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_1),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_124),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_163),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_74),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_81),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_120),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_86),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_3),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_26),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_131),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_13),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_39),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_198),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_116),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_176),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_140),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_92),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_128),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_107),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_183),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_178),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_60),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_184),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_196),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_98),
.Y(n_301)
);

BUFx2_ASAP7_75t_SL g302 ( 
.A(n_197),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_50),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_137),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_138),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_5),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_31),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_166),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_158),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_204),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_208),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_200),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_201),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_248),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_235),
.B(n_0),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_235),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_228),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_243),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_206),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_208),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_253),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_202),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_217),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_219),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_208),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_223),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_227),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_247),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_264),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_203),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_235),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_243),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_205),
.Y(n_346)
);

BUFx2_ASAP7_75t_SL g347 ( 
.A(n_212),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_208),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_294),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_261),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_240),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_207),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_209),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_262),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_240),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_218),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_263),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_274),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_218),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_222),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_222),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_244),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_242),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_242),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_244),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_244),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_244),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_255),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_221),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_210),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_211),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_276),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_252),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_252),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_230),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_230),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_318),
.B(n_230),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_373),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

BUFx8_ASAP7_75t_L g391 ( 
.A(n_383),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_380),
.B(n_290),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_381),
.B(n_289),
.Y(n_394)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_375),
.A2(n_293),
.B1(n_224),
.B2(n_225),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_315),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_316),
.B(n_330),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_319),
.B(n_214),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_329),
.A2(n_365),
.B1(n_322),
.B2(n_352),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_339),
.B(n_346),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_215),
.Y(n_409)
);

BUFx8_ASAP7_75t_L g410 ( 
.A(n_379),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_347),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_355),
.Y(n_414)
);

OA21x2_ASAP7_75t_L g415 ( 
.A1(n_366),
.A2(n_220),
.B(n_216),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_367),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_310),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

AND2x2_ASAP7_75t_SL g419 ( 
.A(n_323),
.B(n_382),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_324),
.A2(n_265),
.B(n_232),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_311),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_341),
.B(n_226),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_321),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_312),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_359),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_327),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_314),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_332),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_334),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_338),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_355),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_364),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_343),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_329),
.A2(n_213),
.B1(n_234),
.B2(n_304),
.Y(n_442)
);

BUFx8_ASAP7_75t_SL g443 ( 
.A(n_362),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_443),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_413),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_413),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_387),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_438),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_431),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_442),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_412),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_435),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_412),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_397),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_399),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_405),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_427),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_414),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_406),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_410),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_406),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_414),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_410),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_410),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_440),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_391),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_436),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_391),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_417),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_406),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_391),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_404),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_386),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_386),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_429),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_419),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_419),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_393),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_402),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_394),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_402),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_421),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

AND3x2_ASAP7_75t_L g492 ( 
.A(n_384),
.B(n_323),
.C(n_313),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_422),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_390),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_422),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_422),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_384),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_R g498 ( 
.A(n_409),
.B(n_377),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_R g499 ( 
.A(n_409),
.B(n_378),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_385),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_385),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_428),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_396),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_415),
.Y(n_504)
);

BUFx10_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_426),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_396),
.A2(n_348),
.B(n_345),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_428),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_R g511 ( 
.A(n_425),
.B(n_362),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_439),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_451),
.B(n_415),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_454),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_474),
.B(n_455),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_469),
.B(n_439),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_486),
.B(n_365),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_472),
.B(n_302),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_475),
.B(n_415),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_444),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_457),
.B(n_361),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_485),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_490),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_415),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_508),
.B(n_320),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_488),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_502),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_509),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_448),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_481),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_448),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_466),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_497),
.B(n_430),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_512),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

BUFx10_ASAP7_75t_L g543 ( 
.A(n_445),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_507),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_460),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_505),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_500),
.B(n_501),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_494),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_489),
.B(n_229),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_463),
.B(n_425),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_494),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_R g552 ( 
.A(n_482),
.B(n_420),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_458),
.B(n_326),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_493),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_492),
.B(n_441),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_459),
.B(n_420),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_461),
.B(n_430),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_511),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_505),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_483),
.B(n_326),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_504),
.A2(n_425),
.B1(n_432),
.B2(n_434),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_488),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_503),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_511),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_510),
.B(n_432),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_495),
.B(n_231),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_513),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_465),
.B(n_432),
.Y(n_569)
);

AO21x2_ASAP7_75t_L g570 ( 
.A1(n_498),
.A2(n_499),
.B(n_476),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_447),
.B(n_344),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_496),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_514),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_480),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_480),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_488),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_491),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_453),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_491),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_491),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_491),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_479),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_452),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_478),
.B(n_344),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_484),
.B(n_441),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_456),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_487),
.Y(n_587)
);

AOI221xp5_ASAP7_75t_L g588 ( 
.A1(n_584),
.A2(n_354),
.B1(n_360),
.B2(n_350),
.C(n_351),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_558),
.B(n_535),
.Y(n_589)
);

AND2x6_ASAP7_75t_SL g590 ( 
.A(n_553),
.B(n_325),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_558),
.B(n_498),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_516),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_537),
.B(n_462),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_537),
.B(n_325),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_540),
.B(n_499),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_583),
.B(n_449),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_563),
.A2(n_392),
.B(n_386),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_556),
.B(n_550),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_576),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_527),
.B(n_464),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_543),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_540),
.B(n_434),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_534),
.B(n_467),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_543),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_518),
.B(n_434),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_528),
.B(n_430),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_530),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_541),
.B(n_468),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_546),
.B(n_471),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_556),
.A2(n_517),
.B1(n_531),
.B2(n_525),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_563),
.A2(n_525),
.B(n_517),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_562),
.B(n_433),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_547),
.B(n_522),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_562),
.B(n_433),
.Y(n_614)
);

NOR2x1p5_ASAP7_75t_L g615 ( 
.A(n_560),
.B(n_473),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_520),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_542),
.Y(n_617)
);

BUFx5_ASAP7_75t_L g618 ( 
.A(n_550),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_578),
.B(n_477),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_552),
.A2(n_437),
.B1(n_433),
.B2(n_292),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_539),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_523),
.B(n_411),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_559),
.B(n_233),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_555),
.B(n_433),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_L g625 ( 
.A(n_586),
.B(n_411),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_523),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_520),
.B(n_433),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_548),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_542),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_565),
.B(n_236),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_549),
.B(n_237),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_586),
.B(n_411),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_587),
.B(n_238),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_523),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_533),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_531),
.B(n_423),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_521),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_582),
.B(n_437),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_561),
.B(n_239),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_570),
.B(n_557),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_564),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_585),
.B(n_376),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_515),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_L g644 ( 
.A(n_571),
.B(n_567),
.C(n_554),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_566),
.B(n_529),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_533),
.Y(n_646)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_601),
.B(n_554),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_611),
.A2(n_577),
.B(n_533),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_636),
.A2(n_577),
.B(n_570),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_595),
.B(n_555),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_610),
.A2(n_607),
.B1(n_592),
.B2(n_640),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_636),
.A2(n_577),
.B(n_544),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_637),
.B(n_585),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_639),
.B(n_519),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_589),
.B(n_519),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_613),
.A2(n_524),
.B1(n_519),
.B2(n_532),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_596),
.B(n_572),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_591),
.A2(n_566),
.B(n_579),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_637),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_642),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_593),
.B(n_572),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_624),
.A2(n_524),
.B(n_532),
.C(n_568),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_594),
.B(n_524),
.Y(n_663)
);

AOI21xp33_ASAP7_75t_L g664 ( 
.A1(n_631),
.A2(n_532),
.B(n_573),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_602),
.B(n_536),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_645),
.B(n_538),
.Y(n_666)
);

O2A1O1Ixp33_ASAP7_75t_SL g667 ( 
.A1(n_612),
.A2(n_581),
.B(n_580),
.C(n_575),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_614),
.A2(n_551),
.B1(n_545),
.B2(n_574),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_598),
.A2(n_398),
.B(n_392),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_623),
.B(n_526),
.Y(n_670)
);

CKINVDCx10_ASAP7_75t_R g671 ( 
.A(n_590),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_645),
.A2(n_398),
.B(n_392),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_605),
.A2(n_353),
.B(n_356),
.C(n_358),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_628),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_625),
.B(n_526),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_634),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_632),
.B(n_246),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_627),
.A2(n_569),
.B(n_550),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_641),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_638),
.A2(n_398),
.B(n_392),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_616),
.B(n_249),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_615),
.B(n_550),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_643),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_644),
.A2(n_569),
.B1(n_298),
.B2(n_295),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_617),
.A2(n_569),
.B1(n_437),
.B2(n_423),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_630),
.B(n_250),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_626),
.A2(n_398),
.B(n_392),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_633),
.B(n_569),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_606),
.A2(n_401),
.B(n_400),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_620),
.A2(n_423),
.B(n_424),
.C(n_416),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_634),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_629),
.B(n_416),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_599),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_650),
.B(n_619),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_671),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_657),
.B(n_621),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_670),
.A2(n_604),
.B1(n_600),
.B2(n_603),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_662),
.A2(n_654),
.B(n_664),
.C(n_656),
.Y(n_698)
);

NAND2x2_ASAP7_75t_L g699 ( 
.A(n_663),
.B(n_608),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_674),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_666),
.B(n_588),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_679),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_661),
.B(n_609),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_653),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_683),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_651),
.A2(n_635),
.B1(n_634),
.B2(n_646),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_659),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_682),
.B(n_655),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_SL g709 ( 
.A(n_686),
.B(n_254),
.C(n_251),
.Y(n_709)
);

O2A1O1Ixp5_ASAP7_75t_L g710 ( 
.A1(n_688),
.A2(n_599),
.B(n_646),
.C(n_597),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_676),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_660),
.B(n_622),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_651),
.A2(n_622),
.B1(n_300),
.B2(n_291),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_665),
.B(n_424),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_682),
.Y(n_715)
);

OAI22x1_ASAP7_75t_L g716 ( 
.A1(n_684),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_681),
.B(n_618),
.Y(n_717)
);

OA22x2_ASAP7_75t_L g718 ( 
.A1(n_675),
.A2(n_260),
.B1(n_267),
.B2(n_268),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_649),
.A2(n_693),
.B1(n_685),
.B2(n_647),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_692),
.B(n_271),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_691),
.B(n_388),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_676),
.B(n_618),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_691),
.B(n_618),
.Y(n_723)
);

O2A1O1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_673),
.A2(n_388),
.B(n_389),
.C(n_408),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_668),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_668),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_658),
.B(n_618),
.Y(n_727)
);

AO21x1_ASAP7_75t_L g728 ( 
.A1(n_648),
.A2(n_408),
.B(n_389),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_677),
.B(n_273),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_690),
.B(n_275),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_667),
.B(n_278),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_652),
.A2(n_618),
.B(n_398),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_678),
.A2(n_437),
.B(n_406),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_672),
.B(n_279),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_680),
.B(n_280),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_689),
.B(n_281),
.Y(n_736)
);

BUFx5_ASAP7_75t_L g737 ( 
.A(n_726),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_702),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_725),
.Y(n_739)
);

AND2x6_ASAP7_75t_L g740 ( 
.A(n_717),
.B(n_708),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_727),
.A2(n_669),
.B(n_687),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_707),
.Y(n_742)
);

OAI21x1_ASAP7_75t_SL g743 ( 
.A1(n_719),
.A2(n_400),
.B(n_401),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_694),
.B(n_696),
.Y(n_744)
);

AO31x2_ASAP7_75t_L g745 ( 
.A1(n_728),
.A2(n_403),
.A3(n_407),
.B(n_2),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_715),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_698),
.B(n_305),
.C(n_285),
.Y(n_747)
);

NAND2x1p5_ASAP7_75t_L g748 ( 
.A(n_711),
.B(n_403),
.Y(n_748)
);

AOI221x1_ASAP7_75t_L g749 ( 
.A1(n_731),
.A2(n_437),
.B1(n_418),
.B2(n_407),
.C(n_4),
.Y(n_749)
);

CKINVDCx11_ASAP7_75t_R g750 ( 
.A(n_699),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_704),
.B(n_283),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_700),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_705),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_721),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_704),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_701),
.B(n_286),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_703),
.B(n_301),
.Y(n_757)
);

AO21x2_ASAP7_75t_L g758 ( 
.A1(n_733),
.A2(n_418),
.B(n_309),
.Y(n_758)
);

AO32x2_ASAP7_75t_L g759 ( 
.A1(n_706),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_759)
);

AO21x2_ASAP7_75t_L g760 ( 
.A1(n_732),
.A2(n_418),
.B(n_395),
.Y(n_760)
);

OAI21x1_ASAP7_75t_L g761 ( 
.A1(n_710),
.A2(n_418),
.B(n_395),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_SL g762 ( 
.A(n_695),
.B(n_418),
.Y(n_762)
);

AOI21xp33_ASAP7_75t_L g763 ( 
.A1(n_734),
.A2(n_6),
.B(n_7),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_697),
.A2(n_395),
.B1(n_7),
.B2(n_8),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_712),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_711),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_736),
.A2(n_395),
.B(n_100),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_706),
.A2(n_97),
.B(n_192),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_721),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_708),
.B(n_6),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_714),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_720),
.B(n_8),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_718),
.B(n_9),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_729),
.B(n_10),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_718),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_709),
.B(n_28),
.Y(n_776)
);

NOR4xp25_ASAP7_75t_L g777 ( 
.A(n_713),
.B(n_11),
.C(n_14),
.D(n_15),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_716),
.B(n_14),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_730),
.B(n_15),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_735),
.B(n_16),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_724),
.B(n_16),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_723),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_722),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_746),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_741),
.A2(n_117),
.B(n_189),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_761),
.A2(n_17),
.B(n_18),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_755),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_749),
.A2(n_118),
.B(n_188),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_752),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_747),
.A2(n_780),
.B(n_772),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_739),
.B(n_19),
.Y(n_791)
);

CKINVDCx6p67_ASAP7_75t_R g792 ( 
.A(n_750),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_743),
.A2(n_768),
.B(n_767),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_774),
.A2(n_20),
.B(n_22),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_739),
.A2(n_119),
.B(n_185),
.Y(n_795)
);

CKINVDCx11_ASAP7_75t_R g796 ( 
.A(n_783),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_766),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_779),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_771),
.B(n_24),
.Y(n_799)
);

AO21x2_ASAP7_75t_L g800 ( 
.A1(n_758),
.A2(n_25),
.B(n_29),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_753),
.A2(n_30),
.B(n_32),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_737),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_742),
.B(n_33),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_752),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_737),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_765),
.Y(n_806)
);

OA21x2_ASAP7_75t_L g807 ( 
.A1(n_753),
.A2(n_34),
.B(n_35),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_738),
.A2(n_37),
.B(n_38),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_737),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_758),
.A2(n_40),
.B(n_41),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_760),
.A2(n_777),
.B(n_781),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_737),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_748),
.A2(n_42),
.B(n_47),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_740),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_754),
.B(n_48),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_751),
.B(n_52),
.Y(n_816)
);

NAND2x1_ASAP7_75t_L g817 ( 
.A(n_740),
.B(n_54),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_766),
.B(n_744),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_769),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_763),
.B(n_58),
.C(n_59),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_770),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_784),
.B(n_757),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_790),
.A2(n_764),
.B1(n_778),
.B2(n_776),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_788),
.A2(n_810),
.B(n_802),
.Y(n_824)
);

INVxp67_ASAP7_75t_SL g825 ( 
.A(n_802),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_793),
.A2(n_775),
.B(n_737),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_810),
.A2(n_773),
.B(n_760),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_788),
.A2(n_762),
.B(n_756),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_789),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_804),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_819),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_809),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_796),
.Y(n_833)
);

NOR2x1_ASAP7_75t_SL g834 ( 
.A(n_812),
.B(n_759),
.Y(n_834)
);

OAI21x1_ASAP7_75t_L g835 ( 
.A1(n_785),
.A2(n_745),
.B(n_782),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_820),
.A2(n_740),
.B(n_759),
.Y(n_836)
);

AO31x2_ASAP7_75t_L g837 ( 
.A1(n_814),
.A2(n_791),
.A3(n_745),
.B(n_786),
.Y(n_837)
);

OAI21x1_ASAP7_75t_SL g838 ( 
.A1(n_794),
.A2(n_791),
.B(n_799),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_821),
.B(n_759),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_787),
.B(n_740),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_805),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_805),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_796),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_819),
.B(n_745),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_798),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_807),
.A2(n_67),
.B(n_68),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_806),
.B(n_70),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_807),
.A2(n_73),
.B(n_76),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_818),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_832),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_824),
.A2(n_786),
.B(n_801),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_829),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_831),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_841),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_830),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_833),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_841),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_842),
.Y(n_858)
);

BUFx2_ASAP7_75t_SL g859 ( 
.A(n_843),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_825),
.Y(n_860)
);

BUFx2_ASAP7_75t_SL g861 ( 
.A(n_843),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_842),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_825),
.B(n_807),
.Y(n_863)
);

INVx8_ASAP7_75t_L g864 ( 
.A(n_833),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_849),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_844),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_866),
.B(n_839),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_859),
.A2(n_823),
.B1(n_845),
.B2(n_836),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_864),
.B(n_822),
.Y(n_869)
);

OAI21xp33_ASAP7_75t_L g870 ( 
.A1(n_863),
.A2(n_845),
.B(n_798),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_864),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_855),
.B(n_837),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_SL g873 ( 
.A1(n_860),
.A2(n_848),
.B(n_846),
.C(n_799),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_859),
.A2(n_818),
.B1(n_828),
.B2(n_792),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_856),
.A2(n_838),
.B1(n_811),
.B2(n_840),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_861),
.A2(n_817),
.B1(n_803),
.B2(n_847),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_857),
.B(n_837),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_871),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_872),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_877),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_874),
.B(n_856),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_867),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_869),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_875),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_881),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_882),
.B(n_852),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_878),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_878),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_880),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_884),
.B(n_870),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_887),
.B(n_883),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_L g892 ( 
.A(n_890),
.B(n_868),
.C(n_881),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_SL g893 ( 
.A1(n_885),
.A2(n_876),
.B(n_863),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_888),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_L g895 ( 
.A(n_889),
.B(n_873),
.C(n_879),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_891),
.B(n_885),
.Y(n_896)
);

NOR2x1_ASAP7_75t_L g897 ( 
.A(n_892),
.B(n_856),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_894),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_893),
.B(n_861),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_895),
.B(n_864),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_896),
.B(n_886),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_898),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_899),
.B(n_869),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_897),
.B(n_864),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_900),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_896),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_902),
.Y(n_907)
);

OAI22xp33_ASAP7_75t_L g908 ( 
.A1(n_906),
.A2(n_866),
.B1(n_853),
.B2(n_865),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_906),
.B(n_855),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_905),
.B(n_852),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_904),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_904),
.A2(n_811),
.B1(n_800),
.B2(n_851),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_901),
.B(n_860),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_901),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_914),
.B(n_903),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_911),
.B(n_854),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_907),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_910),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_909),
.B(n_854),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_913),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_908),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_912),
.B(n_858),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_SL g923 ( 
.A1(n_914),
.A2(n_803),
.B(n_815),
.Y(n_923)
);

OAI22x1_ASAP7_75t_L g924 ( 
.A1(n_921),
.A2(n_815),
.B1(n_853),
.B2(n_797),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_915),
.B(n_854),
.Y(n_925)
);

AOI222xp33_ASAP7_75t_L g926 ( 
.A1(n_917),
.A2(n_816),
.B1(n_834),
.B2(n_851),
.C1(n_827),
.C2(n_835),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_920),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_918),
.A2(n_813),
.B(n_795),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_916),
.B(n_850),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_919),
.B(n_923),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_922),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_915),
.Y(n_932)
);

OAI22xp33_ASAP7_75t_L g933 ( 
.A1(n_921),
.A2(n_831),
.B1(n_850),
.B2(n_862),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_932),
.A2(n_835),
.B(n_826),
.C(n_797),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_927),
.A2(n_930),
.B1(n_933),
.B2(n_924),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_931),
.A2(n_925),
.B(n_929),
.C(n_926),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_926),
.B(n_819),
.C(n_831),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_928),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_932),
.A2(n_800),
.B(n_862),
.C(n_786),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_932),
.A2(n_831),
.B1(n_819),
.B2(n_844),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_932),
.B(n_844),
.Y(n_941)
);

NAND4xp25_ASAP7_75t_L g942 ( 
.A(n_932),
.B(n_77),
.C(n_79),
.D(n_82),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_932),
.A2(n_826),
.B(n_808),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_935),
.A2(n_85),
.B(n_88),
.Y(n_944)
);

AOI322xp5_ASAP7_75t_L g945 ( 
.A1(n_941),
.A2(n_837),
.A3(n_91),
.B1(n_94),
.B2(n_95),
.C1(n_105),
.C2(n_108),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_936),
.B(n_90),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_L g947 ( 
.A(n_942),
.B(n_111),
.C(n_114),
.Y(n_947)
);

AOI322xp5_ASAP7_75t_L g948 ( 
.A1(n_938),
.A2(n_837),
.A3(n_122),
.B1(n_125),
.B2(n_126),
.C1(n_127),
.C2(n_129),
.Y(n_948)
);

AOI221xp5_ASAP7_75t_L g949 ( 
.A1(n_937),
.A2(n_121),
.B1(n_130),
.B2(n_134),
.C(n_135),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_940),
.A2(n_136),
.B(n_139),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_SL g951 ( 
.A(n_944),
.B(n_934),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_946),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_945),
.Y(n_953)
);

NAND3x1_ASAP7_75t_SL g954 ( 
.A(n_952),
.B(n_949),
.C(n_948),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_951),
.A2(n_950),
.B(n_947),
.C(n_939),
.Y(n_955)
);

NOR2x1_ASAP7_75t_L g956 ( 
.A(n_955),
.B(n_953),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_954),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_957),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_956),
.B(n_943),
.Y(n_959)
);

OAI211xp5_ASAP7_75t_L g960 ( 
.A1(n_958),
.A2(n_141),
.B(n_143),
.C(n_144),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_960),
.B(n_959),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_961),
.Y(n_962)
);

BUFx2_ASAP7_75t_SL g963 ( 
.A(n_962),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_SL g964 ( 
.A1(n_963),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_964),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_965),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_965),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_966),
.A2(n_148),
.B(n_149),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_968),
.B(n_967),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_R g970 ( 
.A1(n_969),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_970)
);

AO21x2_ASAP7_75t_L g971 ( 
.A1(n_970),
.A2(n_160),
.B(n_161),
.Y(n_971)
);

OAI22xp33_ASAP7_75t_L g972 ( 
.A1(n_971),
.A2(n_162),
.B1(n_165),
.B2(n_169),
.Y(n_972)
);

AOI211xp5_ASAP7_75t_L g973 ( 
.A1(n_972),
.A2(n_170),
.B(n_171),
.C(n_175),
.Y(n_973)
);


endmodule