module fake_jpeg_31814_n_179 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

INVx8_ASAP7_75t_SL g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_74),
.Y(n_86)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_63),
.Y(n_73)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_23),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_0),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_84),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_48),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_59),
.B1(n_52),
.B2(n_66),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_91),
.B1(n_81),
.B2(n_83),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_59),
.B1(n_65),
.B2(n_51),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_65),
.B1(n_60),
.B2(n_67),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_49),
.B1(n_52),
.B2(n_66),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_93),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_9),
.Y(n_133)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_125),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_131),
.B1(n_129),
.B2(n_115),
.Y(n_143)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_29),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_12),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_55),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_5),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_5),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_7),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_133),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_11),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_42),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_33),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_46),
.B1(n_14),
.B2(n_16),
.Y(n_137)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_141),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_134),
.A2(n_19),
.B(n_20),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_22),
.B(n_24),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_25),
.C(n_26),
.Y(n_147)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_151),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_30),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_34),
.B(n_35),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_37),
.Y(n_158)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_162),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_151),
.C(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_148),
.C(n_143),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_168),
.B(n_169),
.C(n_138),
.D(n_157),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_147),
.C(n_144),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_146),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_166),
.B(n_170),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_156),
.A3(n_159),
.B1(n_164),
.B2(n_139),
.C1(n_120),
.C2(n_136),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_164),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_116),
.Y(n_179)
);


endmodule