module fake_ariane_341_n_1985 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1985);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1985;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_113),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_68),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_35),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_116),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_89),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_65),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_77),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_54),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_115),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_112),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_17),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_96),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_60),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_44),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_19),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_109),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_154),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_158),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_32),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_104),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_91),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_196),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_35),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_64),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_67),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_32),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_127),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_10),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_175),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_141),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_185),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_50),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_166),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_55),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_76),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_59),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_42),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_33),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_95),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_71),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_86),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_143),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_111),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_137),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_6),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_117),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_73),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_130),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_178),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_102),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_120),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_3),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_36),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_203),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_3),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_85),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_192),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_72),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_88),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_74),
.Y(n_282)
);

INVxp33_ASAP7_75t_R g283 ( 
.A(n_197),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_43),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_161),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_200),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_165),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_58),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_25),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_8),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_114),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_169),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_28),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_34),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_157),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_126),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_21),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_78),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_101),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_64),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_40),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_65),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_138),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_17),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_14),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_183),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_56),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_69),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_133),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_69),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_131),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_121),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_29),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_11),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_99),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_53),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_93),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_1),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_31),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_38),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_8),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_62),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_21),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_198),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_10),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_136),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_66),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_43),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_60),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_70),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_63),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_36),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_1),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_181),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_14),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_82),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_68),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_84),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_207),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_180),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_105),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_162),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_13),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_132),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_29),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_46),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_119),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_28),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_128),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_80),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_156),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_147),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_83),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_204),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_7),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_90),
.Y(n_356)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_50),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_144),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_30),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_148),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_20),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_188),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_87),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_155),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_170),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_63),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_5),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_66),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_206),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_54),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_40),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_199),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_110),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_15),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_15),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_81),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_25),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_122),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_16),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_26),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_62),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_168),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_146),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_159),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_135),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_124),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_195),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_58),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_149),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_75),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_67),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_30),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_123),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_201),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_98),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_6),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_12),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_41),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_174),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_145),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_38),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_51),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_49),
.Y(n_403)
);

BUFx4f_ASAP7_75t_SL g404 ( 
.A(n_23),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_152),
.Y(n_405)
);

BUFx5_ASAP7_75t_L g406 ( 
.A(n_12),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_0),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_92),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_160),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_45),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_176),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_20),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_118),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_357),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_297),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_337),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_297),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_357),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_392),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_219),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_225),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_252),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_392),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_229),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_276),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_351),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_229),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_406),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_282),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_229),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_400),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_220),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_267),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_217),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_314),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_323),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_325),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_284),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_331),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_288),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_406),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_229),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_210),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_248),
.B(n_0),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_289),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_229),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_340),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_290),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_241),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_264),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_370),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_241),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_264),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_210),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_294),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_300),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_301),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_266),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_307),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_310),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_274),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_274),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_277),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_316),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_375),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_277),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_213),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_318),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_404),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_243),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_328),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_313),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_329),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_266),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_299),
.B(n_2),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_338),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_313),
.Y(n_489)
);

INVxp33_ASAP7_75t_SL g490 ( 
.A(n_213),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_333),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_338),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_352),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_335),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_352),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_368),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_224),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_224),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_345),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_368),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_401),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_344),
.B(n_2),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_R g505 ( 
.A(n_263),
.B(n_205),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_348),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_390),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_226),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_231),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_390),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_226),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_231),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_355),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_208),
.B(n_4),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_227),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_214),
.B(n_4),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_218),
.Y(n_518)
);

INVx6_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_464),
.B(n_244),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_257),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_429),
.B(n_221),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_432),
.B(n_222),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_414),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_489),
.B(n_265),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_441),
.B(n_223),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_425),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_415),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_425),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_488),
.B(n_230),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_439),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_459),
.B(n_235),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_518),
.B(n_422),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_416),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_418),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_470),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_421),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_423),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_423),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_428),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_428),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_509),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_462),
.B(n_238),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_433),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_433),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_434),
.A2(n_246),
.B(n_245),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_435),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_518),
.B(n_275),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_509),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_459),
.B(n_283),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_436),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_438),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_516),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_462),
.B(n_293),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_438),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_440),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_427),
.B(n_302),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_419),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_440),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_488),
.B(n_255),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_465),
.B(n_258),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_452),
.B(n_235),
.Y(n_574)
);

BUFx8_ASAP7_75t_L g575 ( 
.A(n_465),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_452),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_453),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_453),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_454),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_454),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_510),
.B(n_304),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_510),
.B(n_305),
.Y(n_582)
);

BUFx8_ASAP7_75t_L g583 ( 
.A(n_431),
.Y(n_583)
);

BUFx8_ASAP7_75t_L g584 ( 
.A(n_431),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_458),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_458),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_513),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_513),
.B(n_319),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_492),
.B(n_260),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_444),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_461),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_461),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_473),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_473),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_474),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_474),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_475),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_492),
.B(n_320),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_475),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_466),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_478),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_542),
.Y(n_602)
);

OAI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_589),
.A2(n_508),
.B1(n_455),
.B2(n_490),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_542),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_536),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_540),
.B(n_508),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_540),
.B(n_539),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_589),
.B(n_479),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_542),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_540),
.B(n_417),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_539),
.B(n_449),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_555),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_583),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_535),
.B(n_451),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_539),
.A2(n_487),
.B1(n_504),
.B2(n_456),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_555),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_572),
.B(n_457),
.Y(n_617)
);

INVx4_ASAP7_75t_SL g618 ( 
.A(n_574),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_543),
.B(n_460),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_590),
.B(n_481),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_SL g621 ( 
.A(n_590),
.B(n_467),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_558),
.B(n_420),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_555),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_543),
.B(n_468),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_566),
.A2(n_517),
.B1(n_515),
.B2(n_498),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_543),
.B(n_469),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_557),
.Y(n_627)
);

OR2x6_ASAP7_75t_L g628 ( 
.A(n_569),
.B(n_445),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_557),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_557),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_523),
.B(n_471),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_562),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_SL g633 ( 
.A(n_570),
.B(n_476),
.C(n_472),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_562),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_566),
.A2(n_512),
.B1(n_497),
.B2(n_493),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_567),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_567),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_567),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_527),
.B(n_529),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_570),
.Y(n_641)
);

AND2x4_ASAP7_75t_SL g642 ( 
.A(n_551),
.B(n_486),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_578),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g644 ( 
.A(n_551),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_527),
.B(n_480),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_529),
.B(n_483),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_566),
.A2(n_511),
.B1(n_495),
.B2(n_322),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_547),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_536),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_558),
.B(n_588),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_569),
.B(n_482),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_531),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_547),
.Y(n_653)
);

AND3x1_ASAP7_75t_L g654 ( 
.A(n_559),
.B(n_600),
.C(n_598),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_547),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_560),
.A2(n_559),
.B1(n_600),
.B2(n_379),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_491),
.C(n_485),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_565),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_523),
.B(n_494),
.Y(n_660)
);

INVx4_ASAP7_75t_SL g661 ( 
.A(n_574),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_547),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_558),
.B(n_478),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_598),
.B(n_499),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_578),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_531),
.B(n_507),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_588),
.B(n_484),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_588),
.B(n_484),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_526),
.B(n_514),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_526),
.B(n_424),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_538),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_569),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_225),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_538),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_521),
.B(n_426),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_547),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_536),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_566),
.A2(n_402),
.B1(n_380),
.B2(n_377),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_538),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_588),
.B(n_581),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_530),
.B(n_430),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_547),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_538),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_566),
.A2(n_327),
.B1(n_371),
.B2(n_346),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_521),
.B(n_437),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_588),
.B(n_311),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_533),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_571),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_530),
.B(n_477),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_579),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_583),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_571),
.B(n_225),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_583),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_556),
.B(n_262),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_579),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_521),
.B(n_211),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_528),
.B(n_211),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_571),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_528),
.B(n_212),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_571),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_565),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_580),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_571),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_533),
.B(n_442),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_537),
.B(n_270),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_581),
.A2(n_321),
.B1(n_343),
.B2(n_332),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_537),
.B(n_209),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_585),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_541),
.B(n_250),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_541),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_585),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_586),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_522),
.A2(n_308),
.B1(n_253),
.B2(n_251),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_528),
.B(n_212),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_571),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_571),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_586),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_522),
.B(n_215),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_546),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_544),
.B(n_272),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_577),
.Y(n_722)
);

AND3x2_ASAP7_75t_L g723 ( 
.A(n_560),
.B(n_330),
.C(n_311),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_577),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_544),
.B(n_273),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_545),
.B(n_280),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_545),
.B(n_286),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_548),
.B(n_295),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_581),
.B(n_496),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_548),
.B(n_291),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_549),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_549),
.B(n_393),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_577),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_577),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_577),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_577),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_550),
.B(n_215),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_550),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_577),
.Y(n_739)
);

OR2x6_ASAP7_75t_L g740 ( 
.A(n_581),
.B(n_496),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_546),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_522),
.B(n_582),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_553),
.B(n_292),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_522),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_583),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_575),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_575),
.B(n_216),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_546),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_553),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_575),
.B(n_216),
.Y(n_750)
);

AND2x2_ASAP7_75t_SL g751 ( 
.A(n_556),
.B(n_330),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_546),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_554),
.B(n_228),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_554),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_631),
.B(n_575),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_608),
.B(n_576),
.Y(n_756)
);

BUFx12f_ASAP7_75t_SL g757 ( 
.A(n_628),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_672),
.A2(n_591),
.B1(n_587),
.B2(n_256),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_652),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_659),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_748),
.B(n_576),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_642),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_652),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_748),
.B(n_576),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_L g765 ( 
.A(n_645),
.B(n_576),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_605),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_604),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_604),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_660),
.A2(n_669),
.B1(n_672),
.B2(n_670),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_613),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_748),
.B(n_561),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_741),
.B(n_752),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_687),
.Y(n_773)
);

NAND2x1p5_ASAP7_75t_L g774 ( 
.A(n_746),
.B(n_607),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_687),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_614),
.B(n_561),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_701),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_711),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_617),
.B(n_563),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_646),
.B(n_563),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_741),
.B(n_564),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_689),
.B(n_564),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_623),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_607),
.A2(n_751),
.B1(n_686),
.B2(n_650),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_681),
.B(n_568),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_666),
.B(n_568),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_615),
.A2(n_584),
.B1(n_582),
.B2(n_574),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_606),
.B(n_680),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_752),
.B(n_574),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_611),
.A2(n_584),
.B1(n_582),
.B2(n_574),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_741),
.B(n_711),
.Y(n_791)
);

BUFx6f_ASAP7_75t_SL g792 ( 
.A(n_641),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_628),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_651),
.B(n_582),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_680),
.B(n_591),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_731),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_720),
.A2(n_556),
.B(n_574),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_731),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_623),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_690),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_708),
.B(n_591),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_605),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_658),
.B(n_552),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_710),
.B(n_726),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_727),
.B(n_591),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_605),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_745),
.B(n_584),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_690),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_695),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_695),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_728),
.B(n_552),
.Y(n_811)
);

OR2x6_ASAP7_75t_L g812 ( 
.A(n_628),
.B(n_584),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_732),
.B(n_573),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_751),
.A2(n_556),
.B1(n_587),
.B2(n_574),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_628),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_642),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_702),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_650),
.B(n_573),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_744),
.B(n_593),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_641),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_651),
.B(n_593),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_651),
.B(n_596),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_702),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_738),
.B(n_536),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_664),
.B(n_536),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_705),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_651),
.B(n_596),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_738),
.B(n_536),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_619),
.B(n_536),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_749),
.B(n_754),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_667),
.B(n_597),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_627),
.Y(n_832)
);

NAND2x1_ASAP7_75t_L g833 ( 
.A(n_686),
.B(n_519),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_629),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_705),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_667),
.B(n_597),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_624),
.B(n_594),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_640),
.A2(n_592),
.B(n_501),
.C(n_506),
.Y(n_838)
);

AO221x1_ASAP7_75t_L g839 ( 
.A1(n_657),
.A2(n_279),
.B1(n_225),
.B2(n_386),
.C(n_296),
.Y(n_839)
);

INVx8_ASAP7_75t_L g840 ( 
.A(n_686),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_644),
.B(n_443),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_686),
.Y(n_842)
);

AND2x2_ASAP7_75t_SL g843 ( 
.A(n_751),
.B(n_373),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_749),
.B(n_228),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_709),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_668),
.B(n_592),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_629),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_696),
.B(n_594),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_668),
.B(n_592),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_636),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_636),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_605),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_610),
.B(n_446),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_712),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_686),
.A2(n_556),
.B1(n_574),
.B2(n_595),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_742),
.A2(n_247),
.B1(n_242),
.B2(n_259),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_754),
.B(n_232),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_686),
.A2(n_574),
.B1(n_599),
.B2(n_595),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_729),
.B(n_594),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_663),
.B(n_594),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_643),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_663),
.B(n_594),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_740),
.B(n_594),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_697),
.B(n_595),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_699),
.B(n_595),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_686),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_605),
.B(n_232),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_740),
.A2(n_236),
.B1(n_413),
.B2(n_411),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_712),
.Y(n_869)
);

BUFx8_ASAP7_75t_L g870 ( 
.A(n_610),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_635),
.B(n_675),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_641),
.Y(n_872)
);

NAND2xp33_ASAP7_75t_L g873 ( 
.A(n_674),
.B(n_233),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_740),
.B(n_595),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_713),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_740),
.B(n_595),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_737),
.B(n_595),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_622),
.B(n_704),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_643),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_715),
.B(n_599),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_753),
.B(n_599),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_622),
.B(n_447),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_706),
.B(n_599),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_719),
.B(n_599),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_647),
.B(n_448),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_685),
.B(n_626),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_602),
.A2(n_374),
.B(n_253),
.C(n_251),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_721),
.B(n_599),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_725),
.B(n_599),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_698),
.A2(n_525),
.B(n_524),
.Y(n_890)
);

INVx8_ASAP7_75t_L g891 ( 
.A(n_613),
.Y(n_891)
);

AND2x6_ASAP7_75t_SL g892 ( 
.A(n_620),
.B(n_500),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_655),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_654),
.Y(n_894)
);

OAI221xp5_ASAP7_75t_L g895 ( 
.A1(n_625),
.A2(n_247),
.B1(n_361),
.B2(n_366),
.C(n_367),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_730),
.B(n_601),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_649),
.B(n_233),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_649),
.B(n_234),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_655),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_602),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_L g901 ( 
.A(n_633),
.B(n_621),
.C(n_603),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_L g902 ( 
.A(n_674),
.B(n_679),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_713),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_743),
.B(n_601),
.Y(n_904)
);

NOR2xp67_ASAP7_75t_L g905 ( 
.A(n_693),
.B(n_746),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_714),
.B(n_450),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_718),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_679),
.B(n_601),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_671),
.B(n_601),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_609),
.Y(n_910)
);

AND2x6_ASAP7_75t_SL g911 ( 
.A(n_654),
.B(n_500),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_609),
.A2(n_308),
.B(n_242),
.C(n_237),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_671),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_683),
.B(n_601),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_742),
.A2(n_227),
.B1(n_237),
.B2(n_412),
.Y(n_915)
);

NAND3x1_ASAP7_75t_L g916 ( 
.A(n_714),
.B(n_463),
.C(n_501),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_691),
.B(n_502),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_707),
.B(n_256),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_683),
.B(n_601),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_612),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_612),
.Y(n_921)
);

INVx8_ASAP7_75t_L g922 ( 
.A(n_693),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_691),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_616),
.B(n_601),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_769),
.B(n_723),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_760),
.B(n_603),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_830),
.A2(n_700),
.B(n_698),
.Y(n_927)
);

BUFx4f_ASAP7_75t_L g928 ( 
.A(n_812),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_782),
.B(n_616),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_756),
.B(n_630),
.Y(n_930)
);

AO21x2_ASAP7_75t_L g931 ( 
.A1(n_830),
.A2(n_632),
.B(n_630),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_785),
.A2(n_716),
.B(n_700),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_756),
.B(n_632),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_843),
.A2(n_878),
.B1(n_871),
.B2(n_784),
.Y(n_934)
);

BUFx4f_ASAP7_75t_L g935 ( 
.A(n_812),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_776),
.A2(n_637),
.B(n_665),
.C(n_639),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_777),
.B(n_853),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_800),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_786),
.A2(n_722),
.B(n_716),
.Y(n_939)
);

O2A1O1Ixp5_ASAP7_75t_L g940 ( 
.A1(n_776),
.A2(n_718),
.B(n_703),
.C(n_734),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_779),
.A2(n_634),
.B(n_638),
.C(n_639),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_779),
.A2(n_665),
.B(n_638),
.C(n_662),
.Y(n_942)
);

AOI21x1_ASAP7_75t_L g943 ( 
.A1(n_771),
.A2(n_724),
.B(n_722),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_SL g944 ( 
.A1(n_885),
.A2(n_259),
.B1(n_359),
.B2(n_398),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_L g945 ( 
.A(n_840),
.B(n_648),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_788),
.B(n_747),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_797),
.A2(n_733),
.B(n_724),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_804),
.B(n_750),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_811),
.B(n_678),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_757),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_882),
.B(n_684),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_843),
.A2(n_784),
.B1(n_809),
.B2(n_808),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_810),
.A2(n_703),
.B1(n_734),
.B2(n_648),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_817),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_886),
.A2(n_703),
.B1(n_734),
.B2(n_656),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_772),
.A2(n_735),
.B(n_733),
.Y(n_956)
);

AO21x1_ASAP7_75t_L g957 ( 
.A1(n_829),
.A2(n_694),
.B(n_692),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_812),
.B(n_694),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_813),
.B(n_648),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_803),
.A2(n_682),
.B(n_656),
.C(n_662),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_763),
.B(n_798),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_772),
.A2(n_736),
.B(n_735),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_818),
.B(n_653),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_840),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_823),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_799),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_803),
.B(n_653),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_765),
.A2(n_828),
.B(n_824),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_861),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_763),
.B(n_649),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_895),
.A2(n_361),
.B(n_359),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_794),
.B(n_502),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_758),
.A2(n_682),
.B(n_656),
.C(n_717),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_824),
.A2(n_828),
.B(n_780),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_798),
.B(n_649),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_826),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_835),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_845),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_821),
.B(n_653),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_761),
.A2(n_739),
.B(n_736),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_814),
.A2(n_694),
.B(n_739),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_841),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_761),
.A2(n_764),
.B(n_781),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_L g984 ( 
.A(n_901),
.B(n_367),
.C(n_366),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_822),
.B(n_662),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_807),
.B(n_793),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_827),
.B(n_676),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_861),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_764),
.A2(n_717),
.B(n_682),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_891),
.B(n_503),
.Y(n_990)
);

AOI21xp33_ASAP7_75t_L g991 ( 
.A1(n_755),
.A2(n_688),
.B(n_676),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_SL g992 ( 
.A(n_887),
.B(n_381),
.C(n_374),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_854),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_869),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_875),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_758),
.B(n_649),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_815),
.A2(n_717),
.B1(n_688),
.B2(n_676),
.Y(n_997)
);

NOR3xp33_ASAP7_75t_L g998 ( 
.A(n_894),
.B(n_388),
.C(n_381),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_781),
.A2(n_688),
.B(n_677),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_840),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_819),
.B(n_795),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_831),
.B(n_677),
.Y(n_1002)
);

BUFx12f_ASAP7_75t_L g1003 ( 
.A(n_870),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_836),
.B(n_677),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_829),
.A2(n_673),
.B(n_525),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_903),
.B(n_677),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_891),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_767),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_770),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_886),
.B(n_677),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_907),
.B(n_388),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_846),
.B(n_391),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_902),
.A2(n_525),
.B(n_524),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_906),
.B(n_391),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_877),
.A2(n_524),
.B(n_317),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_849),
.B(n_396),
.Y(n_1016)
);

A2O1A1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_825),
.A2(n_383),
.B(n_315),
.C(n_347),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_766),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_842),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_820),
.B(n_396),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_872),
.B(n_762),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_791),
.A2(n_387),
.B(n_324),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_759),
.B(n_397),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_766),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_842),
.B(n_618),
.Y(n_1025)
);

O2A1O1Ixp5_ASAP7_75t_L g1026 ( 
.A1(n_867),
.A2(n_384),
.B(n_362),
.C(n_363),
.Y(n_1026)
);

NOR3xp33_ASAP7_75t_L g1027 ( 
.A(n_856),
.B(n_915),
.C(n_857),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_860),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_816),
.B(n_397),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_773),
.B(n_398),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_775),
.B(n_407),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_881),
.A2(n_249),
.B(n_236),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_917),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_787),
.A2(n_249),
.B1(n_413),
.B2(n_234),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_801),
.A2(n_254),
.B(n_239),
.Y(n_1035)
);

NOR2x1p5_ASAP7_75t_L g1036 ( 
.A(n_923),
.B(n_407),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_834),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_908),
.A2(n_395),
.B(n_376),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_866),
.B(n_618),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_791),
.A2(n_360),
.B(n_369),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_L g1041 ( 
.A(n_868),
.B(n_410),
.C(n_412),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_862),
.A2(n_534),
.B(n_532),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_834),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_805),
.A2(n_534),
.B(n_532),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_917),
.B(n_918),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_778),
.B(n_410),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_866),
.B(n_618),
.Y(n_1047)
);

NOR2xp67_ASAP7_75t_L g1048 ( 
.A(n_905),
.B(n_503),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_766),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_924),
.A2(n_534),
.B(n_532),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_859),
.A2(n_389),
.B1(n_373),
.B2(n_254),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_796),
.A2(n_389),
.B1(n_261),
.B2(n_240),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_900),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_790),
.B(n_618),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_844),
.B(n_239),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_887),
.A2(n_506),
.B(n_7),
.C(n_9),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_909),
.A2(n_520),
.B(n_534),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_844),
.B(n_240),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_917),
.B(n_661),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_814),
.A2(n_364),
.B(n_261),
.Y(n_1060)
);

BUFx12f_ASAP7_75t_L g1061 ( 
.A(n_892),
.Y(n_1061)
);

AO21x1_ASAP7_75t_L g1062 ( 
.A1(n_837),
.A2(n_661),
.B(n_225),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_825),
.A2(n_411),
.B1(n_364),
.B2(n_365),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_857),
.B(n_365),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_900),
.B(n_372),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_774),
.B(n_372),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_914),
.A2(n_520),
.B(n_534),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_910),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_910),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_919),
.A2(n_520),
.B(n_534),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_920),
.B(n_378),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_766),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_920),
.B(n_378),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_839),
.A2(n_661),
.B1(n_505),
.B2(n_385),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_921),
.B(n_382),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_807),
.B(n_661),
.Y(n_1076)
);

NOR2x2_ASAP7_75t_L g1077 ( 
.A(n_807),
.B(n_5),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_837),
.A2(n_382),
.B(n_385),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_883),
.A2(n_534),
.B(n_532),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_774),
.B(n_394),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_SL g1081 ( 
.A(n_891),
.B(n_922),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_922),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_921),
.B(n_394),
.Y(n_1083)
);

AO21x1_ASAP7_75t_L g1084 ( 
.A1(n_888),
.A2(n_279),
.B(n_519),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_889),
.A2(n_532),
.B(n_520),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_923),
.B(n_399),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_912),
.A2(n_9),
.B(n_11),
.C(n_13),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_896),
.A2(n_520),
.B(n_532),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_848),
.A2(n_399),
.B1(n_405),
.B2(n_408),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_911),
.B(n_405),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_863),
.B(n_408),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_904),
.A2(n_532),
.B(n_520),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_848),
.A2(n_409),
.B(n_326),
.C(n_358),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_874),
.A2(n_409),
.B1(n_268),
.B2(n_312),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_802),
.A2(n_520),
.B(n_334),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_806),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_852),
.A2(n_309),
.B(n_356),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_792),
.B(n_269),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_913),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_876),
.B(n_806),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_792),
.B(n_271),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_833),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_867),
.A2(n_336),
.B(n_354),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_912),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_SL g1105 ( 
.A(n_922),
.B(n_306),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_864),
.A2(n_278),
.B(n_353),
.C(n_281),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_806),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_916),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_806),
.B(n_339),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_948),
.A2(n_864),
.B(n_865),
.C(n_880),
.Y(n_1110)
);

AOI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1014),
.A2(n_838),
.B1(n_865),
.B2(n_880),
.C(n_873),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1027),
.A2(n_884),
.B1(n_898),
.B2(n_897),
.Y(n_1112)
);

AO21x1_ASAP7_75t_L g1113 ( 
.A1(n_996),
.A2(n_898),
.B(n_897),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_934),
.A2(n_855),
.B1(n_858),
.B2(n_884),
.Y(n_1114)
);

XOR2x2_ASAP7_75t_SL g1115 ( 
.A(n_944),
.B(n_18),
.Y(n_1115)
);

INVx6_ASAP7_75t_SL g1116 ( 
.A(n_990),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1001),
.B(n_847),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_972),
.B(n_850),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_SL g1119 ( 
.A1(n_952),
.A2(n_850),
.B(n_851),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_1003),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1105),
.B(n_858),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_951),
.B(n_851),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1028),
.B(n_879),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_938),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_949),
.B(n_879),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_930),
.A2(n_933),
.B(n_929),
.Y(n_1126)
);

BUFx12f_ASAP7_75t_L g1127 ( 
.A(n_1009),
.Y(n_1127)
);

OAI22x1_ASAP7_75t_L g1128 ( 
.A1(n_1033),
.A2(n_899),
.B1(n_893),
.B2(n_768),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_937),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1008),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_954),
.A2(n_855),
.B1(n_832),
.B2(n_783),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_965),
.Y(n_1132)
);

OAI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1081),
.A2(n_341),
.B1(n_285),
.B2(n_287),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_946),
.B(n_342),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1002),
.A2(n_789),
.B(n_890),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1007),
.B(n_22),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1007),
.B(n_22),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1004),
.A2(n_350),
.B(n_349),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1078),
.A2(n_23),
.B(n_24),
.C(n_27),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1045),
.A2(n_303),
.B1(n_298),
.B2(n_279),
.Y(n_1140)
);

OR2x6_ASAP7_75t_SL g1141 ( 
.A(n_1041),
.B(n_24),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_967),
.A2(n_945),
.B(n_959),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1053),
.B(n_27),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_990),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_982),
.B(n_31),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_1000),
.B(n_279),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1068),
.B(n_33),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_SL g1148 ( 
.A1(n_976),
.A2(n_34),
.B(n_37),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_990),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_925),
.B(n_1082),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_984),
.A2(n_37),
.B(n_39),
.C(n_41),
.Y(n_1151)
);

NAND2xp33_ASAP7_75t_SL g1152 ( 
.A(n_1000),
.B(n_279),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_932),
.A2(n_939),
.B(n_968),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_950),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_1021),
.B(n_100),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1069),
.B(n_39),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_971),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1061),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_977),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1018),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_932),
.A2(n_107),
.B(n_193),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_986),
.B(n_46),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_978),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_993),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1086),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1034),
.A2(n_1104),
.B(n_1087),
.C(n_1056),
.Y(n_1166)
);

BUFx5_ASAP7_75t_L g1167 ( 
.A(n_1099),
.Y(n_1167)
);

OAI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_1089),
.A2(n_1063),
.B(n_1020),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1059),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_994),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_926),
.B(n_52),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1018),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_939),
.A2(n_968),
.B(n_941),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_986),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_995),
.B(n_52),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1037),
.Y(n_1176)
);

OAI21xp33_ASAP7_75t_L g1177 ( 
.A1(n_1055),
.A2(n_1064),
.B(n_1058),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1066),
.B(n_53),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_964),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1012),
.B(n_55),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1080),
.B(n_56),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1016),
.B(n_57),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_936),
.A2(n_150),
.B(n_187),
.Y(n_1183)
);

NOR2x1_ASAP7_75t_R g1184 ( 
.A(n_1077),
.B(n_519),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1036),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_942),
.A2(n_57),
.B(n_59),
.C(n_61),
.Y(n_1186)
);

OR2x6_ASAP7_75t_L g1187 ( 
.A(n_958),
.B(n_1076),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1108),
.A2(n_519),
.B1(n_61),
.B2(n_94),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1018),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1043),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1093),
.A2(n_519),
.B(n_97),
.C(n_106),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1017),
.A2(n_79),
.B(n_108),
.C(n_125),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_963),
.A2(n_139),
.B1(n_142),
.B2(n_151),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_928),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1019),
.B(n_998),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_958),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1011),
.A2(n_163),
.B1(n_164),
.B2(n_167),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1090),
.B(n_1029),
.Y(n_1198)
);

INVx4_ASAP7_75t_L g1199 ( 
.A(n_1019),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1024),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_974),
.A2(n_171),
.B(n_179),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_958),
.Y(n_1202)
);

XNOR2xp5_ASAP7_75t_L g1203 ( 
.A(n_992),
.B(n_182),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1048),
.B(n_186),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_974),
.A2(n_973),
.B(n_983),
.C(n_1060),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_961),
.B(n_1023),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1024),
.B(n_1049),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_983),
.A2(n_1040),
.B(n_1026),
.C(n_1038),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1030),
.B(n_1031),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_960),
.A2(n_1046),
.B(n_1106),
.C(n_1075),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1098),
.B(n_1101),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_928),
.B(n_935),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1006),
.A2(n_1044),
.B(n_980),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1024),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1040),
.A2(n_1038),
.B(n_1035),
.C(n_1010),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_979),
.A2(n_987),
.B1(n_985),
.B2(n_955),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_1065),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_964),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1071),
.A2(n_1073),
.B(n_1083),
.C(n_1052),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1044),
.A2(n_927),
.B(n_962),
.Y(n_1220)
);

NAND3xp33_ASAP7_75t_SL g1221 ( 
.A(n_1103),
.B(n_1097),
.C(n_1051),
.Y(n_1221)
);

NOR3xp33_ASAP7_75t_SL g1222 ( 
.A(n_1103),
.B(n_1109),
.C(n_1032),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_966),
.B(n_969),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_935),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_991),
.A2(n_1097),
.B(n_988),
.C(n_1102),
.Y(n_1225)
);

NOR2x1_ASAP7_75t_L g1226 ( 
.A(n_1107),
.B(n_1091),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_931),
.Y(n_1227)
);

NAND3xp33_ASAP7_75t_SL g1228 ( 
.A(n_1094),
.B(n_1074),
.C(n_997),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_927),
.A2(n_962),
.B(n_956),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1102),
.A2(n_940),
.B(n_989),
.C(n_999),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_931),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_981),
.A2(n_1088),
.B(n_1079),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1079),
.A2(n_1088),
.B(n_1085),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1107),
.A2(n_1072),
.B1(n_1096),
.B2(n_1049),
.Y(n_1234)
);

INVx3_ASAP7_75t_SL g1235 ( 
.A(n_1049),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1072),
.B(n_1096),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1072),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_953),
.A2(n_975),
.B(n_970),
.C(n_1100),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1022),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_956),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1085),
.A2(n_1092),
.B(n_947),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1096),
.B(n_989),
.Y(n_1242)
);

AO22x1_ASAP7_75t_L g1243 ( 
.A1(n_1005),
.A2(n_1054),
.B1(n_1047),
.B2(n_1039),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_SL g1244 ( 
.A(n_1025),
.B(n_999),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1015),
.B(n_1042),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_SL g1246 ( 
.A1(n_1095),
.A2(n_1042),
.B(n_1092),
.C(n_1015),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_957),
.B(n_1050),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1062),
.A2(n_1095),
.B1(n_1084),
.B2(n_1050),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_943),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1057),
.A2(n_1067),
.B(n_1070),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1057),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1067),
.A2(n_1070),
.B(n_1013),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1013),
.A2(n_769),
.B1(n_878),
.B2(n_704),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1014),
.A2(n_769),
.B1(n_878),
.B2(n_704),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1008),
.Y(n_1255)
);

AND2x4_ASAP7_75t_SL g1256 ( 
.A(n_1007),
.B(n_812),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_951),
.B(n_878),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_938),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_948),
.B(n_769),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1008),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_951),
.A2(n_1014),
.B1(n_906),
.B2(n_871),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_951),
.B(n_878),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1027),
.A2(n_608),
.B(n_617),
.C(n_614),
.Y(n_1263)
);

AOI22x1_ASAP7_75t_L g1264 ( 
.A1(n_983),
.A2(n_974),
.B1(n_968),
.B2(n_989),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_1205),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1263),
.A2(n_1153),
.B(n_1250),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1245),
.A2(n_1173),
.B(n_1220),
.Y(n_1267)
);

BUFx4f_ASAP7_75t_SL g1268 ( 
.A(n_1127),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1212),
.B(n_1194),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1224),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1168),
.A2(n_1181),
.B(n_1254),
.C(n_1198),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1245),
.A2(n_1213),
.B(n_1216),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1253),
.A2(n_1211),
.B1(n_1112),
.B2(n_1261),
.Y(n_1273)
);

AO21x1_ASAP7_75t_L g1274 ( 
.A1(n_1171),
.A2(n_1139),
.B(n_1157),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1262),
.B(n_1165),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1232),
.A2(n_1252),
.B(n_1233),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1165),
.A2(n_1178),
.B1(n_1145),
.B2(n_1162),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1129),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1264),
.A2(n_1229),
.B(n_1241),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1122),
.B(n_1217),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1235),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1124),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1149),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1247),
.A2(n_1135),
.B(n_1240),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1247),
.A2(n_1242),
.B(n_1161),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1132),
.Y(n_1286)
);

INVx4_ASAP7_75t_L g1287 ( 
.A(n_1120),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1242),
.A2(n_1201),
.B(n_1248),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1216),
.A2(n_1110),
.B(n_1246),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1119),
.A2(n_1183),
.B(n_1239),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1177),
.A2(n_1219),
.B(n_1111),
.C(n_1166),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1209),
.B(n_1174),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1151),
.A2(n_1182),
.B(n_1134),
.C(n_1170),
.Y(n_1293)
);

BUFx10_ASAP7_75t_L g1294 ( 
.A(n_1136),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1163),
.A2(n_1170),
.B(n_1195),
.C(n_1180),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1230),
.A2(n_1225),
.A3(n_1128),
.B(n_1208),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1114),
.A2(n_1228),
.B1(n_1190),
.B2(n_1260),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1152),
.A2(n_1146),
.B(n_1210),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1206),
.A2(n_1186),
.B(n_1121),
.C(n_1155),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1159),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1251),
.A2(n_1238),
.B(n_1234),
.Y(n_1301)
);

BUFx4f_ASAP7_75t_L g1302 ( 
.A(n_1256),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1163),
.A2(n_1148),
.B1(n_1175),
.B2(n_1138),
.C(n_1143),
.Y(n_1303)
);

AND2x6_ASAP7_75t_L g1304 ( 
.A(n_1162),
.B(n_1136),
.Y(n_1304)
);

AO21x1_ASAP7_75t_L g1305 ( 
.A1(n_1197),
.A2(n_1244),
.B(n_1193),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1191),
.A2(n_1221),
.B(n_1175),
.C(n_1215),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_SL g1307 ( 
.A1(n_1192),
.A2(n_1147),
.B(n_1143),
.C(n_1156),
.Y(n_1307)
);

INVx3_ASAP7_75t_SL g1308 ( 
.A(n_1120),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1154),
.Y(n_1309)
);

BUFx8_ASAP7_75t_L g1310 ( 
.A(n_1158),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1118),
.A2(n_1144),
.B1(n_1116),
.B2(n_1137),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1146),
.A2(n_1117),
.B(n_1123),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1164),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1258),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1123),
.A2(n_1243),
.B(n_1114),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1234),
.A2(n_1125),
.B(n_1131),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1176),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1255),
.A2(n_1197),
.A3(n_1193),
.B(n_1156),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1223),
.A2(n_1222),
.B(n_1147),
.C(n_1150),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1169),
.B(n_1137),
.Y(n_1320)
);

NAND2xp33_ASAP7_75t_L g1321 ( 
.A(n_1160),
.B(n_1189),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1236),
.A2(n_1199),
.B(n_1204),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1236),
.A2(n_1199),
.B(n_1207),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1144),
.B(n_1141),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1160),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1179),
.A2(n_1218),
.B(n_1249),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1167),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1185),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1179),
.A2(n_1218),
.B(n_1214),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1116),
.A2(n_1140),
.B1(n_1133),
.B2(n_1188),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1226),
.A2(n_1237),
.B(n_1202),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1214),
.A2(n_1237),
.B(n_1160),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1167),
.A2(n_1203),
.B(n_1200),
.Y(n_1333)
);

A2O1A1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1115),
.A2(n_1196),
.B(n_1172),
.C(n_1189),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1187),
.A2(n_1200),
.B1(n_1172),
.B2(n_1189),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1172),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1167),
.B(n_1184),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1167),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1187),
.B(n_1167),
.Y(n_1339)
);

AO32x2_ASAP7_75t_L g1340 ( 
.A1(n_1187),
.A2(n_1170),
.A3(n_1163),
.B1(n_1216),
.B2(n_952),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1259),
.B(n_878),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1212),
.B(n_1194),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_R g1343 ( 
.A(n_1127),
.B(n_1003),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1113),
.A2(n_1227),
.A3(n_1231),
.B(n_1084),
.Y(n_1344)
);

OAI22x1_ASAP7_75t_L g1345 ( 
.A1(n_1254),
.A2(n_1171),
.B1(n_1181),
.B2(n_1198),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1254),
.A2(n_769),
.B(n_1181),
.Y(n_1346)
);

AOI221xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1168),
.A2(n_1263),
.B1(n_1151),
.B2(n_615),
.C(n_1181),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1259),
.B(n_878),
.Y(n_1348)
);

AO32x2_ASAP7_75t_L g1349 ( 
.A1(n_1163),
.A2(n_1170),
.A3(n_1216),
.B1(n_952),
.B2(n_1114),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1113),
.A2(n_1227),
.A3(n_1231),
.B(n_1084),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1259),
.B(n_1254),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1232),
.A2(n_1252),
.B(n_1233),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1259),
.B(n_1254),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1129),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1168),
.A2(n_1263),
.B1(n_1151),
.B2(n_615),
.C(n_1181),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_933),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_L g1357 ( 
.A(n_1212),
.B(n_1009),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1127),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1116),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_1129),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_SL g1361 ( 
.A1(n_1263),
.A2(n_1259),
.B(n_1166),
.C(n_1205),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_933),
.Y(n_1362)
);

INVxp33_ASAP7_75t_L g1363 ( 
.A(n_1129),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1181),
.A2(n_1198),
.B1(n_1171),
.B2(n_1254),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1259),
.B(n_878),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1263),
.A2(n_1259),
.B(n_1168),
.C(n_1181),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1113),
.A2(n_1227),
.A3(n_1231),
.B(n_1084),
.Y(n_1367)
);

AOI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1254),
.A2(n_769),
.B(n_755),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1224),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_SL g1370 ( 
.A1(n_1210),
.A2(n_1238),
.B(n_952),
.Y(n_1370)
);

O2A1O1Ixp5_ASAP7_75t_L g1371 ( 
.A1(n_1181),
.A2(n_1173),
.B(n_1205),
.C(n_1198),
.Y(n_1371)
);

NAND3xp33_ASAP7_75t_SL g1372 ( 
.A(n_1254),
.B(n_769),
.C(n_1181),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1248),
.A2(n_1231),
.B(n_1227),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1259),
.B(n_878),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1194),
.B(n_928),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1124),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1254),
.B(n_769),
.C(n_1181),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_933),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1127),
.Y(n_1379)
);

AO21x1_ASAP7_75t_L g1380 ( 
.A1(n_1171),
.A2(n_1263),
.B(n_1181),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1259),
.B(n_878),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1232),
.A2(n_1252),
.B(n_1233),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1181),
.A2(n_1198),
.B1(n_1171),
.B2(n_1254),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1110),
.A2(n_952),
.B(n_866),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1224),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_933),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1259),
.B(n_1254),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1263),
.A2(n_769),
.B(n_1254),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1212),
.B(n_1194),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1263),
.A2(n_1259),
.B(n_1168),
.C(n_1181),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1113),
.A2(n_1227),
.A3(n_1231),
.B(n_1084),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1120),
.B(n_812),
.Y(n_1392)
);

OAI21xp33_ASAP7_75t_L g1393 ( 
.A1(n_1168),
.A2(n_769),
.B(n_1254),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1232),
.A2(n_1252),
.B(n_1233),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1259),
.B(n_1198),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1263),
.A2(n_1259),
.B(n_1168),
.C(n_1181),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1136),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1248),
.A2(n_1231),
.B(n_1227),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1124),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1263),
.A2(n_769),
.B(n_1254),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1224),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_933),
.Y(n_1402)
);

OAI21xp33_ASAP7_75t_L g1403 ( 
.A1(n_1168),
.A2(n_769),
.B(n_1254),
.Y(n_1403)
);

AO32x2_ASAP7_75t_L g1404 ( 
.A1(n_1163),
.A2(n_1170),
.A3(n_1216),
.B1(n_952),
.B2(n_1114),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1254),
.B(n_769),
.C(n_1181),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1232),
.A2(n_1252),
.B(n_1233),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1153),
.A2(n_1250),
.B(n_1220),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1200),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1126),
.A2(n_1142),
.B(n_933),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1259),
.B(n_1254),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1153),
.A2(n_1250),
.B(n_1220),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1254),
.B(n_769),
.C(n_1181),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1259),
.B(n_878),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1259),
.B(n_1198),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1113),
.A2(n_1227),
.A3(n_1231),
.B(n_1084),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1130),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1227),
.Y(n_1417)
);

AO31x2_ASAP7_75t_L g1418 ( 
.A1(n_1113),
.A2(n_1227),
.A3(n_1231),
.B(n_1084),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1129),
.B(n_1257),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1200),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1259),
.B(n_878),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1302),
.B(n_1337),
.Y(n_1422)
);

CKINVDCx11_ASAP7_75t_R g1423 ( 
.A(n_1270),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1369),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1345),
.A2(n_1383),
.B1(n_1364),
.B2(n_1380),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1273),
.A2(n_1372),
.B1(n_1377),
.B2(n_1412),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1281),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1405),
.A2(n_1304),
.B1(n_1388),
.B2(n_1400),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1304),
.A2(n_1414),
.B1(n_1395),
.B2(n_1370),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1282),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1304),
.Y(n_1431)
);

INVx6_ASAP7_75t_L g1432 ( 
.A(n_1281),
.Y(n_1432)
);

BUFx2_ASAP7_75t_SL g1433 ( 
.A(n_1385),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1346),
.A2(n_1351),
.B1(n_1410),
.B2(n_1387),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1271),
.A2(n_1403),
.B1(n_1393),
.B2(n_1355),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1341),
.B(n_1348),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1286),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1353),
.A2(n_1274),
.B1(n_1368),
.B2(n_1381),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1401),
.Y(n_1439)
);

INVx11_ASAP7_75t_L g1440 ( 
.A(n_1310),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1300),
.Y(n_1441)
);

CKINVDCx6p67_ASAP7_75t_R g1442 ( 
.A(n_1308),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1304),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1305),
.A2(n_1272),
.B(n_1356),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1365),
.A2(n_1421),
.B1(n_1413),
.B2(n_1374),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1310),
.Y(n_1446)
);

CKINVDCx11_ASAP7_75t_R g1447 ( 
.A(n_1309),
.Y(n_1447)
);

BUFx10_ASAP7_75t_L g1448 ( 
.A(n_1358),
.Y(n_1448)
);

BUFx12f_ASAP7_75t_L g1449 ( 
.A(n_1294),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1366),
.A2(n_1390),
.B1(n_1396),
.B2(n_1291),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1268),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1313),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1324),
.A2(n_1330),
.B1(n_1340),
.B2(n_1404),
.Y(n_1453)
);

CKINVDCx11_ASAP7_75t_R g1454 ( 
.A(n_1379),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1397),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1314),
.Y(n_1456)
);

INVx3_ASAP7_75t_SL g1457 ( 
.A(n_1287),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1362),
.A2(n_1378),
.B(n_1386),
.Y(n_1458)
);

CKINVDCx11_ASAP7_75t_R g1459 ( 
.A(n_1328),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1277),
.A2(n_1295),
.B1(n_1293),
.B2(n_1299),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1347),
.A2(n_1311),
.B1(n_1334),
.B2(n_1320),
.Y(n_1461)
);

CKINVDCx11_ASAP7_75t_R g1462 ( 
.A(n_1397),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1306),
.A2(n_1360),
.B1(n_1278),
.B2(n_1384),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1292),
.B(n_1280),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1416),
.A2(n_1297),
.B1(n_1419),
.B2(n_1317),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1354),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1284),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1363),
.B(n_1269),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1376),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1357),
.A2(n_1289),
.B1(n_1298),
.B2(n_1319),
.Y(n_1470)
);

NAND2x1p5_ASAP7_75t_L g1471 ( 
.A(n_1342),
.B(n_1389),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1287),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1339),
.A2(n_1315),
.B1(n_1265),
.B2(n_1283),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1392),
.A2(n_1404),
.B1(n_1349),
.B2(n_1340),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1339),
.A2(n_1392),
.B1(n_1266),
.B2(n_1375),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1389),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1408),
.B(n_1420),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1359),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1325),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1303),
.A2(n_1361),
.B1(n_1335),
.B2(n_1399),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1349),
.A2(n_1404),
.B1(n_1340),
.B2(n_1417),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1349),
.A2(n_1417),
.B1(n_1312),
.B2(n_1333),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1307),
.A2(n_1338),
.B1(n_1327),
.B2(n_1321),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1336),
.B(n_1420),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1343),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1327),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1316),
.A2(n_1301),
.B1(n_1371),
.B2(n_1290),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1318),
.A2(n_1402),
.B1(n_1409),
.B2(n_1288),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1373),
.A2(n_1398),
.B1(n_1338),
.B2(n_1331),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1408),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1329),
.A2(n_1332),
.B1(n_1322),
.B2(n_1323),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1326),
.A2(n_1285),
.B1(n_1267),
.B2(n_1318),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1296),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1407),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1318),
.A2(n_1296),
.B1(n_1411),
.B2(n_1407),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_SL g1496 ( 
.A(n_1296),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1411),
.A2(n_1279),
.B1(n_1276),
.B2(n_1406),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1344),
.A2(n_1350),
.B1(n_1415),
.B2(n_1391),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1352),
.A2(n_1382),
.B1(n_1394),
.B2(n_1367),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1418),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1391),
.A2(n_1273),
.B1(n_1383),
.B2(n_1364),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1391),
.A2(n_1415),
.B1(n_1418),
.B2(n_1364),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1273),
.A2(n_1383),
.B1(n_1364),
.B2(n_1393),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1281),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1273),
.A2(n_1383),
.B1(n_1364),
.B2(n_1393),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1273),
.A2(n_1383),
.B1(n_1364),
.B2(n_1393),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1282),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1358),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1304),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1273),
.A2(n_1377),
.B1(n_1412),
.B2(n_1405),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1273),
.A2(n_1377),
.B1(n_1412),
.B2(n_1405),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1364),
.A2(n_1383),
.B1(n_1405),
.B2(n_1377),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1270),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1270),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1273),
.A2(n_1377),
.B1(n_1412),
.B2(n_1405),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1310),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1345),
.A2(n_1383),
.B1(n_1364),
.B2(n_1380),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1419),
.B(n_1275),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1282),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1272),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1364),
.A2(n_1383),
.B1(n_1405),
.B2(n_1377),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1345),
.A2(n_1383),
.B1(n_1364),
.B2(n_1380),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1345),
.A2(n_1383),
.B1(n_1364),
.B2(n_1380),
.Y(n_1523)
);

OAI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1364),
.A2(n_1383),
.B1(n_1346),
.B2(n_1377),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_SL g1525 ( 
.A1(n_1346),
.A2(n_1383),
.B(n_1364),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1305),
.A2(n_1272),
.B(n_1356),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1364),
.A2(n_1383),
.B1(n_1405),
.B2(n_1377),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1273),
.A2(n_1377),
.B1(n_1412),
.B2(n_1405),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1364),
.A2(n_1383),
.B1(n_1405),
.B2(n_1377),
.Y(n_1529)
);

INVx6_ASAP7_75t_L g1530 ( 
.A(n_1281),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1364),
.A2(n_1383),
.B1(n_1405),
.B2(n_1377),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1281),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1345),
.A2(n_1383),
.B1(n_1364),
.B2(n_1380),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1310),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1395),
.B(n_1414),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1281),
.Y(n_1536)
);

BUFx12f_ASAP7_75t_L g1537 ( 
.A(n_1310),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1273),
.A2(n_1377),
.B1(n_1412),
.B2(n_1405),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1310),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_1272),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1270),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1282),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1273),
.A2(n_1377),
.B1(n_1412),
.B2(n_1405),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1273),
.A2(n_1377),
.B1(n_1412),
.B2(n_1405),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1345),
.A2(n_1383),
.B1(n_1364),
.B2(n_1380),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1364),
.A2(n_1383),
.B1(n_1414),
.B2(n_1395),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1345),
.A2(n_1383),
.B1(n_1364),
.B2(n_1380),
.Y(n_1547)
);

OAI21xp33_ASAP7_75t_L g1548 ( 
.A1(n_1364),
.A2(n_1383),
.B(n_1346),
.Y(n_1548)
);

CKINVDCx6p67_ASAP7_75t_R g1549 ( 
.A(n_1308),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1281),
.Y(n_1550)
);

CKINVDCx6p67_ASAP7_75t_R g1551 ( 
.A(n_1308),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1444),
.A2(n_1526),
.B(n_1458),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1466),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1503),
.A2(n_1506),
.B1(n_1505),
.B2(n_1546),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1494),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1493),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1481),
.B(n_1453),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1430),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1437),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1459),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1441),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1481),
.B(n_1453),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1452),
.B(n_1456),
.Y(n_1563)
);

NOR2x1_ASAP7_75t_L g1564 ( 
.A(n_1470),
.B(n_1473),
.Y(n_1564)
);

BUFx4f_ASAP7_75t_SL g1565 ( 
.A(n_1516),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1469),
.B(n_1507),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1519),
.B(n_1542),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1432),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1518),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1502),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1496),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1486),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1500),
.Y(n_1573)
);

BUFx2_ASAP7_75t_SL g1574 ( 
.A(n_1443),
.Y(n_1574)
);

NAND2x1p5_ASAP7_75t_L g1575 ( 
.A(n_1443),
.B(n_1431),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1535),
.B(n_1464),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1467),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1467),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1423),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1463),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1474),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1501),
.B(n_1482),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1424),
.B(n_1541),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1474),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_L g1585 ( 
.A(n_1525),
.B(n_1515),
.C(n_1510),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1520),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1501),
.B(n_1512),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1509),
.B(n_1475),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1520),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1540),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1540),
.Y(n_1591)
);

OA21x2_ASAP7_75t_L g1592 ( 
.A1(n_1444),
.A2(n_1526),
.B(n_1458),
.Y(n_1592)
);

AO21x2_ASAP7_75t_L g1593 ( 
.A1(n_1495),
.A2(n_1435),
.B(n_1434),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1548),
.A2(n_1510),
.B1(n_1528),
.B2(n_1538),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1482),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1498),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1491),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1514),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1428),
.B(n_1511),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1432),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1498),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1495),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1489),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1489),
.Y(n_1604)
);

CKINVDCx6p67_ASAP7_75t_R g1605 ( 
.A(n_1485),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1521),
.B(n_1527),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1483),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1428),
.B(n_1511),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1480),
.Y(n_1609)
);

AOI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1450),
.A2(n_1460),
.B(n_1531),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1513),
.B(n_1439),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1515),
.B(n_1528),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1529),
.B(n_1503),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1538),
.B(n_1543),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1488),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1543),
.B(n_1544),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1488),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1492),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1544),
.B(n_1505),
.Y(n_1619)
);

AO21x1_ASAP7_75t_SL g1620 ( 
.A1(n_1506),
.A2(n_1522),
.B(n_1425),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1479),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1477),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1426),
.B(n_1434),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1468),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1497),
.A2(n_1499),
.B(n_1438),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_SL g1626 ( 
.A1(n_1517),
.A2(n_1533),
.B(n_1523),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1524),
.B(n_1547),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1524),
.B(n_1436),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_1454),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1487),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1484),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1487),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1465),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1461),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1490),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1545),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1429),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1432),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1445),
.B(n_1532),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1445),
.B(n_1532),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1550),
.B(n_1471),
.Y(n_1641)
);

OAI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1422),
.A2(n_1476),
.B1(n_1449),
.B2(n_1537),
.Y(n_1642)
);

OA21x2_ASAP7_75t_L g1643 ( 
.A1(n_1427),
.A2(n_1455),
.B(n_1530),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1504),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1622),
.B(n_1536),
.Y(n_1645)
);

INVx5_ASAP7_75t_SL g1646 ( 
.A(n_1605),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1569),
.B(n_1433),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1563),
.B(n_1530),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1585),
.A2(n_1446),
.B(n_1508),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_L g1650 ( 
.A1(n_1612),
.A2(n_1451),
.B(n_1447),
.C(n_1462),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1621),
.B(n_1472),
.Y(n_1651)
);

O2A1O1Ixp33_ASAP7_75t_SL g1652 ( 
.A1(n_1606),
.A2(n_1623),
.B(n_1554),
.C(n_1613),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1597),
.B(n_1504),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1561),
.B(n_1551),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1606),
.B(n_1457),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_SL g1656 ( 
.A1(n_1610),
.A2(n_1440),
.B(n_1539),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1553),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1594),
.A2(n_1442),
.B(n_1549),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1588),
.B(n_1478),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1612),
.A2(n_1614),
.B(n_1616),
.C(n_1599),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1614),
.A2(n_1448),
.B(n_1534),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1558),
.Y(n_1662)
);

BUFx12f_ASAP7_75t_L g1663 ( 
.A(n_1579),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1599),
.A2(n_1448),
.B1(n_1608),
.B2(n_1616),
.Y(n_1664)
);

A2O1A1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1608),
.A2(n_1623),
.B(n_1627),
.C(n_1619),
.Y(n_1665)
);

NAND2xp33_ASAP7_75t_SL g1666 ( 
.A(n_1629),
.B(n_1619),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1588),
.B(n_1571),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1627),
.A2(n_1613),
.B1(n_1636),
.B2(n_1587),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1605),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1566),
.B(n_1567),
.Y(n_1670)
);

CKINVDCx16_ASAP7_75t_R g1671 ( 
.A(n_1572),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1566),
.B(n_1567),
.Y(n_1673)
);

A2O1A1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1587),
.A2(n_1564),
.B(n_1580),
.C(n_1628),
.Y(n_1674)
);

BUFx2_ASAP7_75t_SL g1675 ( 
.A(n_1572),
.Y(n_1675)
);

O2A1O1Ixp33_ASAP7_75t_SL g1676 ( 
.A1(n_1560),
.A2(n_1642),
.B(n_1635),
.C(n_1611),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1590),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1598),
.Y(n_1678)
);

NOR2x1_ASAP7_75t_SL g1679 ( 
.A(n_1593),
.B(n_1572),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1565),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1631),
.B(n_1624),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1644),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1634),
.A2(n_1593),
.B1(n_1637),
.B2(n_1582),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1576),
.B(n_1583),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1620),
.A2(n_1626),
.B1(n_1562),
.B2(n_1557),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1610),
.B(n_1609),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1609),
.A2(n_1607),
.B(n_1552),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1570),
.B(n_1586),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1625),
.A2(n_1632),
.B(n_1630),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1639),
.B(n_1641),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1577),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1556),
.B(n_1573),
.Y(n_1692)
);

AO32x2_ASAP7_75t_L g1693 ( 
.A1(n_1568),
.A2(n_1638),
.A3(n_1600),
.B1(n_1584),
.B2(n_1581),
.Y(n_1693)
);

A2O1A1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1615),
.A2(n_1617),
.B(n_1630),
.C(n_1632),
.Y(n_1694)
);

OR2x6_ASAP7_75t_L g1695 ( 
.A(n_1574),
.B(n_1643),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1602),
.A2(n_1618),
.B(n_1607),
.C(n_1595),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1603),
.A2(n_1604),
.B(n_1591),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1574),
.B(n_1575),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1670),
.B(n_1592),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1673),
.B(n_1592),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1662),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1687),
.B(n_1592),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1687),
.B(n_1693),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1688),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1688),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1659),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1659),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1693),
.B(n_1586),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1672),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1695),
.B(n_1555),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1686),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1686),
.B(n_1589),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1697),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1691),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1677),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1691),
.B(n_1589),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1693),
.B(n_1591),
.Y(n_1717)
);

INVxp33_ASAP7_75t_L g1718 ( 
.A(n_1655),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1692),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1657),
.B(n_1578),
.Y(n_1720)
);

NOR2xp67_ASAP7_75t_L g1721 ( 
.A(n_1653),
.B(n_1578),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1692),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1683),
.B(n_1681),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1682),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1685),
.A2(n_1620),
.B1(n_1626),
.B2(n_1633),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1698),
.Y(n_1726)
);

OAI31xp33_ASAP7_75t_L g1727 ( 
.A1(n_1703),
.A2(n_1660),
.A3(n_1665),
.B(n_1674),
.Y(n_1727)
);

AND2x2_ASAP7_75t_SL g1728 ( 
.A(n_1703),
.B(n_1685),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1716),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1720),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1707),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1710),
.B(n_1679),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1704),
.B(n_1689),
.Y(n_1733)
);

INVx2_ASAP7_75t_R g1734 ( 
.A(n_1702),
.Y(n_1734)
);

OA21x2_ASAP7_75t_L g1735 ( 
.A1(n_1713),
.A2(n_1694),
.B(n_1696),
.Y(n_1735)
);

NAND4xp25_ASAP7_75t_L g1736 ( 
.A(n_1702),
.B(n_1649),
.C(n_1655),
.D(n_1652),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1695),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1713),
.Y(n_1738)
);

AO211x2_ASAP7_75t_L g1739 ( 
.A1(n_1723),
.A2(n_1649),
.B(n_1658),
.C(n_1661),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1714),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1714),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1699),
.B(n_1648),
.Y(n_1742)
);

OAI33xp33_ASAP7_75t_L g1743 ( 
.A1(n_1711),
.A2(n_1601),
.A3(n_1596),
.B1(n_1647),
.B2(n_1654),
.B3(n_1640),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1724),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1700),
.B(n_1690),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1724),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1707),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_SL g1748 ( 
.A(n_1726),
.B(n_1671),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1704),
.B(n_1668),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1711),
.B(n_1668),
.C(n_1664),
.Y(n_1750)
);

INVx4_ASAP7_75t_L g1751 ( 
.A(n_1707),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1700),
.B(n_1708),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1718),
.B(n_1651),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1721),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1703),
.A2(n_1658),
.B1(n_1584),
.B2(n_1581),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1704),
.B(n_1684),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1701),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1708),
.B(n_1717),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1710),
.B(n_1667),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1712),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1705),
.B(n_1645),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1717),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1731),
.Y(n_1763)
);

CKINVDCx16_ASAP7_75t_R g1764 ( 
.A(n_1748),
.Y(n_1764)
);

OR2x6_ASAP7_75t_SL g1765 ( 
.A(n_1750),
.B(n_1723),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1734),
.B(n_1758),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1734),
.B(n_1719),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1732),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1734),
.B(n_1719),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1760),
.B(n_1705),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1758),
.B(n_1722),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1760),
.B(n_1705),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1744),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1757),
.Y(n_1774)
);

INVx4_ASAP7_75t_L g1775 ( 
.A(n_1751),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1758),
.B(n_1722),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1747),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1756),
.B(n_1718),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1752),
.B(n_1702),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1757),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1729),
.B(n_1712),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1729),
.B(n_1709),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1762),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1752),
.B(n_1715),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1746),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1747),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1738),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1762),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1741),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1741),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1740),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1745),
.B(n_1706),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1745),
.B(n_1706),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1749),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1745),
.B(n_1751),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1749),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1730),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1765),
.A2(n_1728),
.B1(n_1750),
.B2(n_1755),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1792),
.B(n_1751),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1781),
.B(n_1756),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1777),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1766),
.B(n_1737),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1778),
.B(n_1728),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1792),
.B(n_1793),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1774),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1781),
.B(n_1730),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1766),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1774),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1770),
.B(n_1761),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1763),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1774),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1763),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1780),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1770),
.B(n_1761),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1772),
.B(n_1733),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1766),
.B(n_1759),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1780),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1778),
.B(n_1728),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1772),
.B(n_1733),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1794),
.B(n_1754),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1771),
.B(n_1759),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1771),
.B(n_1742),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1782),
.B(n_1720),
.Y(n_1823)
);

A2O1A1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1765),
.A2(n_1727),
.B(n_1736),
.C(n_1755),
.Y(n_1824)
);

INVx2_ASAP7_75t_SL g1825 ( 
.A(n_1777),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1780),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1771),
.Y(n_1827)
);

OR2x6_ASAP7_75t_L g1828 ( 
.A(n_1794),
.B(n_1675),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1789),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1776),
.B(n_1764),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1789),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1789),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1790),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1790),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1790),
.Y(n_1835)
);

OAI211xp5_ASAP7_75t_L g1836 ( 
.A1(n_1775),
.A2(n_1736),
.B(n_1727),
.C(n_1664),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1776),
.B(n_1742),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1776),
.B(n_1742),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1791),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1791),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1830),
.B(n_1822),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1800),
.B(n_1783),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1807),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1800),
.B(n_1783),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1830),
.B(n_1795),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1824),
.B(n_1764),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1817),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1807),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1822),
.B(n_1795),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1812),
.B(n_1669),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1837),
.B(n_1795),
.Y(n_1851)
);

OAI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1798),
.A2(n_1836),
.B(n_1818),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1807),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1810),
.B(n_1765),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1810),
.Y(n_1855)
);

INVx1_ASAP7_75t_SL g1856 ( 
.A(n_1801),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1803),
.B(n_1764),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1820),
.B(n_1680),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1817),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1828),
.A2(n_1796),
.B(n_1765),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1827),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1839),
.B(n_1796),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1840),
.B(n_1797),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1801),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1835),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1835),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1827),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1809),
.B(n_1783),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1805),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1809),
.B(n_1788),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1825),
.B(n_1797),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1808),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1811),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1837),
.B(n_1784),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1828),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_SL g1876 ( 
.A1(n_1825),
.A2(n_1650),
.B(n_1786),
.Y(n_1876)
);

OR2x6_ASAP7_75t_L g1877 ( 
.A(n_1828),
.B(n_1656),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1854),
.Y(n_1878)
);

OAI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1860),
.A2(n_1735),
.B1(n_1828),
.B2(n_1748),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1842),
.B(n_1814),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1847),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1847),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1841),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1850),
.B(n_1663),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1841),
.B(n_1838),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1855),
.Y(n_1886)
);

OAI32xp33_ASAP7_75t_L g1887 ( 
.A1(n_1846),
.A2(n_1806),
.A3(n_1819),
.B1(n_1815),
.B2(n_1788),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1842),
.B(n_1814),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1855),
.B(n_1646),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1852),
.B(n_1775),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1857),
.A2(n_1739),
.B1(n_1743),
.B2(n_1735),
.Y(n_1891)
);

A2O1A1Ixp33_ASAP7_75t_L g1892 ( 
.A1(n_1876),
.A2(n_1666),
.B(n_1661),
.C(n_1739),
.Y(n_1892)
);

NAND2xp67_ASAP7_75t_SL g1893 ( 
.A(n_1845),
.B(n_1799),
.Y(n_1893)
);

OAI221xp5_ASAP7_75t_SL g1894 ( 
.A1(n_1876),
.A2(n_1815),
.B1(n_1819),
.B2(n_1806),
.C(n_1739),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1859),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1875),
.A2(n_1802),
.B1(n_1768),
.B2(n_1821),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1845),
.B(n_1838),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1859),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_1864),
.Y(n_1899)
);

OAI21xp33_ASAP7_75t_L g1900 ( 
.A1(n_1862),
.A2(n_1799),
.B(n_1804),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1865),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1865),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1844),
.B(n_1823),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1858),
.A2(n_1743),
.B1(n_1735),
.B2(n_1725),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1892),
.A2(n_1871),
.B(n_1863),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1880),
.B(n_1844),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1892),
.A2(n_1802),
.B1(n_1768),
.B2(n_1874),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1885),
.B(n_1874),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1883),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1899),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1883),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1886),
.B(n_1856),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1904),
.A2(n_1735),
.B1(n_1867),
.B2(n_1861),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1885),
.B(n_1849),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1897),
.B(n_1849),
.Y(n_1915)
);

OAI21xp33_ASAP7_75t_SL g1916 ( 
.A1(n_1890),
.A2(n_1851),
.B(n_1848),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_1878),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1894),
.B(n_1678),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1897),
.B(n_1851),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1880),
.B(n_1888),
.Y(n_1920)
);

OAI332xp33_ASAP7_75t_L g1921 ( 
.A1(n_1890),
.A2(n_1843),
.A3(n_1848),
.B1(n_1853),
.B2(n_1870),
.B3(n_1868),
.C1(n_1867),
.C2(n_1869),
.Y(n_1921)
);

OAI31xp33_ASAP7_75t_L g1922 ( 
.A1(n_1891),
.A2(n_1867),
.A3(n_1861),
.B(n_1868),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1888),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1903),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1881),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1924),
.Y(n_1926)
);

AOI21xp33_ASAP7_75t_L g1927 ( 
.A1(n_1917),
.A2(n_1887),
.B(n_1882),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1924),
.Y(n_1928)
);

INVx3_ASAP7_75t_L g1929 ( 
.A(n_1909),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1906),
.Y(n_1930)
);

INVx2_ASAP7_75t_SL g1931 ( 
.A(n_1909),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1908),
.B(n_1903),
.Y(n_1932)
);

XOR2x2_ASAP7_75t_L g1933 ( 
.A(n_1918),
.B(n_1884),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1906),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1908),
.B(n_1900),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1923),
.B(n_1889),
.Y(n_1936)
);

OAI21xp33_ASAP7_75t_SL g1937 ( 
.A1(n_1905),
.A2(n_1848),
.B(n_1843),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1910),
.B(n_1914),
.Y(n_1938)
);

NOR2x1_ASAP7_75t_L g1939 ( 
.A(n_1929),
.B(n_1912),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1929),
.Y(n_1940)
);

OAI21xp33_ASAP7_75t_L g1941 ( 
.A1(n_1932),
.A2(n_1918),
.B(n_1935),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1928),
.B(n_1920),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1936),
.B(n_1907),
.Y(n_1943)
);

AO22x2_ASAP7_75t_L g1944 ( 
.A1(n_1926),
.A2(n_1925),
.B1(n_1911),
.B2(n_1898),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_SL g1945 ( 
.A1(n_1927),
.A2(n_1922),
.B(n_1919),
.Y(n_1945)
);

NOR2xp67_ASAP7_75t_L g1946 ( 
.A(n_1930),
.B(n_1916),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1936),
.B(n_1921),
.Y(n_1947)
);

INVxp67_ASAP7_75t_L g1948 ( 
.A(n_1934),
.Y(n_1948)
);

AOI211xp5_ASAP7_75t_L g1949 ( 
.A1(n_1937),
.A2(n_1879),
.B(n_1896),
.C(n_1913),
.Y(n_1949)
);

AOI222xp33_ASAP7_75t_L g1950 ( 
.A1(n_1947),
.A2(n_1929),
.B1(n_1931),
.B2(n_1895),
.C1(n_1902),
.C2(n_1901),
.Y(n_1950)
);

AOI211x1_ASAP7_75t_L g1951 ( 
.A1(n_1943),
.A2(n_1941),
.B(n_1942),
.C(n_1938),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1944),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1939),
.B(n_1938),
.Y(n_1953)
);

OAI211xp5_ASAP7_75t_L g1954 ( 
.A1(n_1945),
.A2(n_1946),
.B(n_1949),
.C(n_1948),
.Y(n_1954)
);

O2A1O1Ixp5_ASAP7_75t_L g1955 ( 
.A1(n_1940),
.A2(n_1853),
.B(n_1843),
.C(n_1915),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_SL g1956 ( 
.A(n_1953),
.B(n_1931),
.Y(n_1956)
);

O2A1O1Ixp5_ASAP7_75t_L g1957 ( 
.A1(n_1954),
.A2(n_1853),
.B(n_1944),
.C(n_1866),
.Y(n_1957)
);

AO22x1_ASAP7_75t_L g1958 ( 
.A1(n_1952),
.A2(n_1933),
.B1(n_1869),
.B2(n_1873),
.Y(n_1958)
);

NOR4xp25_ASAP7_75t_L g1959 ( 
.A(n_1951),
.B(n_1933),
.C(n_1866),
.D(n_1873),
.Y(n_1959)
);

OAI221xp5_ASAP7_75t_L g1960 ( 
.A1(n_1950),
.A2(n_1877),
.B1(n_1870),
.B2(n_1872),
.C(n_1788),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1955),
.A2(n_1872),
.B(n_1877),
.Y(n_1961)
);

AOI211xp5_ASAP7_75t_L g1962 ( 
.A1(n_1954),
.A2(n_1802),
.B(n_1893),
.C(n_1676),
.Y(n_1962)
);

AO22x2_ASAP7_75t_L g1963 ( 
.A1(n_1959),
.A2(n_1831),
.B1(n_1834),
.B2(n_1833),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1956),
.B(n_1816),
.Y(n_1964)
);

XNOR2xp5_ASAP7_75t_L g1965 ( 
.A(n_1958),
.B(n_1877),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1957),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1961),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1960),
.Y(n_1968)
);

NOR3xp33_ASAP7_75t_L g1969 ( 
.A(n_1967),
.B(n_1962),
.C(n_1646),
.Y(n_1969)
);

NAND2x1p5_ASAP7_75t_L g1970 ( 
.A(n_1964),
.B(n_1646),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1966),
.B(n_1786),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1969),
.A2(n_1968),
.B1(n_1965),
.B2(n_1963),
.Y(n_1972)
);

AO22x2_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1971),
.B1(n_1963),
.B2(n_1970),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1973),
.A2(n_1877),
.B1(n_1768),
.B2(n_1829),
.Y(n_1974)
);

OAI22x1_ASAP7_75t_L g1975 ( 
.A1(n_1973),
.A2(n_1773),
.B1(n_1785),
.B2(n_1775),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1975),
.Y(n_1976)
);

AOI32xp33_ASAP7_75t_L g1977 ( 
.A1(n_1974),
.A2(n_1816),
.A3(n_1769),
.B1(n_1767),
.B2(n_1779),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_SL g1978 ( 
.A1(n_1976),
.A2(n_1877),
.B1(n_1832),
.B2(n_1777),
.Y(n_1978)
);

OAI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1977),
.A2(n_1826),
.B(n_1813),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_SL g1980 ( 
.A(n_1978),
.B(n_1775),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1979),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1981),
.B(n_1777),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1982),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1983),
.A2(n_1980),
.B1(n_1775),
.B2(n_1787),
.Y(n_1984)
);

AOI211xp5_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1753),
.B(n_1785),
.C(n_1773),
.Y(n_1985)
);


endmodule