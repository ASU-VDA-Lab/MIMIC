module real_aes_6672_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_182;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_L g437 ( .A1(n_0), .A2(n_7), .B1(n_438), .B2(n_709), .C1(n_714), .C2(n_715), .Y(n_437) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_1), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g431 ( .A(n_1), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_2), .A2(n_138), .B(n_143), .C(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_3), .A2(n_133), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g450 ( .A(n_4), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_5), .B(n_157), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_6), .B(n_434), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_7), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g467 ( .A1(n_8), .A2(n_133), .B(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g138 ( .A(n_9), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g167 ( .A(n_10), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_11), .B(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_11), .B(n_44), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_12), .A2(n_245), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_13), .B(n_148), .Y(n_184) );
INVx1_ASAP7_75t_L g472 ( .A(n_14), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_15), .B(n_147), .Y(n_520) );
INVx1_ASAP7_75t_L g131 ( .A(n_16), .Y(n_131) );
INVx1_ASAP7_75t_L g532 ( .A(n_17), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_18), .A2(n_168), .B(n_193), .C(n_195), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_19), .B(n_157), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_20), .B(n_461), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_21), .B(n_133), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_22), .B(n_253), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_23), .A2(n_147), .B(n_149), .C(n_153), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_24), .B(n_157), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_25), .B(n_148), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_26), .A2(n_151), .B(n_195), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_27), .B(n_148), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g213 ( .A(n_28), .Y(n_213) );
INVx1_ASAP7_75t_L g227 ( .A(n_29), .Y(n_227) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_30), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_31), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_32), .B(n_148), .Y(n_451) );
INVx1_ASAP7_75t_L g250 ( .A(n_33), .Y(n_250) );
INVx1_ASAP7_75t_L g485 ( .A(n_34), .Y(n_485) );
INVx2_ASAP7_75t_L g136 ( .A(n_35), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_36), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_37), .A2(n_147), .B(n_206), .C(n_208), .Y(n_205) );
INVxp67_ASAP7_75t_L g251 ( .A(n_38), .Y(n_251) );
CKINVDCx14_ASAP7_75t_R g204 ( .A(n_39), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_40), .A2(n_143), .B(n_226), .C(n_232), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_41), .A2(n_138), .B(n_143), .C(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_42), .A2(n_100), .B1(n_109), .B2(n_720), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_43), .A2(n_116), .B1(n_117), .B2(n_424), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_43), .Y(n_424) );
INVx1_ASAP7_75t_L g103 ( .A(n_44), .Y(n_103) );
INVx1_ASAP7_75t_L g484 ( .A(n_45), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_46), .A2(n_165), .B(n_166), .C(n_169), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_47), .B(n_148), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_48), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_49), .Y(n_247) );
INVx1_ASAP7_75t_L g141 ( .A(n_50), .Y(n_141) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_51), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_52), .B(n_133), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_53), .A2(n_143), .B1(n_153), .B2(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_54), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_55), .Y(n_447) );
CKINVDCx14_ASAP7_75t_R g163 ( .A(n_56), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_57), .A2(n_165), .B(n_208), .C(n_471), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_58), .Y(n_513) );
INVx1_ASAP7_75t_L g469 ( .A(n_59), .Y(n_469) );
INVx1_ASAP7_75t_L g139 ( .A(n_60), .Y(n_139) );
INVx1_ASAP7_75t_L g130 ( .A(n_61), .Y(n_130) );
INVx1_ASAP7_75t_SL g207 ( .A(n_62), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_63), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_64), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g216 ( .A(n_65), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_SL g460 ( .A1(n_66), .A2(n_208), .B(n_461), .C(n_462), .Y(n_460) );
INVxp67_ASAP7_75t_L g463 ( .A(n_67), .Y(n_463) );
INVx1_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_69), .A2(n_133), .B(n_162), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_70), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_71), .A2(n_133), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_72), .Y(n_488) );
INVx1_ASAP7_75t_L g507 ( .A(n_73), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_74), .A2(n_245), .B(n_246), .Y(n_244) );
INVx1_ASAP7_75t_L g191 ( .A(n_75), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_76), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_77), .A2(n_138), .B(n_143), .C(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g132 ( .A1(n_78), .A2(n_133), .B(n_140), .Y(n_132) );
INVx1_ASAP7_75t_L g194 ( .A(n_79), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_80), .B(n_228), .Y(n_501) );
INVx2_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
INVx1_ASAP7_75t_L g181 ( .A(n_82), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_83), .B(n_461), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_84), .A2(n_138), .B(n_143), .C(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g105 ( .A(n_85), .Y(n_105) );
OR2x2_ASAP7_75t_L g428 ( .A(n_85), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g708 ( .A(n_85), .B(n_430), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_86), .A2(n_143), .B(n_215), .C(n_218), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_87), .B(n_160), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_88), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_89), .A2(n_138), .B(n_143), .C(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_90), .Y(n_524) );
INVx1_ASAP7_75t_L g459 ( .A(n_91), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_92), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_93), .B(n_228), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_94), .B(n_126), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_95), .B(n_126), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_98), .A2(n_133), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
BUFx2_ASAP7_75t_L g720 ( .A(n_101), .Y(n_720) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
OR2x2_ASAP7_75t_L g707 ( .A(n_105), .B(n_430), .Y(n_707) );
NOR2x2_ASAP7_75t_L g717 ( .A(n_105), .B(n_429), .Y(n_717) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_436), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g719 ( .A(n_113), .Y(n_719) );
OAI21xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_425), .B(n_433), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g438 ( .A1(n_118), .A2(n_439), .B1(n_707), .B2(n_708), .Y(n_438) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g713 ( .A(n_119), .Y(n_713) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_350), .Y(n_119) );
NOR4xp25_ASAP7_75t_L g120 ( .A(n_121), .B(n_292), .C(n_322), .D(n_332), .Y(n_120) );
OAI211xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_197), .B(n_255), .C(n_282), .Y(n_121) );
OAI222xp33_ASAP7_75t_L g377 ( .A1(n_122), .A2(n_297), .B1(n_378), .B2(n_379), .C1(n_380), .C2(n_381), .Y(n_377) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_172), .Y(n_122) );
AOI33xp33_ASAP7_75t_L g303 ( .A1(n_123), .A2(n_290), .A3(n_291), .B1(n_304), .B2(n_309), .B3(n_311), .Y(n_303) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_123), .A2(n_361), .B(n_363), .C(n_365), .Y(n_360) );
OR2x2_ASAP7_75t_L g376 ( .A(n_123), .B(n_362), .Y(n_376) );
INVx1_ASAP7_75t_L g409 ( .A(n_123), .Y(n_409) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_159), .Y(n_123) );
INVx2_ASAP7_75t_L g286 ( .A(n_124), .Y(n_286) );
AND2x2_ASAP7_75t_L g302 ( .A(n_124), .B(n_188), .Y(n_302) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_124), .Y(n_337) );
AND2x2_ASAP7_75t_L g366 ( .A(n_124), .B(n_159), .Y(n_366) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_132), .B(n_156), .Y(n_124) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_125), .A2(n_189), .B(n_196), .Y(n_188) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_125), .A2(n_202), .B(n_210), .Y(n_201) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g158 ( .A(n_126), .Y(n_158) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_126), .A2(n_457), .B(n_464), .Y(n_456) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g243 ( .A(n_127), .Y(n_243) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_128), .B(n_129), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
BUFx2_ASAP7_75t_L g245 ( .A(n_133), .Y(n_245) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_134), .B(n_138), .Y(n_178) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g231 ( .A(n_135), .Y(n_231) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g154 ( .A(n_136), .Y(n_154) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_137), .Y(n_152) );
INVx3_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g461 ( .A(n_137), .Y(n_461) );
INVx4_ASAP7_75t_SL g155 ( .A(n_138), .Y(n_155) );
BUFx3_ASAP7_75t_L g232 ( .A(n_138), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_142), .B(n_146), .C(n_155), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_SL g162 ( .A1(n_142), .A2(n_155), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_142), .A2(n_155), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_142), .A2(n_155), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_SL g246 ( .A1(n_142), .A2(n_155), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_142), .A2(n_155), .B(n_459), .C(n_460), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_142), .A2(n_155), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_142), .A2(n_155), .B(n_529), .C(n_530), .Y(n_528) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_144), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_147), .B(n_207), .Y(n_206) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_151), .B(n_194), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g249 ( .A1(n_151), .A2(n_228), .B1(n_250), .B2(n_251), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_151), .B(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_152), .A2(n_183), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g452 ( .A(n_153), .Y(n_452) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g218 ( .A(n_155), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_155), .A2(n_178), .B1(n_482), .B2(n_486), .Y(n_481) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_157), .A2(n_467), .B(n_473), .Y(n_466) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_158), .B(n_187), .Y(n_186) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_212), .B(n_219), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_158), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_SL g503 ( .A(n_158), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g266 ( .A(n_159), .Y(n_266) );
BUFx3_ASAP7_75t_L g274 ( .A(n_159), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_159), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g285 ( .A(n_159), .B(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_159), .B(n_173), .Y(n_314) );
AND2x2_ASAP7_75t_L g383 ( .A(n_159), .B(n_317), .Y(n_383) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_171), .Y(n_159) );
INVx1_ASAP7_75t_L g175 ( .A(n_160), .Y(n_175) );
INVx2_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_160), .A2(n_178), .B(n_224), .C(n_225), .Y(n_223) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_160), .A2(n_527), .B(n_533), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx5_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_168), .B(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_168), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
INVx2_ASAP7_75t_SL g277 ( .A(n_172), .Y(n_277) );
OR2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_188), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_173), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g319 ( .A(n_173), .Y(n_319) );
AND2x2_ASAP7_75t_L g330 ( .A(n_173), .B(n_286), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_173), .B(n_315), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_173), .B(n_317), .Y(n_362) );
AND2x2_ASAP7_75t_L g421 ( .A(n_173), .B(n_366), .Y(n_421) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g291 ( .A(n_174), .B(n_188), .Y(n_291) );
AND2x2_ASAP7_75t_L g301 ( .A(n_174), .B(n_302), .Y(n_301) );
BUFx3_ASAP7_75t_L g323 ( .A(n_174), .Y(n_323) );
AND3x2_ASAP7_75t_L g382 ( .A(n_174), .B(n_383), .C(n_384), .Y(n_382) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_186), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_175), .B(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_175), .B(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_175), .B(n_524), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_178), .A2(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_178), .A2(n_447), .B(n_448), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_178), .A2(n_507), .B(n_508), .Y(n_506) );
O2A1O1Ixp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_184), .C(n_185), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_182), .A2(n_185), .B(n_216), .C(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_185), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_185), .A2(n_510), .B(n_511), .Y(n_509) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_188), .Y(n_273) );
INVx1_ASAP7_75t_SL g317 ( .A(n_188), .Y(n_317) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_188), .B(n_266), .C(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_235), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_198), .A2(n_301), .B(n_353), .C(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_200), .B(n_222), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_200), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_SL g369 ( .A(n_200), .Y(n_369) );
AND2x2_ASAP7_75t_L g390 ( .A(n_200), .B(n_237), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_200), .B(n_299), .Y(n_418) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AND2x2_ASAP7_75t_L g263 ( .A(n_201), .B(n_254), .Y(n_263) );
INVx2_ASAP7_75t_L g270 ( .A(n_201), .Y(n_270) );
AND2x2_ASAP7_75t_L g290 ( .A(n_201), .B(n_237), .Y(n_290) );
AND2x2_ASAP7_75t_L g340 ( .A(n_201), .B(n_222), .Y(n_340) );
INVx1_ASAP7_75t_L g344 ( .A(n_201), .Y(n_344) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_209), .Y(n_521) );
INVx2_ASAP7_75t_SL g254 ( .A(n_211), .Y(n_254) );
BUFx2_ASAP7_75t_L g280 ( .A(n_211), .Y(n_280) );
AND2x2_ASAP7_75t_L g407 ( .A(n_211), .B(n_222), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
INVx1_ASAP7_75t_L g253 ( .A(n_221), .Y(n_253) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_221), .A2(n_516), .B(n_523), .Y(n_515) );
INVx3_ASAP7_75t_SL g237 ( .A(n_222), .Y(n_237) );
AND2x2_ASAP7_75t_L g262 ( .A(n_222), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g269 ( .A(n_222), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g299 ( .A(n_222), .B(n_259), .Y(n_299) );
OR2x2_ASAP7_75t_L g308 ( .A(n_222), .B(n_254), .Y(n_308) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_222), .Y(n_326) );
AND2x2_ASAP7_75t_L g331 ( .A(n_222), .B(n_284), .Y(n_331) );
AND2x2_ASAP7_75t_L g359 ( .A(n_222), .B(n_239), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_222), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g397 ( .A(n_222), .B(n_238), .Y(n_397) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_233), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_229), .C(n_230), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_228), .A2(n_450), .B(n_451), .C(n_452), .Y(n_449) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_231), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g321 ( .A(n_237), .B(n_270), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_237), .B(n_263), .Y(n_349) );
AND2x2_ASAP7_75t_L g367 ( .A(n_237), .B(n_284), .Y(n_367) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_254), .Y(n_238) );
AND2x2_ASAP7_75t_L g268 ( .A(n_239), .B(n_254), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_239), .B(n_297), .Y(n_296) );
BUFx3_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
OR2x2_ASAP7_75t_L g354 ( .A(n_239), .B(n_274), .Y(n_354) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_244), .B(n_252), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_241), .A2(n_260), .B(n_261), .Y(n_259) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_241), .A2(n_506), .B(n_512), .Y(n_505) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_SL g497 ( .A1(n_242), .A2(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_243), .A2(n_446), .B(n_453), .Y(n_445) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_243), .A2(n_481), .B(n_487), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_243), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g260 ( .A(n_244), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_252), .Y(n_261) );
AND2x2_ASAP7_75t_L g289 ( .A(n_254), .B(n_259), .Y(n_289) );
INVx1_ASAP7_75t_L g297 ( .A(n_254), .Y(n_297) );
AND2x2_ASAP7_75t_L g392 ( .A(n_254), .B(n_270), .Y(n_392) );
AOI222xp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_264), .B1(n_267), .B2(n_271), .C1(n_275), .C2(n_278), .Y(n_255) );
INVx1_ASAP7_75t_L g387 ( .A(n_256), .Y(n_387) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_262), .Y(n_256) );
AND2x2_ASAP7_75t_L g283 ( .A(n_257), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g294 ( .A(n_257), .B(n_263), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_257), .B(n_285), .Y(n_310) );
OAI222xp33_ASAP7_75t_L g332 ( .A1(n_257), .A2(n_333), .B1(n_338), .B2(n_339), .C1(n_347), .C2(n_349), .Y(n_332) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g320 ( .A(n_259), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_259), .B(n_340), .Y(n_380) );
AND2x2_ASAP7_75t_L g391 ( .A(n_259), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g399 ( .A(n_262), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_264), .B(n_315), .Y(n_378) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_266), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g336 ( .A(n_266), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx3_ASAP7_75t_L g281 ( .A(n_269), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g371 ( .A1(n_269), .A2(n_372), .B(n_375), .C(n_377), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_269), .B(n_306), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_269), .B(n_289), .Y(n_411) );
AND2x2_ASAP7_75t_L g284 ( .A(n_270), .B(n_280), .Y(n_284) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g311 ( .A(n_273), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_274), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g363 ( .A(n_274), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g402 ( .A(n_274), .B(n_302), .Y(n_402) );
INVx1_ASAP7_75t_L g414 ( .A(n_274), .Y(n_414) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_277), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g395 ( .A(n_280), .Y(n_395) );
A2O1A1Ixp33_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_285), .B(n_287), .C(n_291), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_283), .A2(n_313), .B1(n_328), .B2(n_331), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_284), .B(n_298), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_284), .B(n_306), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_285), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g348 ( .A(n_285), .Y(n_348) );
AND2x2_ASAP7_75t_L g355 ( .A(n_285), .B(n_335), .Y(n_355) );
INVx2_ASAP7_75t_L g316 ( .A(n_286), .Y(n_316) );
INVxp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NOR4xp25_ASAP7_75t_L g293 ( .A(n_290), .B(n_294), .C(n_295), .D(n_298), .Y(n_293) );
INVx1_ASAP7_75t_SL g364 ( .A(n_291), .Y(n_364) );
AND2x2_ASAP7_75t_L g408 ( .A(n_291), .B(n_409), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_300), .B(n_303), .C(n_312), .Y(n_292) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_299), .B(n_369), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_301), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_419) );
INVx1_ASAP7_75t_SL g374 ( .A(n_302), .Y(n_374) );
AND2x2_ASAP7_75t_L g413 ( .A(n_302), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_306), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_310), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_311), .B(n_336), .Y(n_396) );
OAI21xp5_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_318), .B(n_320), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g388 ( .A(n_315), .Y(n_388) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g416 ( .A(n_316), .Y(n_416) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_317), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B(n_327), .Y(n_322) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_323), .Y(n_335) );
OR2x2_ASAP7_75t_L g373 ( .A(n_323), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI21xp33_ASAP7_75t_SL g368 ( .A1(n_326), .A2(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_330), .A2(n_357), .B1(n_360), .B2(n_367), .C(n_368), .Y(n_356) );
INVx1_ASAP7_75t_SL g400 ( .A(n_331), .Y(n_400) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
OR2x2_ASAP7_75t_L g347 ( .A(n_335), .B(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g384 ( .A(n_337), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_344), .B2(n_345), .Y(n_339) );
INVx1_ASAP7_75t_L g379 ( .A(n_340), .Y(n_379) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_343), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR4xp25_ASAP7_75t_L g350 ( .A(n_351), .B(n_385), .C(n_398), .D(n_410), .Y(n_350) );
NAND3xp33_ASAP7_75t_SL g351 ( .A(n_352), .B(n_356), .C(n_371), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_354), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_361), .B(n_366), .Y(n_370) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI221xp5_ASAP7_75t_SL g398 ( .A1(n_373), .A2(n_399), .B1(n_400), .B2(n_401), .C(n_403), .Y(n_398) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_375), .A2(n_390), .B(n_391), .C(n_393), .Y(n_389) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_376), .A2(n_394), .B1(n_396), .B2(n_397), .Y(n_393) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_388), .C(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g404 ( .A(n_397), .Y(n_404) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_405), .B(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B1(n_415), .B2(n_417), .C(n_419), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_428), .Y(n_435) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_433), .A2(n_437), .B(n_718), .Y(n_436) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g710 ( .A(n_439), .Y(n_710) );
NAND2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_623), .Y(n_439) );
NOR5xp2_ASAP7_75t_L g440 ( .A(n_441), .B(n_546), .C(n_578), .D(n_593), .E(n_610), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_474), .B(n_493), .C(n_534), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_455), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_443), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_443), .B(n_598), .Y(n_661) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_444), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_444), .B(n_490), .Y(n_547) );
AND2x2_ASAP7_75t_L g588 ( .A(n_444), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_444), .B(n_557), .Y(n_592) );
OR2x2_ASAP7_75t_L g629 ( .A(n_444), .B(n_480), .Y(n_629) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g479 ( .A(n_445), .B(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g537 ( .A(n_445), .Y(n_537) );
OR2x2_ASAP7_75t_L g700 ( .A(n_445), .B(n_540), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_455), .A2(n_603), .B1(n_604), .B2(n_607), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_455), .B(n_537), .Y(n_686) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .Y(n_455) );
AND2x2_ASAP7_75t_L g492 ( .A(n_456), .B(n_480), .Y(n_492) );
AND2x2_ASAP7_75t_L g539 ( .A(n_456), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g544 ( .A(n_456), .Y(n_544) );
INVx3_ASAP7_75t_L g557 ( .A(n_456), .Y(n_557) );
OR2x2_ASAP7_75t_L g577 ( .A(n_456), .B(n_540), .Y(n_577) );
AND2x2_ASAP7_75t_L g596 ( .A(n_456), .B(n_466), .Y(n_596) );
BUFx2_ASAP7_75t_L g628 ( .A(n_456), .Y(n_628) );
AND2x4_ASAP7_75t_L g543 ( .A(n_465), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g478 ( .A(n_466), .Y(n_478) );
INVx2_ASAP7_75t_L g491 ( .A(n_466), .Y(n_491) );
OR2x2_ASAP7_75t_L g559 ( .A(n_466), .B(n_540), .Y(n_559) );
AND2x2_ASAP7_75t_L g589 ( .A(n_466), .B(n_480), .Y(n_589) );
AND2x2_ASAP7_75t_L g606 ( .A(n_466), .B(n_537), .Y(n_606) );
AND2x2_ASAP7_75t_L g646 ( .A(n_466), .B(n_557), .Y(n_646) );
AND2x2_ASAP7_75t_SL g682 ( .A(n_466), .B(n_492), .Y(n_682) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp33_ASAP7_75t_SL g475 ( .A(n_476), .B(n_489), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_477), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
OAI21xp33_ASAP7_75t_L g620 ( .A1(n_478), .A2(n_492), .B(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_478), .B(n_480), .Y(n_676) );
AND2x2_ASAP7_75t_L g612 ( .A(n_479), .B(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g540 ( .A(n_480), .Y(n_540) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_480), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_489), .B(n_537), .Y(n_705) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_490), .A2(n_648), .B1(n_649), .B2(n_654), .Y(n_647) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x2_ASAP7_75t_L g538 ( .A(n_491), .B(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g576 ( .A(n_491), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g613 ( .A(n_491), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_492), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g667 ( .A(n_492), .Y(n_667) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_514), .Y(n_494) );
INVx4_ASAP7_75t_L g553 ( .A(n_495), .Y(n_553) );
AND2x2_ASAP7_75t_L g631 ( .A(n_495), .B(n_598), .Y(n_631) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_505), .Y(n_495) );
INVx3_ASAP7_75t_L g550 ( .A(n_496), .Y(n_550) );
AND2x2_ASAP7_75t_L g564 ( .A(n_496), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g568 ( .A(n_496), .Y(n_568) );
INVx2_ASAP7_75t_L g582 ( .A(n_496), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_496), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g639 ( .A(n_496), .B(n_634), .Y(n_639) );
AND2x2_ASAP7_75t_L g704 ( .A(n_496), .B(n_674), .Y(n_704) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
AND2x2_ASAP7_75t_L g545 ( .A(n_505), .B(n_526), .Y(n_545) );
INVx2_ASAP7_75t_L g565 ( .A(n_505), .Y(n_565) );
INVx1_ASAP7_75t_L g570 ( .A(n_514), .Y(n_570) );
AND2x2_ASAP7_75t_L g616 ( .A(n_514), .B(n_564), .Y(n_616) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_525), .Y(n_514) );
INVx2_ASAP7_75t_L g555 ( .A(n_515), .Y(n_555) );
INVx1_ASAP7_75t_L g563 ( .A(n_515), .Y(n_563) );
AND2x2_ASAP7_75t_L g581 ( .A(n_515), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_515), .B(n_565), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_522), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_521), .Y(n_518) );
AND2x2_ASAP7_75t_L g598 ( .A(n_525), .B(n_555), .Y(n_598) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g551 ( .A(n_526), .Y(n_551) );
AND2x2_ASAP7_75t_L g634 ( .A(n_526), .B(n_565), .Y(n_634) );
OAI21xp5_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_541), .B(n_545), .Y(n_534) );
INVx1_ASAP7_75t_SL g579 ( .A(n_535), .Y(n_579) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_536), .B(n_543), .Y(n_636) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g585 ( .A(n_537), .B(n_540), .Y(n_585) );
AND2x2_ASAP7_75t_L g614 ( .A(n_537), .B(n_558), .Y(n_614) );
OR2x2_ASAP7_75t_L g617 ( .A(n_537), .B(n_577), .Y(n_617) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_538), .A2(n_630), .B1(n_682), .B2(n_683), .C1(n_685), .C2(n_687), .Y(n_681) );
BUFx2_ASAP7_75t_L g595 ( .A(n_540), .Y(n_595) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g584 ( .A(n_543), .B(n_585), .Y(n_584) );
INVx3_ASAP7_75t_SL g601 ( .A(n_543), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_543), .B(n_595), .Y(n_655) );
AND2x2_ASAP7_75t_L g590 ( .A(n_545), .B(n_550), .Y(n_590) );
INVx1_ASAP7_75t_L g609 ( .A(n_545), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_548), .B1(n_552), .B2(n_556), .C(n_560), .Y(n_546) );
OR2x2_ASAP7_75t_L g618 ( .A(n_548), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x2_ASAP7_75t_L g603 ( .A(n_550), .B(n_573), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_550), .B(n_563), .Y(n_643) );
AND2x2_ASAP7_75t_L g648 ( .A(n_550), .B(n_598), .Y(n_648) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_550), .Y(n_658) );
NAND2x1_ASAP7_75t_SL g669 ( .A(n_550), .B(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g554 ( .A(n_551), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g574 ( .A(n_551), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_551), .B(n_569), .Y(n_600) );
INVx1_ASAP7_75t_L g666 ( .A(n_551), .Y(n_666) );
INVx1_ASAP7_75t_L g641 ( .A(n_552), .Y(n_641) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g653 ( .A(n_553), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g665 ( .A(n_553), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g670 ( .A(n_554), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_554), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g573 ( .A(n_555), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_555), .B(n_565), .Y(n_586) );
INVx1_ASAP7_75t_L g652 ( .A(n_555), .Y(n_652) );
INVx1_ASAP7_75t_L g673 ( .A(n_556), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI21xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_566), .B(n_575), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
AND2x2_ASAP7_75t_L g706 ( .A(n_562), .B(n_639), .Y(n_706) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g674 ( .A(n_563), .B(n_634), .Y(n_674) );
AOI32xp33_ASAP7_75t_L g587 ( .A1(n_564), .A2(n_570), .A3(n_588), .B1(n_590), .B2(n_591), .Y(n_587) );
AOI322xp5_ASAP7_75t_L g689 ( .A1(n_564), .A2(n_596), .A3(n_679), .B1(n_690), .B2(n_691), .C1(n_692), .C2(n_694), .Y(n_689) );
INVx2_ASAP7_75t_L g569 ( .A(n_565), .Y(n_569) );
INVx1_ASAP7_75t_L g679 ( .A(n_565), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_570), .B1(n_571), .B2(n_572), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_567), .B(n_573), .Y(n_622) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_568), .B(n_634), .Y(n_684) );
INVx1_ASAP7_75t_L g571 ( .A(n_569), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_569), .B(n_598), .Y(n_688) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_577), .B(n_672), .Y(n_671) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_580), .B1(n_583), .B2(n_586), .C(n_587), .Y(n_578) );
OR2x2_ASAP7_75t_L g599 ( .A(n_580), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g608 ( .A(n_580), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g633 ( .A(n_581), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g637 ( .A(n_591), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_597), .B1(n_599), .B2(n_601), .C(n_602), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_595), .A2(n_626), .B1(n_630), .B2(n_631), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_596), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g701 ( .A(n_596), .Y(n_701) );
INVx1_ASAP7_75t_L g695 ( .A(n_598), .Y(n_695) );
INVx1_ASAP7_75t_SL g630 ( .A(n_599), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_601), .B(n_629), .Y(n_691) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_606), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g672 ( .A(n_606), .Y(n_672) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g610 ( .A1(n_611), .A2(n_615), .B1(n_617), .B2(n_618), .C(n_620), .Y(n_610) );
NOR2xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_614), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_612), .A2(n_630), .B1(n_676), .B2(n_677), .Y(n_675) );
CKINVDCx14_ASAP7_75t_R g615 ( .A(n_616), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_617), .A2(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR3xp33_ASAP7_75t_SL g623 ( .A(n_624), .B(n_656), .C(n_680), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_625), .B(n_632), .C(n_640), .D(n_647), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g703 ( .A(n_628), .Y(n_703) );
INVx3_ASAP7_75t_SL g697 ( .A(n_629), .Y(n_697) );
OR2x2_ASAP7_75t_L g702 ( .A(n_629), .B(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B1(n_637), .B2(n_639), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_634), .B(n_652), .Y(n_693) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_642), .B(n_644), .Y(n_640) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_659), .B(n_662), .C(n_675), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g690 ( .A(n_661), .Y(n_690) );
AOI222xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_667), .B1(n_668), .B2(n_671), .C1(n_673), .C2(n_674), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND4xp25_ASAP7_75t_SL g699 ( .A(n_672), .B(n_700), .C(n_701), .D(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND3xp33_ASAP7_75t_SL g680 ( .A(n_681), .B(n_689), .C(n_698), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_707), .A2(n_710), .B1(n_711), .B2(n_713), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_708), .Y(n_712) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
endmodule