module fake_ibex_9_n_2114 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_366, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_2114);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_366;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_2114;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_766;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_1930;
wire n_452;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_1971;
wire n_879;
wire n_1957;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_2112;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1936;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2076;
wire n_1036;
wire n_974;
wire n_1831;
wire n_608;
wire n_864;
wire n_412;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_2077;
wire n_517;
wire n_817;
wire n_2095;
wire n_555;
wire n_951;
wire n_2053;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1952;
wire n_785;
wire n_1624;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_2108;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_2078;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_2093;
wire n_786;
wire n_505;
wire n_2043;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1433;
wire n_1314;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_2083;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2013;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_665;
wire n_1101;
wire n_2079;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1992;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_2104;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2092;
wire n_566;
wire n_416;
wire n_581;
wire n_1472;
wire n_1365;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2016;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_519;
wire n_1843;
wire n_408;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_1902;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_SL g397 ( 
.A(n_265),
.Y(n_397)
);

INVxp33_ASAP7_75t_L g398 ( 
.A(n_380),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_247),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_275),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_157),
.Y(n_404)
);

BUFx5_ASAP7_75t_L g405 ( 
.A(n_105),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_350),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_305),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_220),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_233),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_234),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_133),
.Y(n_412)
);

INVxp33_ASAP7_75t_SL g413 ( 
.A(n_0),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_205),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_144),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_354),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_156),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_201),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_322),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_166),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_26),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_16),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_318),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_126),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_41),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_174),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_121),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_17),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_39),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_300),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_321),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_278),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_317),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_346),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_101),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_227),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_56),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_189),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_327),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_181),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_196),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_193),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_237),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_99),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_289),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_84),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_193),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_86),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_352),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_365),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_92),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_292),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_357),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_335),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_102),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_307),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_276),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_170),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_366),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_386),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_6),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_344),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_177),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_373),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_343),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_383),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_198),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_51),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_18),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_390),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_280),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_272),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_147),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_210),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_R g476 ( 
.A(n_308),
.B(n_328),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_297),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_140),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_26),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_283),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_356),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_107),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_80),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_315),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_231),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_160),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_330),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_329),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_149),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_89),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_296),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_202),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_293),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_22),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_21),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_89),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_359),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_13),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_178),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_225),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_270),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_29),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_145),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_41),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_374),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_215),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_360),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_391),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_12),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_164),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_301),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_302),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_164),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_252),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_70),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_110),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_113),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_342),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_290),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_334),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_19),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_368),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_117),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_232),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_370),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_254),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_371),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_148),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_331),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_176),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_134),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_246),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_254),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_65),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_158),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_175),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_159),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_336),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_148),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_298),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_195),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_123),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_393),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_168),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_340),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_355),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_157),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_2),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_205),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_222),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_122),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_187),
.Y(n_553)
);

CKINVDCx14_ASAP7_75t_R g554 ( 
.A(n_105),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_79),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_143),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_294),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_81),
.B(n_162),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_1),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_231),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_200),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_323),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_268),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_27),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_332),
.Y(n_565)
);

NOR2xp67_ASAP7_75t_L g566 ( 
.A(n_118),
.B(n_115),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_337),
.Y(n_567)
);

INVxp33_ASAP7_75t_SL g568 ( 
.A(n_364),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_54),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_291),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_358),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_32),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_58),
.Y(n_573)
);

NOR2xp67_ASAP7_75t_L g574 ( 
.A(n_320),
.B(n_255),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_247),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_326),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_97),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_378),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_353),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_99),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_117),
.Y(n_581)
);

BUFx8_ASAP7_75t_SL g582 ( 
.A(n_13),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_351),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_256),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_382),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_165),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_129),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_3),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_190),
.Y(n_589)
);

CKINVDCx14_ASAP7_75t_R g590 ( 
.A(n_167),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_129),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_339),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_208),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_376),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_220),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_216),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_299),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_349),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_224),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_369),
.Y(n_600)
);

BUFx5_ASAP7_75t_L g601 ( 
.A(n_138),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_319),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_218),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_361),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_248),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_54),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_375),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_202),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_138),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_21),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_377),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_4),
.Y(n_612)
);

BUFx8_ASAP7_75t_SL g613 ( 
.A(n_381),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_214),
.Y(n_614)
);

CKINVDCx14_ASAP7_75t_R g615 ( 
.A(n_372),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_295),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_215),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_85),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_104),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_385),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_387),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_250),
.Y(n_622)
);

INVxp33_ASAP7_75t_L g623 ( 
.A(n_250),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_181),
.Y(n_624)
);

BUFx10_ASAP7_75t_L g625 ( 
.A(n_345),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_199),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_341),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_175),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_266),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_217),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_31),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_261),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_35),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_186),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_379),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_395),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_241),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_7),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_242),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_103),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_394),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_38),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_76),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_249),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_244),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_240),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_167),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_253),
.Y(n_648)
);

BUFx5_ASAP7_75t_L g649 ( 
.A(n_114),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_333),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_229),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_120),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_43),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_132),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_392),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_259),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_1),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_52),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_151),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_285),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_131),
.Y(n_661)
);

INVxp33_ASAP7_75t_L g662 ( 
.A(n_258),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_232),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_282),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_103),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_388),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_312),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_169),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_257),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_6),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_623),
.B(n_0),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_405),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_612),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g674 ( 
.A(n_399),
.B(n_2),
.Y(n_674)
);

OA21x2_ASAP7_75t_L g675 ( 
.A1(n_401),
.A2(n_262),
.B(n_260),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_405),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_612),
.Y(n_677)
);

NOR2x1_ASAP7_75t_L g678 ( 
.A(n_612),
.B(n_670),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_405),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_434),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_434),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_434),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_434),
.Y(n_683)
);

OAI22x1_ASAP7_75t_SL g684 ( 
.A1(n_399),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_419),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_521),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_405),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_405),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_405),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_601),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_601),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_601),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_601),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_601),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_423),
.B(n_5),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_521),
.Y(n_696)
);

BUFx8_ASAP7_75t_L g697 ( 
.A(n_655),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_521),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_601),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_649),
.Y(n_700)
);

OA21x2_ASAP7_75t_L g701 ( 
.A1(n_401),
.A2(n_264),
.B(n_263),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_649),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_521),
.Y(n_703)
);

NAND2x1p5_ASAP7_75t_L g704 ( 
.A(n_423),
.B(n_267),
.Y(n_704)
);

OAI22x1_ASAP7_75t_R g705 ( 
.A1(n_410),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_448),
.B(n_8),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_649),
.Y(n_708)
);

CKINVDCx6p67_ASAP7_75t_R g709 ( 
.A(n_492),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_649),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_649),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_649),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_412),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_500),
.B(n_9),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_606),
.B(n_10),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_412),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_421),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_431),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_421),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_565),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_431),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_436),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_565),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_617),
.B(n_11),
.Y(n_724)
);

BUFx8_ASAP7_75t_L g725 ( 
.A(n_397),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_448),
.B(n_14),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_455),
.A2(n_271),
.B(n_269),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_511),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_455),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_511),
.B(n_15),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_484),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_419),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_565),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_436),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_484),
.Y(n_735)
);

BUFx12f_ASAP7_75t_L g736 ( 
.A(n_625),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_670),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_438),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_438),
.Y(n_739)
);

CKINVDCx11_ASAP7_75t_R g740 ( 
.A(n_410),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_512),
.A2(n_274),
.B(n_273),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_462),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_512),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_623),
.B(n_15),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_570),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_646),
.B(n_277),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_470),
.Y(n_747)
);

AND2x2_ASAP7_75t_SL g748 ( 
.A(n_409),
.B(n_396),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_563),
.B(n_16),
.Y(n_749)
);

NOR2x1_ASAP7_75t_L g750 ( 
.A(n_574),
.B(n_17),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_570),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_571),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_650),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_440),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_571),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_440),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_462),
.B(n_18),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_475),
.B(n_19),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_475),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_487),
.Y(n_760)
);

OA21x2_ASAP7_75t_L g761 ( 
.A1(n_592),
.A2(n_281),
.B(n_279),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_592),
.A2(n_286),
.B(n_284),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_411),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_604),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_487),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_662),
.B(n_398),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_490),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_554),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_768)
);

OA21x2_ASAP7_75t_L g769 ( 
.A1(n_636),
.A2(n_288),
.B(n_287),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_490),
.B(n_24),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_636),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_662),
.B(n_27),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_650),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_497),
.B(n_28),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_554),
.B(n_29),
.Y(n_775)
);

BUFx8_ASAP7_75t_SL g776 ( 
.A(n_582),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_666),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_757),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_766),
.B(n_519),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_754),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_672),
.Y(n_781)
);

INVxp33_ASAP7_75t_L g782 ( 
.A(n_766),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_754),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_685),
.B(n_416),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_673),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_757),
.A2(n_415),
.B1(n_417),
.B2(n_408),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_757),
.A2(n_426),
.B1(n_430),
.B2(n_427),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_747),
.B(n_404),
.Y(n_788)
);

AND3x2_ASAP7_75t_L g789 ( 
.A(n_685),
.B(n_504),
.C(n_480),
.Y(n_789)
);

OR2x6_ASAP7_75t_L g790 ( 
.A(n_736),
.B(n_566),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_736),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_673),
.B(n_585),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_758),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_695),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_775),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_676),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_758),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_758),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_775),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_673),
.B(n_590),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_758),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_676),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_679),
.Y(n_803)
);

INVxp33_ASAP7_75t_L g804 ( 
.A(n_671),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_679),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_768),
.A2(n_422),
.B1(n_491),
.B2(n_411),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_709),
.B(n_596),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_756),
.Y(n_808)
);

OAI21xp33_ASAP7_75t_SL g809 ( 
.A1(n_748),
.A2(n_441),
.B(n_439),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_695),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_687),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_770),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_764),
.B(n_557),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_774),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_SL g815 ( 
.A(n_671),
.B(n_446),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_707),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_687),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_L g818 ( 
.A1(n_714),
.A2(n_422),
.B1(n_543),
.B2(n_491),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_689),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_707),
.B(n_666),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_726),
.B(n_402),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_726),
.B(n_403),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_689),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_690),
.Y(n_824)
);

BUFx10_ASAP7_75t_L g825 ( 
.A(n_748),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_744),
.B(n_471),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_748),
.A2(n_413),
.B1(n_568),
.B2(n_451),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_726),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_692),
.Y(n_829)
);

INVxp33_ASAP7_75t_L g830 ( 
.A(n_744),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_SL g831 ( 
.A1(n_763),
.A2(n_543),
.B1(n_561),
.B2(n_556),
.Y(n_831)
);

INVxp67_ASAP7_75t_SL g832 ( 
.A(n_772),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_681),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_730),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_730),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_728),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_730),
.Y(n_837)
);

AND3x1_ASAP7_75t_L g838 ( 
.A(n_772),
.B(n_443),
.C(n_442),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_730),
.B(n_406),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_697),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_715),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_697),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_677),
.Y(n_843)
);

INVx4_ASAP7_75t_L g844 ( 
.A(n_704),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_678),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_737),
.B(n_458),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_776),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_704),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_678),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_693),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_725),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_697),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_737),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_688),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_688),
.B(n_418),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_725),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_691),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_691),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_725),
.B(n_502),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_694),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_694),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_724),
.B(n_608),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_706),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_699),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_765),
.B(n_497),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_706),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_711),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_711),
.Y(n_868)
);

BUFx4f_ASAP7_75t_L g869 ( 
.A(n_704),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_700),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_681),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_732),
.Y(n_872)
);

AND2x6_ASAP7_75t_L g873 ( 
.A(n_750),
.B(n_424),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_746),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_681),
.Y(n_875)
);

INVx5_ASAP7_75t_L g876 ( 
.A(n_680),
.Y(n_876)
);

BUFx10_ASAP7_75t_L g877 ( 
.A(n_749),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_712),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_700),
.B(n_432),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_725),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_702),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_708),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_708),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_710),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_718),
.A2(n_444),
.B1(n_452),
.B2(n_445),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_765),
.B(n_767),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_682),
.Y(n_887)
);

AO22x2_ASAP7_75t_L g888 ( 
.A1(n_684),
.A2(n_558),
.B1(n_525),
.B2(n_536),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_718),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_746),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_721),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_740),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_721),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_682),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_765),
.B(n_458),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_729),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_682),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_683),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_746),
.B(n_400),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_731),
.B(n_453),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_680),
.Y(n_901)
);

AND2x6_ASAP7_75t_L g902 ( 
.A(n_750),
.B(n_454),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_675),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_767),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_713),
.B(n_460),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_731),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_735),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_713),
.B(n_457),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_743),
.B(n_461),
.Y(n_909)
);

AO21x2_ASAP7_75t_L g910 ( 
.A1(n_727),
.A2(n_477),
.B(n_463),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_745),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_716),
.B(n_607),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_716),
.B(n_481),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_705),
.B(n_582),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_751),
.A2(n_413),
.B1(n_451),
.B2(n_446),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_686),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_717),
.B(n_719),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_751),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_752),
.A2(n_568),
.B1(n_583),
.B2(n_576),
.Y(n_919)
);

NAND2xp33_ASAP7_75t_R g920 ( 
.A(n_675),
.B(n_665),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_752),
.B(n_486),
.Y(n_921)
);

AND2x6_ASAP7_75t_L g922 ( 
.A(n_755),
.B(n_488),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_771),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_717),
.B(n_489),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_777),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_719),
.B(n_514),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_777),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_686),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_686),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_680),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_675),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_722),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_734),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_701),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_842),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_869),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_832),
.B(n_607),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_832),
.B(n_826),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_792),
.B(n_738),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_821),
.A2(n_741),
.B(n_701),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_841),
.B(n_611),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_788),
.B(n_674),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_804),
.B(n_738),
.Y(n_943)
);

NOR2x1p5_ASAP7_75t_L g944 ( 
.A(n_892),
.B(n_674),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_800),
.B(n_471),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_780),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_804),
.B(n_739),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_830),
.B(n_739),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_851),
.B(n_625),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_813),
.B(n_615),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_784),
.B(n_742),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_795),
.Y(n_952)
);

OAI22xp33_ASAP7_75t_L g953 ( 
.A1(n_827),
.A2(n_583),
.B1(n_597),
.B2(n_576),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_801),
.A2(n_759),
.B1(n_760),
.B2(n_742),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_795),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_880),
.B(n_629),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_830),
.B(n_759),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_783),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_784),
.B(n_760),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_880),
.B(n_629),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_856),
.B(n_629),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_779),
.B(n_407),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_782),
.A2(n_664),
.B1(n_667),
.B2(n_597),
.Y(n_963)
);

NAND2x1_ASAP7_75t_L g964 ( 
.A(n_794),
.B(n_701),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_862),
.B(n_414),
.Y(n_965)
);

O2A1O1Ixp5_ASAP7_75t_L g966 ( 
.A1(n_903),
.A2(n_578),
.B(n_498),
.C(n_506),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_859),
.B(n_494),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_818),
.B(n_425),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_809),
.A2(n_667),
.B1(n_664),
.B2(n_428),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_859),
.B(n_890),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_799),
.B(n_420),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_890),
.B(n_508),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_808),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_799),
.B(n_433),
.Y(n_974)
);

AND2x4_ASAP7_75t_SL g975 ( 
.A(n_840),
.B(n_852),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_905),
.B(n_435),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_845),
.B(n_509),
.Y(n_977)
);

BUFx6f_ASAP7_75t_SL g978 ( 
.A(n_914),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_844),
.B(n_450),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_844),
.B(n_465),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_918),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_886),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_912),
.B(n_466),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_785),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_816),
.A2(n_741),
.B(n_459),
.C(n_464),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_846),
.B(n_467),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_849),
.B(n_513),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_848),
.B(n_472),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_895),
.B(n_473),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_791),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_904),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_917),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_853),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_838),
.A2(n_437),
.B1(n_449),
.B2(n_429),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_874),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_810),
.B(n_933),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_874),
.B(n_523),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_786),
.B(n_528),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_787),
.B(n_530),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_787),
.B(n_778),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_801),
.A2(n_456),
.B1(n_469),
.B2(n_468),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_904),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_915),
.Y(n_1003)
);

NOR3xp33_ASAP7_75t_L g1004 ( 
.A(n_806),
.B(n_559),
.C(n_550),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_793),
.B(n_539),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_797),
.B(n_541),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_889),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_798),
.B(n_547),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_865),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_785),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_807),
.B(n_919),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_815),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_836),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_891),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_822),
.B(n_520),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_828),
.Y(n_1016)
);

AND2x2_ASAP7_75t_SL g1017 ( 
.A(n_899),
.B(n_701),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_839),
.B(n_526),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_839),
.B(n_812),
.Y(n_1019)
);

OAI21xp33_ASAP7_75t_L g1020 ( 
.A1(n_837),
.A2(n_478),
.B(n_474),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_926),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_926),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_789),
.B(n_447),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_814),
.A2(n_482),
.B1(n_483),
.B2(n_479),
.Y(n_1024)
);

CKINVDCx11_ASAP7_75t_R g1025 ( 
.A(n_914),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_843),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_877),
.B(n_820),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_834),
.A2(n_495),
.B1(n_499),
.B2(n_493),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_834),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_932),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_877),
.B(n_544),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_893),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_789),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_896),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_L g1035 ( 
.A(n_835),
.B(n_546),
.Y(n_1035)
);

AOI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_818),
.A2(n_684),
.B1(n_510),
.B2(n_515),
.C(n_507),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_906),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_907),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_914),
.B(n_447),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_911),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_820),
.B(n_485),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_885),
.A2(n_790),
.B1(n_888),
.B2(n_923),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_825),
.B(n_562),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_873),
.B(n_496),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_825),
.B(n_567),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_790),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_815),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_L g1048 ( 
.A(n_873),
.B(n_579),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_925),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_873),
.B(n_501),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_927),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_902),
.B(n_505),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_902),
.A2(n_529),
.B1(n_532),
.B2(n_527),
.Y(n_1053)
);

BUFx3_ASAP7_75t_L g1054 ( 
.A(n_790),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_902),
.A2(n_538),
.B1(n_545),
.B2(n_537),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_900),
.Y(n_1056)
);

NAND2xp33_ASAP7_75t_L g1057 ( 
.A(n_922),
.B(n_594),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_872),
.B(n_573),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_922),
.Y(n_1059)
);

NOR3xp33_ASAP7_75t_L g1060 ( 
.A(n_806),
.B(n_609),
.C(n_552),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_908),
.B(n_564),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_900),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_888),
.B(n_705),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_908),
.B(n_598),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_913),
.B(n_600),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_909),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_903),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_924),
.B(n_855),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_924),
.B(n_569),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_855),
.B(n_572),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_L g1071 ( 
.A(n_847),
.B(n_30),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_909),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_931),
.B(n_613),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_879),
.B(n_602),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_921),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_931),
.A2(n_503),
.B1(n_517),
.B2(n_516),
.Y(n_1076)
);

BUFx8_ASAP7_75t_L g1077 ( 
.A(n_888),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_854),
.B(n_616),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_921),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_934),
.B(n_514),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_934),
.A2(n_762),
.B(n_761),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_781),
.Y(n_1082)
);

BUFx5_ASAP7_75t_L g1083 ( 
.A(n_857),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_901),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_858),
.B(n_614),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_864),
.B(n_619),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_870),
.B(n_881),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_881),
.B(n_620),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_910),
.A2(n_883),
.B(n_882),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_910),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_883),
.B(n_624),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_884),
.B(n_633),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_884),
.B(n_639),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_796),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_802),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_803),
.B(n_621),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_803),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_860),
.B(n_627),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_805),
.B(n_632),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_811),
.B(n_647),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_817),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_831),
.A2(n_657),
.B1(n_654),
.B2(n_518),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_831),
.B(n_524),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_819),
.B(n_533),
.C(n_531),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_823),
.B(n_635),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_824),
.B(n_641),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_824),
.B(n_660),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_861),
.B(n_534),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_901),
.Y(n_1109)
);

NOR2xp67_ASAP7_75t_L g1110 ( 
.A(n_876),
.B(n_30),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_920),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_863),
.A2(n_762),
.B(n_761),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_829),
.B(n_555),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_850),
.B(n_555),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_866),
.B(n_535),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_867),
.B(n_540),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_868),
.B(n_542),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_850),
.B(n_560),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_878),
.B(n_560),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_930),
.B(n_586),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_930),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_887),
.A2(n_549),
.B1(n_553),
.B2(n_548),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_SL g1123 ( 
.A1(n_929),
.A2(n_556),
.B1(n_575),
.B2(n_561),
.Y(n_1123)
);

O2A1O1Ixp5_ASAP7_75t_L g1124 ( 
.A1(n_887),
.A2(n_595),
.B(n_618),
.C(n_591),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_935),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_964),
.A2(n_762),
.B(n_761),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1082),
.Y(n_1127)
);

BUFx8_ASAP7_75t_L g1128 ( 
.A(n_978),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_992),
.A2(n_605),
.B1(n_610),
.B2(n_575),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1083),
.B(n_643),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1011),
.A2(n_610),
.B1(n_626),
.B2(n_605),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1003),
.A2(n_968),
.B(n_1004),
.C(n_938),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1081),
.A2(n_940),
.B(n_1112),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_952),
.B(n_955),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1004),
.B(n_476),
.C(n_762),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1016),
.A2(n_640),
.B1(n_644),
.B2(n_626),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_970),
.B(n_640),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1089),
.A2(n_1087),
.B(n_1017),
.Y(n_1138)
);

NOR2xp67_ASAP7_75t_L g1139 ( 
.A(n_1033),
.B(n_31),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1017),
.A2(n_769),
.B(n_894),
.Y(n_1140)
);

AOI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1090),
.A2(n_769),
.B(n_894),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1083),
.B(n_643),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_937),
.B(n_577),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_996),
.A2(n_769),
.B(n_898),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_959),
.B(n_580),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_963),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1067),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_959),
.B(n_982),
.Y(n_1148)
);

NOR2x1_ASAP7_75t_R g1149 ( 
.A(n_1025),
.B(n_1054),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1060),
.A2(n_581),
.B(n_587),
.C(n_584),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1068),
.A2(n_589),
.B(n_593),
.C(n_588),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_970),
.B(n_613),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1058),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1083),
.B(n_652),
.Y(n_1154)
);

AOI33xp33_ASAP7_75t_L g1155 ( 
.A1(n_1001),
.A2(n_630),
.A3(n_622),
.B1(n_634),
.B2(n_631),
.B3(n_628),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_945),
.A2(n_928),
.B(n_916),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1060),
.A2(n_645),
.B(n_648),
.C(n_637),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1103),
.A2(n_653),
.B(n_656),
.C(n_651),
.Y(n_1158)
);

INVx4_ASAP7_75t_L g1159 ( 
.A(n_975),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_966),
.A2(n_928),
.B(n_659),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_995),
.B(n_618),
.Y(n_1161)
);

AO22x1_ASAP7_75t_L g1162 ( 
.A1(n_1077),
.A2(n_661),
.B1(n_668),
.B2(n_658),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_L g1163 ( 
.A(n_953),
.B(n_652),
.C(n_476),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_L g1164 ( 
.A(n_953),
.B(n_652),
.C(n_32),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1104),
.A2(n_696),
.B(n_686),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1019),
.A2(n_551),
.B(n_599),
.C(n_522),
.Y(n_1166)
);

AND2x6_ASAP7_75t_L g1167 ( 
.A(n_1059),
.B(n_522),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_R g1168 ( 
.A(n_978),
.B(n_33),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_1080),
.Y(n_1169)
);

OAI22x1_ASAP7_75t_L g1170 ( 
.A1(n_969),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1170)
);

AOI21xp33_ASAP7_75t_L g1171 ( 
.A1(n_1027),
.A2(n_599),
.B(n_551),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1047),
.A2(n_1042),
.B1(n_1027),
.B2(n_1012),
.Y(n_1172)
);

AOI21xp33_ASAP7_75t_L g1173 ( 
.A1(n_1047),
.A2(n_599),
.B(n_551),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_939),
.B(n_599),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1111),
.B(n_603),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1080),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1080),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_1063),
.B(n_638),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_939),
.B(n_638),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1073),
.B(n_941),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_1007),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1000),
.A2(n_663),
.B(n_669),
.C(n_642),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1014),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1029),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1076),
.A2(n_669),
.B1(n_663),
.B2(n_680),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_1049),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_967),
.A2(n_669),
.B(n_663),
.C(n_686),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1123),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1029),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_943),
.B(n_669),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_967),
.A2(n_698),
.B(n_703),
.C(n_696),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_947),
.B(n_948),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_966),
.A2(n_871),
.B(n_833),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_957),
.B(n_36),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1046),
.B(n_37),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1026),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_957),
.B(n_37),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1063),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_990),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_1039),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1124),
.A2(n_875),
.B(n_871),
.Y(n_1201)
);

BUFx4_ASAP7_75t_SL g1202 ( 
.A(n_958),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_972),
.B(n_40),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_972),
.B(n_42),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1076),
.A2(n_703),
.B1(n_720),
.B2(n_698),
.Y(n_1205)
);

BUFx4f_ASAP7_75t_L g1206 ( 
.A(n_936),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_951),
.B(n_44),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1109),
.Y(n_1208)
);

CKINVDCx6p67_ASAP7_75t_R g1209 ( 
.A(n_997),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_994),
.B(n_45),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1028),
.B(n_45),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1124),
.A2(n_897),
.B(n_723),
.Y(n_1212)
);

OAI21xp33_ASAP7_75t_L g1213 ( 
.A1(n_1061),
.A2(n_733),
.B(n_723),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_973),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_R g1215 ( 
.A(n_1077),
.B(n_46),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1023),
.B(n_46),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1005),
.A2(n_1008),
.B(n_1006),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1024),
.B(n_47),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_971),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1031),
.B(n_47),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1021),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_998),
.A2(n_773),
.B1(n_753),
.B2(n_50),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1022),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_993),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1015),
.A2(n_1018),
.B(n_1074),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_1036),
.B(n_48),
.C(n_49),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1069),
.B(n_48),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1018),
.A2(n_773),
.B(n_52),
.C(n_49),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1064),
.A2(n_773),
.B(n_56),
.C(n_53),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_999),
.A2(n_773),
.B1(n_57),
.B2(n_53),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_950),
.A2(n_58),
.B1(n_55),
.B2(n_57),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1065),
.B(n_55),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1102),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_954),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_979),
.B(n_980),
.Y(n_1235)
);

OAI21xp33_ASAP7_75t_L g1236 ( 
.A1(n_974),
.A2(n_62),
.B(n_63),
.Y(n_1236)
);

AO21x1_ASAP7_75t_L g1237 ( 
.A1(n_1088),
.A2(n_63),
.B(n_64),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_954),
.A2(n_1078),
.B1(n_1088),
.B2(n_1032),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_944),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1053),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1085),
.B(n_64),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1009),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1020),
.A2(n_1041),
.B(n_1086),
.C(n_1048),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1078),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1244)
);

AO32x2_ASAP7_75t_L g1245 ( 
.A1(n_1062),
.A2(n_68),
.A3(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1034),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1246)
);

BUFx8_ASAP7_75t_L g1247 ( 
.A(n_1075),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1074),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1248)
);

OR2x2_ASAP7_75t_SL g1249 ( 
.A(n_1044),
.B(n_72),
.Y(n_1249)
);

BUFx8_ASAP7_75t_L g1250 ( 
.A(n_1056),
.Y(n_1250)
);

CKINVDCx10_ASAP7_75t_R g1251 ( 
.A(n_1071),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1037),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1252)
);

NOR3xp33_ASAP7_75t_L g1253 ( 
.A(n_1043),
.B(n_76),
.C(n_77),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1030),
.Y(n_1254)
);

OR2x6_ASAP7_75t_SL g1255 ( 
.A(n_1050),
.B(n_77),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_976),
.B(n_78),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1038),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1109),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_977),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_962),
.B(n_1091),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1092),
.B(n_82),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1040),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_991),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1084),
.Y(n_1264)
);

BUFx2_ASAP7_75t_SL g1265 ( 
.A(n_1110),
.Y(n_1265)
);

NAND2x1_ASAP7_75t_L g1266 ( 
.A(n_1084),
.B(n_303),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1045),
.B(n_86),
.Y(n_1267)
);

AND2x6_ASAP7_75t_L g1268 ( 
.A(n_1066),
.B(n_304),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1093),
.B(n_87),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1094),
.A2(n_1097),
.B(n_1095),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1072),
.A2(n_90),
.B1(n_87),
.B2(n_88),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_977),
.A2(n_91),
.B(n_88),
.C(n_90),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_988),
.B(n_961),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1051),
.A2(n_1114),
.B1(n_1118),
.B2(n_1113),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1119),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_987),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_983),
.A2(n_310),
.B(n_309),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1100),
.A2(n_100),
.B(n_96),
.C(n_98),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1070),
.B(n_96),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1101),
.A2(n_107),
.B1(n_104),
.B2(n_106),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1121),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1055),
.B(n_106),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1079),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_986),
.A2(n_313),
.B(n_311),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1052),
.B(n_111),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_989),
.A2(n_316),
.B(n_314),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_981),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1108),
.B(n_112),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_949),
.B(n_956),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1115),
.B(n_116),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1116),
.B(n_118),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1120),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1116),
.B(n_1117),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_960),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1117),
.B(n_119),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1107),
.A2(n_123),
.B(n_120),
.C(n_122),
.Y(n_1296)
);

BUFx8_ASAP7_75t_L g1297 ( 
.A(n_984),
.Y(n_1297)
);

OAI21xp33_ASAP7_75t_L g1298 ( 
.A1(n_1098),
.A2(n_124),
.B(n_125),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1013),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1002),
.B(n_127),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1122),
.A2(n_131),
.B1(n_128),
.B2(n_130),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_R g1302 ( 
.A(n_1035),
.B(n_130),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_L g1303 ( 
.A(n_946),
.B(n_338),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1096),
.A2(n_1099),
.B1(n_1106),
.B2(n_1105),
.Y(n_1304)
);

OR2x6_ASAP7_75t_SL g1305 ( 
.A(n_1010),
.B(n_135),
.Y(n_1305)
);

NOR3xp33_ASAP7_75t_L g1306 ( 
.A(n_1057),
.B(n_136),
.C(n_137),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_940),
.A2(n_348),
.B(n_347),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_992),
.B(n_139),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1082),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_965),
.B(n_139),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1003),
.A2(n_140),
.B(n_141),
.C(n_142),
.Y(n_1311)
);

NOR2x1_ASAP7_75t_L g1312 ( 
.A(n_935),
.B(n_143),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_935),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1138),
.A2(n_1237),
.A3(n_1140),
.B(n_1166),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1126),
.A2(n_146),
.A3(n_147),
.B(n_149),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1137),
.B(n_150),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1148),
.B(n_152),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1192),
.B(n_152),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1144),
.A2(n_1260),
.B(n_1217),
.Y(n_1319)
);

NOR2xp67_ASAP7_75t_L g1320 ( 
.A(n_1159),
.B(n_153),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1235),
.B(n_153),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1136),
.B(n_154),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1147),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1191),
.A2(n_155),
.A3(n_159),
.B(n_160),
.Y(n_1324)
);

AO21x2_ASAP7_75t_L g1325 ( 
.A1(n_1307),
.A2(n_363),
.B(n_362),
.Y(n_1325)
);

NOR2x1_ASAP7_75t_L g1326 ( 
.A(n_1178),
.B(n_161),
.Y(n_1326)
);

AO22x1_ASAP7_75t_L g1327 ( 
.A1(n_1128),
.A2(n_163),
.B1(n_166),
.B2(n_168),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1160),
.A2(n_1225),
.B(n_1193),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1224),
.Y(n_1329)
);

OAI22x1_ASAP7_75t_L g1330 ( 
.A1(n_1131),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1153),
.B(n_172),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1238),
.A2(n_179),
.A3(n_180),
.B(n_182),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1297),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_1167),
.Y(n_1334)
);

AND2x6_ASAP7_75t_SL g1335 ( 
.A(n_1178),
.B(n_183),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1297),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1238),
.A2(n_184),
.A3(n_185),
.B(n_186),
.Y(n_1337)
);

AOI211x1_ASAP7_75t_L g1338 ( 
.A1(n_1225),
.A2(n_184),
.B(n_185),
.C(n_187),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1136),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1184),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1147),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1146),
.B(n_191),
.Y(n_1342)
);

OAI21xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1178),
.A2(n_192),
.B(n_194),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1125),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1305),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1308),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1313),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1128),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1240),
.B(n_197),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1152),
.B(n_198),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1160),
.A2(n_199),
.B(n_200),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1134),
.B(n_203),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1274),
.A2(n_203),
.B(n_204),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1187),
.A2(n_204),
.A3(n_206),
.B(n_207),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1281),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1274),
.A2(n_1156),
.B(n_1270),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1189),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1229),
.A2(n_1228),
.A3(n_1185),
.B(n_1190),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1263),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1155),
.B(n_209),
.Y(n_1360)
);

INVx8_ASAP7_75t_L g1361 ( 
.A(n_1169),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1185),
.A2(n_211),
.B(n_212),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1159),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1293),
.B(n_213),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1188),
.B(n_213),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1174),
.A2(n_214),
.A3(n_217),
.B(n_219),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1254),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1172),
.B(n_221),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1130),
.A2(n_223),
.B(n_226),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1292),
.B(n_1151),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1142),
.A2(n_228),
.B(n_229),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1129),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1158),
.B(n_230),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1143),
.B(n_235),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1154),
.A2(n_235),
.B(n_236),
.Y(n_1375)
);

OAI22x1_ASAP7_75t_L g1376 ( 
.A1(n_1300),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1219),
.B(n_239),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1221),
.B(n_1223),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1232),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1145),
.B(n_243),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1235),
.B(n_245),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1179),
.A2(n_251),
.B(n_253),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_R g1383 ( 
.A(n_1239),
.B(n_255),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1242),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1181),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1194),
.A2(n_1197),
.B(n_1207),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1277),
.A2(n_1286),
.B(n_1284),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1202),
.Y(n_1388)
);

BUFx4f_ASAP7_75t_L g1389 ( 
.A(n_1209),
.Y(n_1389)
);

AO31x2_ASAP7_75t_L g1390 ( 
.A1(n_1259),
.A2(n_1276),
.A3(n_1272),
.B(n_1205),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1310),
.B(n_1164),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1288),
.B(n_1203),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1204),
.B(n_1227),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1226),
.B(n_1211),
.Y(n_1394)
);

O2A1O1Ixp5_ASAP7_75t_L g1395 ( 
.A1(n_1171),
.A2(n_1256),
.B(n_1241),
.C(n_1285),
.Y(n_1395)
);

NOR2xp67_ASAP7_75t_SL g1396 ( 
.A(n_1181),
.B(n_1183),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1289),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1247),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1173),
.A2(n_1165),
.B(n_1213),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1200),
.A2(n_1177),
.B1(n_1176),
.B2(n_1210),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1168),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1299),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1218),
.B(n_1279),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1161),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1287),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1282),
.A2(n_1150),
.B(n_1157),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1216),
.B(n_1290),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1186),
.B(n_1273),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1291),
.B(n_1295),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1246),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1311),
.A2(n_1233),
.B(n_1278),
.C(n_1220),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1267),
.A2(n_1195),
.B1(n_1199),
.B2(n_1253),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1261),
.B(n_1269),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1198),
.B(n_1214),
.Y(n_1414)
);

INVxp67_ASAP7_75t_SL g1415 ( 
.A(n_1186),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1273),
.B(n_1294),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1149),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1231),
.A2(n_1249),
.B1(n_1230),
.B2(n_1248),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1273),
.B(n_1312),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_L g1420 ( 
.A(n_1306),
.B(n_1296),
.C(n_1222),
.Y(n_1420)
);

NOR4xp25_ASAP7_75t_L g1421 ( 
.A(n_1244),
.B(n_1252),
.C(n_1246),
.D(n_1257),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1127),
.B(n_1309),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1206),
.Y(n_1423)
);

AO21x1_ASAP7_75t_L g1424 ( 
.A1(n_1303),
.A2(n_1244),
.B(n_1257),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1170),
.B(n_1304),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1206),
.B(n_1302),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1247),
.B(n_1264),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1250),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1162),
.B(n_1301),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1234),
.A2(n_1275),
.B(n_1283),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1215),
.A2(n_1301),
.B1(n_1252),
.B2(n_1262),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1275),
.A2(n_1271),
.B(n_1268),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1250),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1255),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1262),
.A2(n_1139),
.B1(n_1175),
.B2(n_1280),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1265),
.B(n_1258),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1208),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1245),
.Y(n_1438)
);

AND3x2_ASAP7_75t_L g1439 ( 
.A(n_1251),
.B(n_842),
.C(n_1060),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_SL g1440 ( 
.A1(n_1268),
.A2(n_1178),
.B(n_1185),
.Y(n_1440)
);

AO32x2_ASAP7_75t_L g1441 ( 
.A1(n_1275),
.A2(n_1244),
.A3(n_1185),
.B1(n_1252),
.B2(n_1246),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1133),
.A2(n_1141),
.B(n_1126),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1133),
.A2(n_1141),
.B(n_1126),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1148),
.B(n_832),
.Y(n_1444)
);

CKINVDCx6p67_ASAP7_75t_R g1445 ( 
.A(n_1125),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1148),
.B(n_851),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1184),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1243),
.A2(n_1217),
.B(n_1132),
.C(n_1260),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1128),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1126),
.A2(n_1133),
.B(n_964),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1153),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1148),
.A2(n_1238),
.B1(n_1111),
.B2(n_1274),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1133),
.A2(n_1212),
.B(n_1201),
.Y(n_1455)
);

AOI221x1_ASAP7_75t_L g1456 ( 
.A1(n_1133),
.A2(n_1298),
.B1(n_1236),
.B2(n_1138),
.C(n_1135),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1134),
.Y(n_1457)
);

AO32x2_ASAP7_75t_L g1458 ( 
.A1(n_1275),
.A2(n_1244),
.A3(n_1185),
.B1(n_1252),
.B2(n_1246),
.Y(n_1458)
);

NAND3xp33_ASAP7_75t_SL g1459 ( 
.A(n_1163),
.B(n_892),
.C(n_872),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1136),
.B(n_1129),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1196),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1126),
.A2(n_1133),
.B(n_964),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1133),
.A2(n_1212),
.B(n_1201),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1178),
.A2(n_1185),
.B(n_1274),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1148),
.B(n_851),
.Y(n_1468)
);

NAND3x1_ASAP7_75t_L g1469 ( 
.A(n_1164),
.B(n_1004),
.C(n_1060),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1470)
);

NOR2xp67_ASAP7_75t_SL g1471 ( 
.A(n_1169),
.B(n_935),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1196),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1196),
.Y(n_1473)
);

AOI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1132),
.A2(n_1182),
.B(n_1238),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1138),
.A2(n_1089),
.B(n_940),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1148),
.A2(n_1238),
.B1(n_1111),
.B2(n_1274),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1133),
.A2(n_1212),
.B(n_1201),
.Y(n_1477)
);

NOR2x1_ASAP7_75t_SL g1478 ( 
.A(n_1178),
.B(n_1169),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1297),
.Y(n_1480)
);

AOI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1141),
.A2(n_1133),
.B(n_1126),
.Y(n_1481)
);

NAND3x1_ASAP7_75t_L g1482 ( 
.A(n_1164),
.B(n_1004),
.C(n_1060),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1153),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1147),
.Y(n_1485)
);

NAND2xp33_ASAP7_75t_L g1486 ( 
.A(n_1169),
.B(n_1083),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1243),
.A2(n_1217),
.B(n_1132),
.C(n_1260),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1297),
.Y(n_1489)
);

OAI22x1_ASAP7_75t_L g1490 ( 
.A1(n_1131),
.A2(n_674),
.B1(n_919),
.B2(n_827),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1135),
.B(n_1182),
.C(n_1230),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1297),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1137),
.B(n_942),
.Y(n_1493)
);

A2O1A1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1243),
.A2(n_1217),
.B(n_1132),
.C(n_1260),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1148),
.A2(n_1238),
.B1(n_1111),
.B2(n_1274),
.Y(n_1495)
);

O2A1O1Ixp5_ASAP7_75t_L g1496 ( 
.A1(n_1180),
.A2(n_1171),
.B(n_1193),
.C(n_1133),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1148),
.B(n_832),
.Y(n_1497)
);

AOI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1141),
.A2(n_1133),
.B(n_1126),
.Y(n_1498)
);

O2A1O1Ixp33_ASAP7_75t_SL g1499 ( 
.A1(n_1266),
.A2(n_985),
.B(n_1166),
.C(n_1191),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1184),
.Y(n_1500)
);

NAND3x1_ASAP7_75t_L g1501 ( 
.A(n_1164),
.B(n_1004),
.C(n_1060),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1184),
.Y(n_1502)
);

OA22x2_ASAP7_75t_L g1503 ( 
.A1(n_1178),
.A2(n_1063),
.B1(n_914),
.B2(n_827),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1148),
.B(n_832),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1196),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1153),
.B(n_832),
.Y(n_1506)
);

AO21x2_ASAP7_75t_L g1507 ( 
.A1(n_1133),
.A2(n_1212),
.B(n_1201),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1297),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1196),
.Y(n_1509)
);

O2A1O1Ixp5_ASAP7_75t_L g1510 ( 
.A1(n_1180),
.A2(n_1171),
.B(n_1193),
.C(n_1133),
.Y(n_1510)
);

NOR3xp33_ASAP7_75t_SL g1511 ( 
.A(n_1239),
.B(n_892),
.C(n_847),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1137),
.B(n_942),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1153),
.B(n_832),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1297),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1196),
.Y(n_1516)
);

OAI22x1_ASAP7_75t_L g1517 ( 
.A1(n_1131),
.A2(n_674),
.B1(n_919),
.B2(n_827),
.Y(n_1517)
);

INVx8_ASAP7_75t_L g1518 ( 
.A(n_1178),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1243),
.A2(n_1217),
.B(n_1132),
.C(n_1260),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1196),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1148),
.B(n_1192),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1163),
.A2(n_827),
.B(n_1164),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1125),
.Y(n_1523)
);

AOI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1141),
.A2(n_1133),
.B(n_1126),
.Y(n_1524)
);

BUFx2_ASAP7_75t_R g1525 ( 
.A(n_1348),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1456),
.A2(n_1443),
.B(n_1442),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1336),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1493),
.B(n_1512),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1431),
.A2(n_1503),
.B1(n_1429),
.B2(n_1391),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1340),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1480),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1519),
.A2(n_1328),
.B(n_1356),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1357),
.Y(n_1533)
);

INVx8_ASAP7_75t_L g1534 ( 
.A(n_1361),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1489),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1319),
.A2(n_1464),
.B(n_1450),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1449),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1447),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1361),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1492),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1500),
.Y(n_1541)
);

AO31x2_ASAP7_75t_L g1542 ( 
.A1(n_1453),
.A2(n_1476),
.A3(n_1495),
.B(n_1438),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1518),
.B(n_1361),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1444),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_R g1545 ( 
.A(n_1508),
.B(n_1428),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1502),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1461),
.B(n_1457),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1524),
.A2(n_1498),
.B(n_1481),
.Y(n_1548)
);

INVx2_ASAP7_75t_SL g1549 ( 
.A(n_1389),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1329),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1506),
.B(n_1514),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1495),
.A2(n_1387),
.B(n_1475),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1462),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1472),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1503),
.A2(n_1410),
.B1(n_1424),
.B2(n_1394),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1394),
.A2(n_1406),
.B1(n_1418),
.B2(n_1322),
.Y(n_1556)
);

AO21x1_ASAP7_75t_L g1557 ( 
.A1(n_1432),
.A2(n_1435),
.B(n_1362),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1496),
.A2(n_1510),
.B(n_1474),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_SL g1559 ( 
.A1(n_1478),
.A2(n_1362),
.B(n_1351),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1460),
.B(n_1463),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1473),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1505),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1460),
.B(n_1463),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1509),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1467),
.B(n_1470),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1470),
.B(n_1479),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1516),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_1363),
.B(n_1333),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1406),
.A2(n_1418),
.B1(n_1430),
.B2(n_1316),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1491),
.A2(n_1432),
.B(n_1399),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1479),
.B(n_1483),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1404),
.Y(n_1572)
);

NOR2xp67_ASAP7_75t_L g1573 ( 
.A(n_1515),
.B(n_1417),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1520),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1483),
.B(n_1487),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1404),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1518),
.B(n_1440),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1513),
.B(n_1521),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1402),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1345),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1396),
.B(n_1389),
.Y(n_1581)
);

BUFx8_ASAP7_75t_SL g1582 ( 
.A(n_1355),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1398),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1403),
.A2(n_1491),
.B(n_1370),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1497),
.B(n_1504),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1386),
.A2(n_1409),
.B(n_1393),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1452),
.B(n_1484),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1518),
.B(n_1466),
.Y(n_1588)
);

BUFx8_ASAP7_75t_L g1589 ( 
.A(n_1433),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1409),
.A2(n_1393),
.B(n_1413),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1372),
.B(n_1377),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1384),
.Y(n_1592)
);

A2O1A1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1411),
.A2(n_1522),
.B(n_1430),
.C(n_1392),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1413),
.A2(n_1403),
.B(n_1499),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1415),
.B(n_1419),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1445),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1455),
.A2(n_1477),
.B(n_1465),
.Y(n_1597)
);

NOR2xp67_ASAP7_75t_L g1598 ( 
.A(n_1388),
.B(n_1423),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1359),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1367),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1522),
.B(n_1400),
.Y(n_1601)
);

BUFx2_ASAP7_75t_SL g1602 ( 
.A(n_1401),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1405),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1378),
.Y(n_1604)
);

INVx6_ASAP7_75t_L g1605 ( 
.A(n_1436),
.Y(n_1605)
);

NOR2x1_ASAP7_75t_SL g1606 ( 
.A(n_1436),
.B(n_1334),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1353),
.A2(n_1350),
.B(n_1395),
.C(n_1346),
.Y(n_1607)
);

BUFx4f_ASAP7_75t_L g1608 ( 
.A(n_1321),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1360),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1365),
.B(n_1321),
.Y(n_1610)
);

BUFx2_ASAP7_75t_R g1611 ( 
.A(n_1434),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1344),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1347),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1318),
.B(n_1421),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1381),
.B(n_1349),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1422),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1317),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1459),
.B(n_1414),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1317),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1318),
.B(n_1421),
.Y(n_1620)
);

CKINVDCx11_ASAP7_75t_R g1621 ( 
.A(n_1335),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1422),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1385),
.B(n_1523),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1364),
.A2(n_1420),
.B(n_1368),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1408),
.B(n_1426),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1352),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1381),
.B(n_1416),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1339),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1376),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1507),
.A2(n_1407),
.B(n_1486),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1407),
.B(n_1380),
.Y(n_1631)
);

AO21x2_ASAP7_75t_L g1632 ( 
.A1(n_1325),
.A2(n_1425),
.B(n_1420),
.Y(n_1632)
);

NOR2xp67_ASAP7_75t_L g1633 ( 
.A(n_1490),
.B(n_1517),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1326),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1379),
.Y(n_1635)
);

BUFx8_ASAP7_75t_L g1636 ( 
.A(n_1441),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1331),
.B(n_1441),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1368),
.A2(n_1342),
.B(n_1380),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1374),
.A2(n_1446),
.B(n_1468),
.Y(n_1639)
);

AOI22x1_ASAP7_75t_L g1640 ( 
.A1(n_1369),
.A2(n_1375),
.B1(n_1371),
.B2(n_1382),
.Y(n_1640)
);

AND2x6_ASAP7_75t_L g1641 ( 
.A(n_1323),
.B(n_1485),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1469),
.A2(n_1501),
.B(n_1482),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1383),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1427),
.B(n_1320),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1343),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1412),
.B(n_1358),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1330),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1366),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1366),
.Y(n_1649)
);

BUFx12f_ASAP7_75t_L g1650 ( 
.A(n_1397),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1358),
.B(n_1373),
.Y(n_1651)
);

INVxp67_ASAP7_75t_SL g1652 ( 
.A(n_1437),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1358),
.B(n_1390),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1441),
.B(n_1458),
.Y(n_1654)
);

INVx6_ASAP7_75t_L g1655 ( 
.A(n_1397),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1390),
.B(n_1314),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1332),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1332),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1327),
.B(n_1337),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1332),
.B(n_1337),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1439),
.B(n_1341),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1315),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1511),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1337),
.A2(n_1315),
.B(n_1338),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1458),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1324),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1354),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1354),
.A2(n_1488),
.B(n_1448),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1361),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1431),
.A2(n_1004),
.B1(n_1476),
.B2(n_1453),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1493),
.B(n_942),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1672)
);

OR2x6_ASAP7_75t_L g1673 ( 
.A(n_1518),
.B(n_1361),
.Y(n_1673)
);

BUFx2_ASAP7_75t_R g1674 ( 
.A(n_1348),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1319),
.A2(n_1133),
.B(n_1450),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1448),
.A2(n_1494),
.B(n_1488),
.Y(n_1676)
);

NAND2x1p5_ASAP7_75t_L g1677 ( 
.A(n_1471),
.B(n_1169),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1448),
.A2(n_1494),
.B(n_1488),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1448),
.A2(n_1494),
.B(n_1488),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1493),
.B(n_942),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1448),
.A2(n_1494),
.B(n_1488),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1448),
.A2(n_1494),
.B(n_1488),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1361),
.Y(n_1683)
);

INVx4_ASAP7_75t_L g1684 ( 
.A(n_1361),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1336),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1361),
.Y(n_1686)
);

NAND2x1p5_ASAP7_75t_L g1687 ( 
.A(n_1471),
.B(n_1169),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1577),
.B(n_1588),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1571),
.B(n_1575),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1534),
.Y(n_1690)
);

AO21x2_ASAP7_75t_L g1691 ( 
.A1(n_1558),
.A2(n_1668),
.B(n_1676),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1600),
.Y(n_1692)
);

AO21x2_ASAP7_75t_L g1693 ( 
.A1(n_1558),
.A2(n_1668),
.B(n_1676),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1603),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1550),
.Y(n_1695)
);

INVx5_ASAP7_75t_SL g1696 ( 
.A(n_1543),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1562),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1564),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1574),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1553),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1528),
.A2(n_1670),
.B1(n_1601),
.B2(n_1529),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1554),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1613),
.Y(n_1703)
);

OA21x2_ASAP7_75t_L g1704 ( 
.A1(n_1548),
.A2(n_1536),
.B(n_1678),
.Y(n_1704)
);

INVxp67_ASAP7_75t_L g1705 ( 
.A(n_1613),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1561),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1684),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1567),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1534),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1534),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1527),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1592),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1560),
.B(n_1565),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1616),
.Y(n_1714)
);

BUFx8_ASAP7_75t_SL g1715 ( 
.A(n_1582),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1576),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1530),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1576),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1533),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1684),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1563),
.B(n_1566),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1539),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1539),
.Y(n_1723)
);

OA21x2_ASAP7_75t_L g1724 ( 
.A1(n_1536),
.A2(n_1679),
.B(n_1678),
.Y(n_1724)
);

NAND2x1_ASAP7_75t_L g1725 ( 
.A(n_1559),
.B(n_1588),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1578),
.B(n_1622),
.Y(n_1726)
);

OA21x2_ASAP7_75t_L g1727 ( 
.A1(n_1679),
.A2(n_1682),
.B(n_1681),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1681),
.A2(n_1682),
.B(n_1675),
.Y(n_1728)
);

BUFx8_ASAP7_75t_SL g1729 ( 
.A(n_1537),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1538),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1671),
.B(n_1680),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1541),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1546),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1579),
.Y(n_1734)
);

INVx5_ASAP7_75t_L g1735 ( 
.A(n_1543),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1608),
.A2(n_1670),
.B1(n_1556),
.B2(n_1569),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_SL g1737 ( 
.A(n_1599),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1563),
.B(n_1566),
.Y(n_1738)
);

BUFx4f_ASAP7_75t_SL g1739 ( 
.A(n_1589),
.Y(n_1739)
);

AO21x2_ASAP7_75t_L g1740 ( 
.A1(n_1552),
.A2(n_1532),
.B(n_1675),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1669),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1652),
.Y(n_1742)
);

AO21x2_ASAP7_75t_L g1743 ( 
.A1(n_1552),
.A2(n_1532),
.B(n_1597),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1669),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1672),
.B(n_1604),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1652),
.Y(n_1746)
);

BUFx4f_ASAP7_75t_SL g1747 ( 
.A(n_1589),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1547),
.B(n_1614),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1593),
.B(n_1590),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1590),
.B(n_1654),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1526),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1587),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1551),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1629),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1647),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1556),
.B(n_1555),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1544),
.Y(n_1757)
);

INVxp67_ASAP7_75t_SL g1758 ( 
.A(n_1608),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1544),
.B(n_1586),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1644),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1636),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1644),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1543),
.Y(n_1763)
);

BUFx4f_ASAP7_75t_SL g1764 ( 
.A(n_1540),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1555),
.B(n_1617),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1623),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1644),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1633),
.A2(n_1628),
.B1(n_1569),
.B2(n_1557),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1612),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1614),
.B(n_1620),
.Y(n_1770)
);

OAI21xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1577),
.A2(n_1588),
.B(n_1631),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1683),
.Y(n_1772)
);

OR2x6_ASAP7_75t_L g1773 ( 
.A(n_1577),
.B(n_1673),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1634),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1662),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1619),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1631),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1586),
.B(n_1665),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1581),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1673),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1581),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1683),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1641),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1591),
.B(n_1620),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1627),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1637),
.B(n_1609),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1585),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1585),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1572),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1764),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1738),
.B(n_1635),
.Y(n_1791)
);

OR2x2_ASAP7_75t_SL g1792 ( 
.A(n_1783),
.B(n_1659),
.Y(n_1792)
);

OAI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1701),
.A2(n_1642),
.B1(n_1731),
.B2(n_1768),
.C(n_1736),
.Y(n_1793)
);

BUFx2_ASAP7_75t_L g1794 ( 
.A(n_1742),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1692),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1731),
.B(n_1689),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1694),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1738),
.B(n_1642),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1745),
.B(n_1610),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1748),
.B(n_1784),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1750),
.B(n_1542),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1695),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1697),
.Y(n_1803)
);

INVx4_ASAP7_75t_R g1804 ( 
.A(n_1739),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1769),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1786),
.B(n_1542),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1748),
.B(n_1646),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1688),
.B(n_1646),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1726),
.B(n_1667),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1726),
.B(n_1666),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1727),
.B(n_1657),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1745),
.B(n_1615),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1727),
.B(n_1658),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1759),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1721),
.B(n_1636),
.Y(n_1815)
);

INVx11_ASAP7_75t_L g1816 ( 
.A(n_1747),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1778),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1727),
.B(n_1648),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1770),
.B(n_1653),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1775),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1742),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1716),
.B(n_1718),
.Y(n_1822)
);

AND2x4_ASAP7_75t_SL g1823 ( 
.A(n_1773),
.B(n_1673),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1766),
.Y(n_1824)
);

INVx2_ASAP7_75t_SL g1825 ( 
.A(n_1735),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1711),
.Y(n_1826)
);

NOR4xp25_ASAP7_75t_SL g1827 ( 
.A(n_1760),
.B(n_1580),
.C(n_1645),
.D(n_1663),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1698),
.Y(n_1828)
);

OR2x2_ASAP7_75t_SL g1829 ( 
.A(n_1783),
.B(n_1605),
.Y(n_1829)
);

AND2x2_ASAP7_75t_SL g1830 ( 
.A(n_1688),
.B(n_1660),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1699),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1757),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1749),
.B(n_1649),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1717),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1787),
.B(n_1638),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1719),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1756),
.B(n_1656),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1775),
.Y(n_1838)
);

INVx4_ASAP7_75t_L g1839 ( 
.A(n_1735),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1756),
.B(n_1651),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1713),
.B(n_1651),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1788),
.B(n_1638),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1751),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1773),
.B(n_1630),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1713),
.B(n_1632),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1730),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1737),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1714),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1691),
.B(n_1664),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1691),
.B(n_1664),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1732),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1693),
.B(n_1570),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1746),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1693),
.B(n_1765),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1693),
.B(n_1570),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1773),
.B(n_1606),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1765),
.B(n_1584),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1690),
.Y(n_1858)
);

AOI33xp33_ASAP7_75t_L g1859 ( 
.A1(n_1755),
.A2(n_1626),
.A3(n_1583),
.B1(n_1625),
.B2(n_1549),
.B3(n_1595),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1794),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1859),
.B(n_1771),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1817),
.B(n_1728),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1796),
.B(n_1621),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1794),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1817),
.B(n_1728),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1840),
.B(n_1728),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1843),
.Y(n_1867)
);

NAND2x1p5_ASAP7_75t_L g1868 ( 
.A(n_1839),
.B(n_1856),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1840),
.B(n_1754),
.Y(n_1869)
);

OR2x6_ASAP7_75t_L g1870 ( 
.A(n_1844),
.B(n_1725),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1816),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1856),
.B(n_1707),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1837),
.B(n_1724),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1814),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1837),
.B(n_1845),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1821),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1845),
.B(n_1841),
.Y(n_1877)
);

AND2x4_ASAP7_75t_SL g1878 ( 
.A(n_1856),
.B(n_1773),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1841),
.B(n_1740),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1814),
.Y(n_1880)
);

NAND2x1p5_ASAP7_75t_L g1881 ( 
.A(n_1839),
.B(n_1725),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1854),
.B(n_1740),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1821),
.Y(n_1883)
);

INVx2_ASAP7_75t_SL g1884 ( 
.A(n_1853),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1857),
.B(n_1718),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1854),
.B(n_1740),
.Y(n_1886)
);

NOR3xp33_ASAP7_75t_L g1887 ( 
.A(n_1793),
.B(n_1618),
.C(n_1762),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1801),
.B(n_1743),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1801),
.B(n_1743),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1806),
.B(n_1743),
.Y(n_1890)
);

AND2x2_ASAP7_75t_SL g1891 ( 
.A(n_1830),
.B(n_1761),
.Y(n_1891)
);

CKINVDCx20_ASAP7_75t_R g1892 ( 
.A(n_1790),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1848),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1820),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1820),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1833),
.B(n_1704),
.Y(n_1896)
);

NOR2xp67_ASAP7_75t_L g1897 ( 
.A(n_1839),
.B(n_1767),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1838),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1800),
.B(n_1761),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1833),
.B(n_1704),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1853),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1857),
.B(n_1704),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1800),
.B(n_1777),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1807),
.B(n_1753),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1809),
.B(n_1810),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1826),
.B(n_1531),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1818),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1810),
.B(n_1811),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1905),
.B(n_1824),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1882),
.B(n_1813),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1861),
.A2(n_1607),
.B(n_1703),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1908),
.B(n_1849),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1894),
.Y(n_1913)
);

INVxp67_ASAP7_75t_L g1914 ( 
.A(n_1893),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1905),
.B(n_1832),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1894),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1908),
.B(n_1849),
.Y(n_1917)
);

NAND2x1_ASAP7_75t_SL g1918 ( 
.A(n_1897),
.B(n_1852),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_1864),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1873),
.B(n_1850),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1895),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1875),
.B(n_1795),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1873),
.B(n_1850),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1907),
.B(n_1807),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1879),
.B(n_1813),
.Y(n_1925)
);

INVxp67_ASAP7_75t_SL g1926 ( 
.A(n_1864),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1907),
.B(n_1819),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1895),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1879),
.B(n_1852),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1875),
.B(n_1797),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1898),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1867),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1868),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1882),
.B(n_1855),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1869),
.B(n_1802),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1886),
.B(n_1855),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1867),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1886),
.B(n_1808),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1870),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1874),
.Y(n_1940)
);

NAND2xp33_ASAP7_75t_R g1941 ( 
.A(n_1871),
.B(n_1545),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1874),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1909),
.B(n_1892),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1929),
.B(n_1877),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1912),
.B(n_1902),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1940),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1932),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1940),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1939),
.B(n_1870),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1932),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1929),
.B(n_1877),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1942),
.Y(n_1952)
);

INVx1_ASAP7_75t_SL g1953 ( 
.A(n_1915),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1912),
.B(n_1902),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1934),
.B(n_1890),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1942),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1910),
.B(n_1925),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1917),
.B(n_1896),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1917),
.B(n_1896),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1913),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1913),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1932),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1910),
.B(n_1885),
.Y(n_1963)
);

OAI21xp33_ASAP7_75t_L g1964 ( 
.A1(n_1934),
.A2(n_1887),
.B(n_1890),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1919),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1916),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1925),
.B(n_1885),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1916),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1936),
.B(n_1888),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1920),
.B(n_1900),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1921),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1921),
.Y(n_1972)
);

AND2x2_ASAP7_75t_SL g1973 ( 
.A(n_1939),
.B(n_1891),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1914),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1937),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1911),
.A2(n_1887),
.B1(n_1891),
.B2(n_1798),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1936),
.B(n_1888),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1928),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1952),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1952),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1965),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1957),
.B(n_1967),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1957),
.B(n_1922),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1956),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1949),
.B(n_1939),
.Y(n_1985)
);

OAI32xp33_ASAP7_75t_L g1986 ( 
.A1(n_1964),
.A2(n_1939),
.A3(n_1868),
.B1(n_1899),
.B2(n_1941),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1963),
.B(n_1920),
.Y(n_1987)
);

OAI22xp33_ASAP7_75t_L g1988 ( 
.A1(n_1976),
.A2(n_1933),
.B1(n_1868),
.B2(n_1897),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1973),
.B(n_1891),
.Y(n_1989)
);

OAI31xp33_ASAP7_75t_L g1990 ( 
.A1(n_1974),
.A2(n_1933),
.A3(n_1878),
.B(n_1823),
.Y(n_1990)
);

OAI32xp33_ASAP7_75t_L g1991 ( 
.A1(n_1953),
.A2(n_1899),
.A3(n_1906),
.B1(n_1881),
.B2(n_1924),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1973),
.A2(n_1911),
.B1(n_1938),
.B2(n_1930),
.Y(n_1992)
);

AOI21xp33_ASAP7_75t_SL g1993 ( 
.A1(n_1943),
.A2(n_1881),
.B(n_1847),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1963),
.B(n_1923),
.Y(n_1994)
);

OAI32xp33_ASAP7_75t_L g1995 ( 
.A1(n_1967),
.A2(n_1944),
.A3(n_1951),
.B1(n_1969),
.B2(n_1955),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1946),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1970),
.B(n_1923),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1947),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1956),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1949),
.A2(n_1938),
.B1(n_1889),
.B2(n_1830),
.Y(n_2000)
);

OAI33xp33_ASAP7_75t_L g2001 ( 
.A1(n_1977),
.A2(n_1935),
.A3(n_1805),
.B1(n_1869),
.B2(n_1752),
.B3(n_1903),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1961),
.Y(n_2002)
);

NAND4xp25_ASAP7_75t_L g2003 ( 
.A(n_1949),
.B(n_1863),
.C(n_1573),
.D(n_1643),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1970),
.B(n_1924),
.Y(n_2004)
);

OAI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1958),
.A2(n_1872),
.B(n_1926),
.Y(n_2005)
);

XNOR2xp5_ASAP7_75t_L g2006 ( 
.A(n_1958),
.B(n_1602),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1961),
.Y(n_2007)
);

OAI32xp33_ASAP7_75t_L g2008 ( 
.A1(n_1959),
.A2(n_1881),
.A3(n_1927),
.B1(n_1883),
.B2(n_1876),
.Y(n_2008)
);

INVxp67_ASAP7_75t_L g2009 ( 
.A(n_1948),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1966),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1966),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1985),
.B(n_1945),
.Y(n_2012)
);

AOI211xp5_ASAP7_75t_L g2013 ( 
.A1(n_1986),
.A2(n_1568),
.B(n_1661),
.C(n_1598),
.Y(n_2013)
);

AOI21xp33_ASAP7_75t_L g2014 ( 
.A1(n_1991),
.A2(n_1774),
.B(n_1705),
.Y(n_2014)
);

INVxp33_ASAP7_75t_L g2015 ( 
.A(n_2006),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1985),
.B(n_1945),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1990),
.B(n_1959),
.Y(n_2017)
);

OR2x2_ASAP7_75t_L g2018 ( 
.A(n_1987),
.B(n_1954),
.Y(n_2018)
);

AOI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1992),
.A2(n_1954),
.B1(n_1889),
.B2(n_1960),
.Y(n_2019)
);

O2A1O1Ixp33_ASAP7_75t_L g2020 ( 
.A1(n_1981),
.A2(n_1791),
.B(n_1842),
.C(n_1835),
.Y(n_2020)
);

O2A1O1Ixp33_ASAP7_75t_L g2021 ( 
.A1(n_2003),
.A2(n_1828),
.B(n_1831),
.C(n_1803),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1996),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1997),
.B(n_1900),
.Y(n_2023)
);

A2O1A1Ixp33_ASAP7_75t_L g2024 ( 
.A1(n_1993),
.A2(n_1823),
.B(n_1878),
.C(n_1918),
.Y(n_2024)
);

AOI221xp5_ASAP7_75t_L g2025 ( 
.A1(n_2001),
.A2(n_1972),
.B1(n_1971),
.B2(n_1978),
.C(n_1968),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_2001),
.A2(n_1968),
.B1(n_1978),
.B2(n_1927),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1989),
.A2(n_1860),
.B(n_1918),
.Y(n_2027)
);

OAI221xp5_ASAP7_75t_L g2028 ( 
.A1(n_2005),
.A2(n_1860),
.B1(n_1870),
.B2(n_1901),
.C(n_1884),
.Y(n_2028)
);

OAI322xp33_ASAP7_75t_L g2029 ( 
.A1(n_1982),
.A2(n_1904),
.A3(n_1903),
.B1(n_1815),
.B2(n_1866),
.C1(n_1884),
.C2(n_1822),
.Y(n_2029)
);

INVxp67_ASAP7_75t_L g2030 ( 
.A(n_1979),
.Y(n_2030)
);

OAI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_2027),
.A2(n_2005),
.B1(n_2000),
.B2(n_2009),
.C(n_1994),
.Y(n_2031)
);

AOI221xp5_ASAP7_75t_L g2032 ( 
.A1(n_2029),
.A2(n_1995),
.B1(n_2020),
.B2(n_2015),
.C(n_2017),
.Y(n_2032)
);

AOI221xp5_ASAP7_75t_L g2033 ( 
.A1(n_2022),
.A2(n_2008),
.B1(n_1988),
.B2(n_1994),
.C(n_1987),
.Y(n_2033)
);

AOI222xp33_ASAP7_75t_L g2034 ( 
.A1(n_2022),
.A2(n_1980),
.B1(n_2010),
.B2(n_2007),
.C1(n_2002),
.C2(n_1999),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_2021),
.A2(n_2011),
.B1(n_1984),
.B2(n_1998),
.C(n_1983),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_2013),
.A2(n_1878),
.B(n_2004),
.Y(n_2036)
);

AOI211xp5_ASAP7_75t_SL g2037 ( 
.A1(n_2028),
.A2(n_1720),
.B(n_1707),
.C(n_1804),
.Y(n_2037)
);

NAND4xp25_ASAP7_75t_L g2038 ( 
.A(n_2024),
.B(n_1685),
.C(n_1535),
.D(n_1596),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2014),
.A2(n_1690),
.B(n_1710),
.C(n_1709),
.Y(n_2039)
);

O2A1O1Ixp5_ASAP7_75t_L g2040 ( 
.A1(n_2012),
.A2(n_1880),
.B(n_1950),
.C(n_1947),
.Y(n_2040)
);

O2A1O1Ixp33_ASAP7_75t_L g2041 ( 
.A1(n_2030),
.A2(n_1707),
.B(n_1720),
.C(n_1779),
.Y(n_2041)
);

AOI221xp5_ASAP7_75t_L g2042 ( 
.A1(n_2025),
.A2(n_2030),
.B1(n_2019),
.B2(n_2026),
.C(n_2018),
.Y(n_2042)
);

OAI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_2016),
.A2(n_1901),
.B(n_1883),
.Y(n_2043)
);

OAI211xp5_ASAP7_75t_L g2044 ( 
.A1(n_2023),
.A2(n_1827),
.B(n_1710),
.C(n_1709),
.Y(n_2044)
);

AOI221xp5_ASAP7_75t_L g2045 ( 
.A1(n_2029),
.A2(n_1836),
.B1(n_1851),
.B2(n_1846),
.C(n_1834),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2026),
.B(n_1950),
.Y(n_2046)
);

O2A1O1Ixp5_ASAP7_75t_L g2047 ( 
.A1(n_2015),
.A2(n_1880),
.B(n_1975),
.C(n_1962),
.Y(n_2047)
);

OAI21xp33_ASAP7_75t_L g2048 ( 
.A1(n_2017),
.A2(n_1866),
.B(n_1865),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_2017),
.A2(n_1829),
.B1(n_1792),
.B2(n_1870),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_2022),
.Y(n_2050)
);

OAI211xp5_ASAP7_75t_SL g2051 ( 
.A1(n_2013),
.A2(n_1781),
.B(n_1904),
.C(n_1812),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2050),
.Y(n_2052)
);

NAND3xp33_ASAP7_75t_L g2053 ( 
.A(n_2032),
.B(n_1624),
.C(n_1789),
.Y(n_2053)
);

AOI211xp5_ASAP7_75t_SL g2054 ( 
.A1(n_2049),
.A2(n_1720),
.B(n_1816),
.C(n_1611),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_2038),
.B(n_1715),
.Y(n_2055)
);

NOR3xp33_ASAP7_75t_L g2056 ( 
.A(n_2042),
.B(n_1624),
.C(n_1758),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2043),
.B(n_1862),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_2033),
.B(n_1594),
.C(n_1584),
.Y(n_2058)
);

NAND5xp2_ASAP7_75t_L g2059 ( 
.A(n_2037),
.B(n_1715),
.C(n_1674),
.D(n_1525),
.E(n_1611),
.Y(n_2059)
);

NOR3xp33_ASAP7_75t_L g2060 ( 
.A(n_2048),
.B(n_1741),
.C(n_1722),
.Y(n_2060)
);

NOR4xp25_ASAP7_75t_L g2061 ( 
.A(n_2031),
.B(n_1733),
.C(n_1702),
.D(n_1706),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2045),
.B(n_1962),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_L g2063 ( 
.A(n_2041),
.B(n_1858),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2036),
.B(n_1862),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2035),
.B(n_2034),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2046),
.B(n_1975),
.Y(n_2066)
);

NAND3xp33_ASAP7_75t_L g2067 ( 
.A(n_2065),
.B(n_2052),
.C(n_2054),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2063),
.Y(n_2068)
);

NOR2xp33_ASAP7_75t_L g2069 ( 
.A(n_2055),
.B(n_1729),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2064),
.B(n_2039),
.Y(n_2070)
);

NAND3x1_ASAP7_75t_L g2071 ( 
.A(n_2056),
.B(n_2047),
.C(n_2040),
.Y(n_2071)
);

NOR3xp33_ASAP7_75t_L g2072 ( 
.A(n_2053),
.B(n_2044),
.C(n_2051),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_2059),
.B(n_1729),
.Y(n_2073)
);

NOR2xp67_ASAP7_75t_L g2074 ( 
.A(n_2062),
.B(n_1650),
.Y(n_2074)
);

NAND3xp33_ASAP7_75t_L g2075 ( 
.A(n_2054),
.B(n_1594),
.C(n_1640),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2061),
.B(n_1928),
.Y(n_2076)
);

NAND4xp75_ASAP7_75t_L g2077 ( 
.A(n_2066),
.B(n_1525),
.C(n_1674),
.D(n_1737),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2057),
.B(n_1931),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2058),
.Y(n_2079)
);

NOR2x1_ASAP7_75t_L g2080 ( 
.A(n_2060),
.B(n_1737),
.Y(n_2080)
);

OAI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_2067),
.A2(n_2072),
.B(n_2074),
.Y(n_2081)
);

INVxp33_ASAP7_75t_L g2082 ( 
.A(n_2069),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_2067),
.B(n_1655),
.Y(n_2083)
);

NOR4xp25_ASAP7_75t_L g2084 ( 
.A(n_2079),
.B(n_1780),
.C(n_1763),
.D(n_1708),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2076),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_2077),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_2073),
.B(n_1858),
.Y(n_2087)
);

NOR3xp33_ASAP7_75t_L g2088 ( 
.A(n_2068),
.B(n_1686),
.C(n_1722),
.Y(n_2088)
);

OAI221xp5_ASAP7_75t_L g2089 ( 
.A1(n_2080),
.A2(n_1780),
.B1(n_1763),
.B2(n_1870),
.C(n_1825),
.Y(n_2089)
);

NAND3xp33_ASAP7_75t_L g2090 ( 
.A(n_2070),
.B(n_1639),
.C(n_1700),
.Y(n_2090)
);

OAI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_2086),
.A2(n_2071),
.B1(n_2078),
.B2(n_2075),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_2087),
.Y(n_2092)
);

BUFx3_ASAP7_75t_L g2093 ( 
.A(n_2087),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_2083),
.Y(n_2094)
);

INVxp67_ASAP7_75t_L g2095 ( 
.A(n_2081),
.Y(n_2095)
);

NOR4xp25_ASAP7_75t_L g2096 ( 
.A(n_2085),
.B(n_1776),
.C(n_1712),
.D(n_1734),
.Y(n_2096)
);

XOR2x2_ASAP7_75t_L g2097 ( 
.A(n_2088),
.B(n_1799),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_2090),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2084),
.B(n_1884),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2097),
.Y(n_2100)
);

OAI22x1_ASAP7_75t_L g2101 ( 
.A1(n_2095),
.A2(n_2082),
.B1(n_2089),
.B2(n_1686),
.Y(n_2101)
);

OAI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2091),
.A2(n_1829),
.B1(n_1696),
.B2(n_1655),
.Y(n_2102)
);

XOR2xp5_ASAP7_75t_L g2103 ( 
.A(n_2094),
.B(n_1785),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_2092),
.Y(n_2104)
);

INVx4_ASAP7_75t_L g2105 ( 
.A(n_2093),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_2098),
.A2(n_1744),
.B(n_1723),
.Y(n_2106)
);

OAI22x1_ASAP7_75t_L g2107 ( 
.A1(n_2105),
.A2(n_2092),
.B1(n_2099),
.B2(n_2096),
.Y(n_2107)
);

OAI22x1_ASAP7_75t_L g2108 ( 
.A1(n_2104),
.A2(n_2096),
.B1(n_1677),
.B2(n_1687),
.Y(n_2108)
);

BUFx2_ASAP7_75t_L g2109 ( 
.A(n_2101),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2107),
.Y(n_2110)
);

AOI21xp33_ASAP7_75t_L g2111 ( 
.A1(n_2110),
.A2(n_2109),
.B(n_2100),
.Y(n_2111)
);

OAI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2111),
.A2(n_2102),
.B(n_2103),
.Y(n_2112)
);

OA21x2_ASAP7_75t_L g2113 ( 
.A1(n_2112),
.A2(n_2106),
.B(n_2108),
.Y(n_2113)
);

A2O1A1Ixp33_ASAP7_75t_L g2114 ( 
.A1(n_2113),
.A2(n_1782),
.B(n_1772),
.C(n_1723),
.Y(n_2114)
);


endmodule