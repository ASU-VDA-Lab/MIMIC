module fake_jpeg_8623_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_43),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_18),
.B1(n_40),
.B2(n_35),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_58),
.Y(n_75)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_69),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_8),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_30),
.B(n_27),
.C(n_31),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_67),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_18),
.B1(n_33),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_66),
.B1(n_33),
.B2(n_42),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_18),
.B1(n_33),
.B2(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_21),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_43),
.C(n_26),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_43),
.C(n_26),
.Y(n_112)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_25),
.B1(n_29),
.B2(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_33),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_21),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_88),
.B1(n_94),
.B2(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_31),
.Y(n_122)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_35),
.B1(n_40),
.B2(n_51),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_49),
.B(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_103),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_77),
.B(n_30),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_111),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_68),
.B1(n_51),
.B2(n_46),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_84),
.B1(n_75),
.B2(n_70),
.Y(n_133)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_26),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_113),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_22),
.B(n_21),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_88),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_118),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_30),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_119),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_123),
.B1(n_25),
.B2(n_29),
.Y(n_144)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_27),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_30),
.B(n_27),
.C(n_31),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_124),
.B(n_126),
.Y(n_154)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_86),
.B1(n_91),
.B2(n_46),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_138),
.B1(n_140),
.B2(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_137),
.B1(n_143),
.B2(n_149),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_75),
.B1(n_83),
.B2(n_70),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_79),
.B1(n_59),
.B2(n_90),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_59),
.B1(n_93),
.B2(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_83),
.B1(n_89),
.B2(n_55),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_38),
.B1(n_57),
.B2(n_45),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_36),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_148),
.B(n_141),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_104),
.A2(n_55),
.B1(n_74),
.B2(n_73),
.Y(n_149)
);

INVx2_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_98),
.B(n_119),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_158),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_153),
.A2(n_157),
.B(n_165),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_111),
.C(n_112),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_164),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_156),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_116),
.C(n_99),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_106),
.B1(n_103),
.B2(n_121),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_178),
.B1(n_163),
.B2(n_129),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_129),
.A2(n_96),
.B1(n_25),
.B2(n_29),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_170),
.B1(n_22),
.B2(n_149),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_72),
.B1(n_19),
.B2(n_27),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_97),
.B1(n_96),
.B2(n_101),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_0),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_147),
.B(n_22),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_32),
.A3(n_22),
.B1(n_16),
.B2(n_23),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

AOI32xp33_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_71),
.A3(n_52),
.B1(n_47),
.B2(n_72),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_24),
.B(n_23),
.C(n_16),
.D(n_41),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_178),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_71),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_181),
.B(n_185),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_145),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_146),
.B1(n_144),
.B2(n_166),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_183),
.A2(n_195),
.B1(n_202),
.B2(n_204),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_143),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_186),
.C(n_193),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_147),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_153),
.B(n_133),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_24),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_137),
.B1(n_127),
.B2(n_141),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_136),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_19),
.B(n_47),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_17),
.B(n_24),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_52),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_156),
.C(n_19),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_19),
.B1(n_64),
.B2(n_36),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_203),
.A2(n_168),
.B1(n_174),
.B2(n_171),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_165),
.B1(n_158),
.B2(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_212),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_224),
.B1(n_226),
.B2(n_229),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_162),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_171),
.C(n_167),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_222),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_12),
.C(n_14),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_215),
.B(n_221),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_160),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_223),
.C(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_156),
.Y(n_218)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_194),
.B(n_156),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_219),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_201),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_184),
.C(n_186),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_41),
.C(n_36),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_17),
.B(n_41),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_203),
.B1(n_200),
.B2(n_179),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_198),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_237),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_219),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_221),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_182),
.B1(n_205),
.B2(n_198),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_247),
.B1(n_228),
.B2(n_229),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_183),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_225),
.C(n_208),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_185),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_214),
.Y(n_257)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_206),
.B(n_193),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_41),
.B1(n_17),
.B2(n_23),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_248)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_257),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_232),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_267),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_217),
.C(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_261),
.C(n_1),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_227),
.C(n_207),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_10),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_245),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_247),
.Y(n_275)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_234),
.A3(n_246),
.B1(n_236),
.B2(n_239),
.C1(n_250),
.C2(n_242),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_238),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_17),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_7),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

AO221x1_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_241),
.B1(n_231),
.B2(n_232),
.C(n_237),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_259),
.B(n_11),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_285),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_14),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_284),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_0),
.B(n_1),
.Y(n_282)
);

OAI321xp33_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_12),
.A3(n_11),
.B1(n_8),
.B2(n_4),
.C(n_5),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_254),
.C(n_261),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_13),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_13),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_262),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_290),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_257),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_293),
.C(n_2),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_255),
.B1(n_259),
.B2(n_12),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_276),
.B(n_282),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_11),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_1),
.C(n_2),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_3),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_302),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_294),
.A2(n_274),
.B(n_272),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_305),
.C(n_308),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_272),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_298),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_8),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_307),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_1),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_292),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_310),
.C(n_313),
.Y(n_318)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_290),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_306),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_315),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_302),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_291),
.B(n_295),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_319),
.A2(n_311),
.B(n_3),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_3),
.C(n_5),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_321),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_318),
.Y(n_324)
);

OAI21xp33_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_323),
.B(n_317),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_6),
.B(n_309),
.Y(n_326)
);


endmodule