module real_jpeg_33149_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_0),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_0),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_0),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_0),
.Y(n_508)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_1),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_1),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_1),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_1),
.B(n_76),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_1),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_1),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_1),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_1),
.B(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_2),
.B(n_278),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_2),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_3),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_3),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_3),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_3),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_3),
.B(n_203),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g451 ( 
.A(n_3),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_3),
.B(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_4),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_6),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_7),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_7),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_7),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_7),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_7),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_SL g346 ( 
.A(n_7),
.B(n_347),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_7),
.B(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_8),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_9),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_9),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_9),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_9),
.B(n_152),
.Y(n_151)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_240),
.Y(n_239)
);

NAND2x1_ASAP7_75t_L g248 ( 
.A(n_9),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_9),
.B(n_116),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_10),
.B(n_44),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_10),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_10),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_10),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_10),
.B(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_SL g474 ( 
.A(n_10),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_10),
.B(n_489),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_11),
.Y(n_154)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_11),
.Y(n_205)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_13),
.Y(n_251)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_13),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_14),
.B(n_80),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_14),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_14),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_14),
.B(n_144),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_14),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_14),
.B(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_14),
.B(n_507),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_15),
.Y(n_162)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_15),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_36),
.Y(n_35)
);

AND2x4_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_16),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_16),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_16),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_16),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_16),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_17),
.B(n_51),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_17),
.B(n_189),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g319 ( 
.A(n_17),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_17),
.B(n_342),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_17),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_17),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_17),
.B(n_423),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_17),
.B(n_455),
.Y(n_454)
);

OAI311xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_175),
.A3(n_279),
.B1(n_283),
.C1(n_557),
.Y(n_18)
);

AOI331xp33_ASAP7_75t_L g283 ( 
.A1(n_19),
.A2(n_20),
.A3(n_176),
.B1(n_276),
.B2(n_284),
.B3(n_553),
.C1(n_554),
.Y(n_283)
);

NAND4xp25_ASAP7_75t_L g557 ( 
.A(n_19),
.B(n_276),
.C(n_279),
.D(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_173),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_22),
.B(n_102),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_82),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_46),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.C(n_42),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_35),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_36),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_37),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_37),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_38),
.B(n_91),
.C(n_95),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_38),
.A2(n_39),
.B1(n_95),
.B2(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_38),
.B(n_307),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_38),
.B(n_147),
.C(n_308),
.Y(n_375)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_40),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_41),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_43),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_47),
.B(n_137),
.C(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_47),
.B(n_228),
.Y(n_377)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_49),
.A2(n_50),
.B1(n_129),
.B2(n_139),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_49),
.A2(n_50),
.B1(n_141),
.B2(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_50),
.B(n_130),
.C(n_138),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_54),
.B(n_237),
.C(n_247),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_54),
.A2(n_55),
.B1(n_247),
.B2(n_248),
.Y(n_400)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_56),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g82 ( 
.A(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_75),
.C(n_77),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_60),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.C(n_70),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_61),
.A2(n_62),
.B1(n_68),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_68),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_68),
.A2(n_107),
.B1(n_201),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2x2_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_75),
.A2(n_88),
.B1(n_120),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_75),
.A2(n_88),
.B1(n_206),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_81),
.Y(n_231)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJx2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.C(n_99),
.Y(n_84)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_85),
.B(n_172),
.Y(n_171)
);

INVxp33_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_110),
.C(n_119),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_88),
.B(n_200),
.C(n_206),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_90),
.B(n_99),
.Y(n_172)
);

XOR2x2_ASAP7_75t_L g165 ( 
.A(n_91),
.B(n_166),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_93),
.B(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_111),
.C(n_158),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_95),
.B(n_316),
.Y(n_315)
);

MAJx2_ASAP7_75t_L g358 ( 
.A(n_95),
.B(n_316),
.C(n_319),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_96),
.Y(n_420)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_97),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_98),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_98),
.Y(n_503)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_163),
.C(n_170),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_103),
.B(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_126),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_264)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_107),
.B(n_201),
.C(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_110),
.B(n_209),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_117),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_112),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_111),
.A2(n_112),
.B1(n_117),
.B2(n_196),
.Y(n_195)
);

OAI221xp5_ASAP7_75t_L g197 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_117),
.C(n_196),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_112),
.B(n_243),
.Y(n_417)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_114),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_115),
.B(n_191),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_195),
.B(n_197),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_115),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_115),
.A2(n_223),
.B1(n_422),
.B2(n_459),
.Y(n_458)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_116),
.Y(n_336)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_125),
.Y(n_310)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_127),
.B(n_264),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_140),
.C(n_155),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_132),
.Y(n_322)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_137),
.B(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_139),
.B(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_141),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.C(n_150),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_146),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_148),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_147),
.A2(n_148),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_161),
.Y(n_292)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_164),
.B(n_171),
.Y(n_273)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_165),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_168),
.B(n_169),
.Y(n_267)
);

INVxp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_276),
.Y(n_176)
);

INVxp33_ASAP7_75t_SL g553 ( 
.A(n_177),
.Y(n_553)
);

OA21x2_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_268),
.B(n_274),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_258),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_179),
.B(n_258),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_212),
.C(n_218),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_181),
.B(n_213),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_198),
.Y(n_181)
);

INVxp33_ASAP7_75t_SL g260 ( 
.A(n_182),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_194),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_183),
.B(n_186),
.Y(n_531)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B(n_193),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_191),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_191),
.A2(n_225),
.B1(n_334),
.B2(n_337),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_191),
.B(n_337),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_192),
.Y(n_489)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_193),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_193),
.A2(n_296),
.B1(n_414),
.B2(n_415),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_194),
.B(n_531),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_207),
.B1(n_208),
.B2(n_211),
.Y(n_198)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_260),
.C(n_261),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_219),
.B(n_525),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_235),
.C(n_252),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_220),
.B(n_529),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.C(n_232),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_222),
.B(n_227),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_223),
.B(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_232),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_235),
.A2(n_236),
.B1(n_254),
.B2(n_255),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_237),
.A2(n_238),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.C(n_246),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_239),
.B(n_383),
.Y(n_382)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_243),
.B(n_246),
.Y(n_383)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_266),
.C(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_275),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g275 ( 
.A(n_272),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_277),
.B(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_284),
.Y(n_558)
);

OA21x2_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_522),
.B(n_546),
.Y(n_284)
);

NAND3xp33_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_386),
.C(n_406),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_360),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_287),
.B(n_360),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_312),
.C(n_338),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_288),
.B(n_313),
.Y(n_410)
);

XOR2x2_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_306),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_290),
.B(n_306),
.C(n_385),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_293),
.B(n_294),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_293),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_294),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_294),
.B(n_380),
.C(n_382),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_295),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.C(n_304),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_297),
.A2(n_298),
.B1(n_304),
.B2(n_305),
.Y(n_414)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_308),
.Y(n_311)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_323),
.C(n_333),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_314),
.B(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_318),
.B(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_323),
.B(n_333),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_329),
.C(n_330),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_325),
.B(n_331),
.Y(n_464)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_329),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_334),
.Y(n_337)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_338),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_340),
.B1(n_354),
.B2(n_359),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_355),
.C(n_358),
.Y(n_362)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_344),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_346),
.C(n_350),
.Y(n_380)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_350),
.B2(n_351),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_349),
.Y(n_453)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_354),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_378),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_379),
.C(n_384),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_364),
.C(n_376),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_376),
.Y(n_363)
);

XNOR2x2_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_375),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_371),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_SL g396 ( 
.A(n_366),
.B(n_371),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_371),
.Y(n_397)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_375),
.A2(n_396),
.B(n_397),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_384),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

AOI21x1_ASAP7_75t_L g547 ( 
.A1(n_387),
.A2(n_548),
.B(n_549),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_388),
.B(n_389),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_390),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_402),
.B2(n_403),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_392),
.Y(n_542)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_395),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_398),
.Y(n_536)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g534 ( 
.A(n_401),
.Y(n_534)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_403),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_431),
.B(n_521),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_408),
.B(n_411),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_416),
.B(n_425),
.C(n_428),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_412),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_413),
.A2(n_416),
.B1(n_429),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_413),
.Y(n_519)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_414),
.Y(n_415)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_416),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.C(n_421),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_417),
.A2(n_418),
.B1(n_419),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_421),
.B(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_422),
.Y(n_459)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_425),
.A2(n_426),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_513),
.B(n_520),
.Y(n_431)
);

OAI21xp33_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_470),
.B(n_512),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_460),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_434),
.B(n_460),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_450),
.C(n_457),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_435),
.A2(n_436),
.B1(n_482),
.B2(n_483),
.Y(n_481)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_444),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_439),
.B1(n_442),
.B2(n_443),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_443),
.C(n_444),
.Y(n_462)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_442),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_450),
.A2(n_457),
.B1(n_458),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_454),
.Y(n_473)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

BUFx4f_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_467),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_465),
.B2(n_466),
.Y(n_461)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_462),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_463),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_463),
.B(n_465),
.C(n_515),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_467),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_485),
.B(n_511),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_481),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_481),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.C(n_477),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_496),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_474),
.A2(n_477),
.B1(n_478),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_486),
.A2(n_498),
.B(n_510),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_495),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_487),
.B(n_495),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_490),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_490),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_488),
.B(n_506),
.Y(n_505)
);

INVx3_ASAP7_75t_SL g491 ( 
.A(n_492),
.Y(n_491)
);

INVx8_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_505),
.B(n_509),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_504),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_504),
.Y(n_509)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_516),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_516),
.Y(n_520)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_537),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_526),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_524),
.A2(n_526),
.B1(n_538),
.B2(n_540),
.Y(n_551)
);

NOR2x1_ASAP7_75t_SL g552 ( 
.A(n_524),
.B(n_526),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_530),
.C(n_532),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_530),
.Y(n_539)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_533),
.B(n_539),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_535),
.C(n_536),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_540),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_540),
.Y(n_550)
);

MAJx2_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_543),
.C(n_545),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

O2A1O1Ixp33_ASAP7_75t_SL g546 ( 
.A1(n_547),
.A2(n_550),
.B(n_551),
.C(n_552),
.Y(n_546)
);

INVx6_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);


endmodule