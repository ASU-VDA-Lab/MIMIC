module real_aes_508_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_0), .A2(n_115), .B1(n_414), .B2(n_567), .Y(n_566) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_1), .A2(n_65), .B1(n_217), .B2(n_251), .C1(n_285), .C2(n_288), .Y(n_323) );
OA22x2_ASAP7_75t_L g405 ( .A1(n_2), .A2(n_406), .B1(n_407), .B2(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_2), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_3), .A2(n_99), .B1(n_602), .B2(n_603), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_4), .A2(n_218), .B1(n_459), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_5), .A2(n_50), .B1(n_278), .B2(n_325), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_6), .A2(n_129), .B1(n_303), .B2(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g238 ( .A(n_7), .Y(n_238) );
AO22x2_ASAP7_75t_L g265 ( .A1(n_7), .A2(n_160), .B1(n_255), .B2(n_266), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_8), .A2(n_132), .B1(n_297), .B2(n_298), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_9), .A2(n_203), .B1(n_285), .B2(n_288), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_10), .A2(n_93), .B1(n_363), .B2(n_365), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_11), .A2(n_131), .B1(n_385), .B2(n_451), .Y(n_491) );
XOR2x2_ASAP7_75t_L g469 ( .A(n_12), .B(n_470), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_13), .A2(n_94), .B1(n_305), .B2(n_306), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_14), .A2(n_159), .B1(n_269), .B2(n_273), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_15), .A2(n_77), .B1(n_389), .B2(n_392), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_16), .A2(n_90), .B1(n_422), .B2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_17), .A2(n_27), .B1(n_278), .B2(n_325), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_18), .A2(n_97), .B1(n_453), .B2(n_455), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_19), .B(n_237), .Y(n_236) );
AO22x2_ASAP7_75t_L g262 ( .A1(n_19), .A2(n_47), .B1(n_255), .B2(n_263), .Y(n_262) );
AOI22xp33_ASAP7_75t_SL g277 ( .A1(n_20), .A2(n_68), .B1(n_278), .B2(n_281), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_21), .A2(n_221), .B1(n_369), .B2(n_445), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_22), .A2(n_106), .B1(n_529), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_23), .A2(n_29), .B1(n_293), .B2(n_294), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_24), .A2(n_196), .B1(n_375), .B2(n_430), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_25), .A2(n_89), .B1(n_376), .B2(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_26), .A2(n_193), .B1(n_285), .B2(n_288), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_28), .A2(n_79), .B1(n_429), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_30), .A2(n_194), .B1(n_269), .B2(n_273), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_31), .A2(n_147), .B1(n_374), .B2(n_584), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_32), .A2(n_62), .B1(n_422), .B2(n_423), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_33), .A2(n_128), .B1(n_510), .B2(n_513), .Y(n_509) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_34), .A2(n_71), .B1(n_103), .B2(n_385), .C1(n_451), .C2(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_35), .A2(n_213), .B1(n_303), .B2(n_319), .Y(n_351) );
XOR2x2_ASAP7_75t_L g568 ( .A(n_36), .B(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_37), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_38), .A2(n_144), .B1(n_423), .B2(n_438), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_39), .A2(n_140), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_40), .A2(n_127), .B1(n_414), .B2(n_567), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_41), .A2(n_211), .B1(n_565), .B2(n_606), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_42), .A2(n_67), .B1(n_473), .B2(n_572), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_43), .A2(n_312), .B1(n_313), .B2(n_327), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_43), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_44), .A2(n_75), .B1(n_297), .B2(n_298), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_45), .A2(n_49), .B1(n_389), .B2(n_482), .Y(n_481) );
AOI222xp33_ASAP7_75t_L g608 ( .A1(n_46), .A2(n_51), .B1(n_210), .B2(n_412), .C1(n_609), .C2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_48), .A2(n_167), .B1(n_269), .B2(n_273), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_52), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_53), .A2(n_85), .B1(n_580), .B2(n_581), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_54), .Y(n_619) );
AOI222xp33_ASAP7_75t_L g652 ( .A1(n_55), .A2(n_123), .B1(n_188), .B2(n_383), .C1(n_385), .C2(n_609), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_56), .A2(n_152), .B1(n_305), .B2(n_306), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_57), .A2(n_116), .B1(n_489), .B2(n_490), .Y(n_488) );
INVx3_ASAP7_75t_L g255 ( .A(n_58), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_59), .A2(n_122), .B1(n_278), .B2(n_325), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_60), .A2(n_109), .B1(n_374), .B2(n_376), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_61), .A2(n_138), .B1(n_443), .B2(n_445), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_63), .A2(n_121), .B1(n_297), .B2(n_298), .Y(n_350) );
OA22x2_ASAP7_75t_L g593 ( .A1(n_64), .A2(n_594), .B1(n_595), .B2(n_611), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_64), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_66), .A2(n_102), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_69), .A2(n_101), .B1(n_285), .B2(n_414), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_70), .B(n_98), .Y(n_239) );
INVx1_ASAP7_75t_SL g256 ( .A(n_70), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_72), .A2(n_182), .B1(n_396), .B2(n_398), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_73), .A2(n_142), .B1(n_372), .B2(n_521), .Y(n_634) );
INVx2_ASAP7_75t_L g229 ( .A(n_74), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_76), .A2(n_130), .B1(n_298), .B2(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_78), .A2(n_223), .B(n_232), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_80), .A2(n_111), .B1(n_458), .B2(n_459), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_81), .A2(n_209), .B1(n_294), .B2(n_347), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_82), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_82), .B(n_441), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_82), .A2(n_462), .B(n_463), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g292 ( .A1(n_83), .A2(n_148), .B1(n_293), .B2(n_294), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_84), .A2(n_178), .B1(n_269), .B2(n_412), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_86), .A2(n_212), .B1(n_363), .B2(n_365), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_87), .A2(n_205), .B1(n_389), .B2(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_88), .A2(n_173), .B1(n_399), .B2(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_91), .A2(n_104), .B1(n_506), .B2(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g501 ( .A(n_92), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g324 ( .A1(n_95), .A2(n_161), .B1(n_278), .B2(n_325), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_96), .A2(n_175), .B1(n_575), .B2(n_576), .Y(n_574) );
AO22x2_ASAP7_75t_L g258 ( .A1(n_98), .A2(n_169), .B1(n_255), .B2(n_259), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_100), .A2(n_184), .B1(n_383), .B2(n_385), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_105), .A2(n_174), .B1(n_516), .B2(n_517), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_107), .A2(n_151), .B1(n_383), .B2(n_385), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_108), .A2(n_157), .B1(n_297), .B2(n_298), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_110), .A2(n_145), .B1(n_396), .B2(n_473), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_112), .Y(n_544) );
AOI22xp33_ASAP7_75t_SL g525 ( .A1(n_113), .A2(n_168), .B1(n_526), .B2(n_529), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_114), .A2(n_125), .B1(n_422), .B2(n_430), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_117), .A2(n_206), .B1(n_556), .B2(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g257 ( .A(n_118), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_119), .A2(n_172), .B1(n_431), .B2(n_535), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_120), .A2(n_219), .B1(n_429), .B2(n_431), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g356 ( .A1(n_124), .A2(n_190), .B1(n_357), .B2(n_360), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_126), .B(n_251), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_133), .A2(n_149), .B1(n_385), .B2(n_451), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_134), .A2(n_136), .B1(n_302), .B2(n_303), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_135), .A2(n_201), .B1(n_294), .B2(n_347), .Y(n_346) );
XNOR2x1_ASAP7_75t_L g353 ( .A(n_137), .B(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_R g537 ( .A(n_139), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_141), .A2(n_187), .B1(n_521), .B2(n_524), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_143), .A2(n_171), .B1(n_479), .B2(n_480), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_146), .B(n_416), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_150), .A2(n_181), .B1(n_503), .B2(n_505), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_153), .A2(n_214), .B1(n_581), .B2(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_154), .A2(n_216), .B1(n_363), .B2(n_365), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_155), .A2(n_199), .B1(n_305), .B2(n_306), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_156), .B(n_379), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_158), .A2(n_170), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_162), .A2(n_179), .B1(n_285), .B2(n_414), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_163), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_164), .A2(n_202), .B1(n_369), .B2(n_372), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_165), .A2(n_220), .B1(n_365), .B2(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_166), .A2(n_192), .B1(n_297), .B2(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_176), .B(n_588), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_177), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g241 ( .A(n_177), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_180), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_183), .A2(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
AND2x2_ASAP7_75t_R g310 ( .A(n_185), .B(n_241), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_186), .A2(n_207), .B1(n_303), .B2(n_319), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_189), .B(n_379), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_191), .A2(n_208), .B1(n_479), .B2(n_586), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_195), .A2(n_200), .B1(n_363), .B2(n_565), .Y(n_564) );
INVxp67_ASAP7_75t_L g231 ( .A(n_197), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_198), .Y(n_561) );
NAND2xp33_ASAP7_75t_SL g628 ( .A(n_204), .B(n_629), .Y(n_628) );
XNOR2xp5_ASAP7_75t_L g246 ( .A(n_215), .B(n_247), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_215), .A2(n_308), .B1(n_311), .B2(n_328), .Y(n_307) );
BUFx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NOR2x1_ASAP7_75t_R g224 ( .A(n_225), .B(n_227), .Y(n_224) );
OR2x2_ASAP7_75t_L g329 ( .A(n_225), .B(n_228), .Y(n_329) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_226), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
OAI211xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_242), .B(n_307), .C(n_330), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
CKINVDCx6p67_ASAP7_75t_R g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
INVx1_ASAP7_75t_L g660 ( .A(n_236), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g659 ( .A(n_240), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_248), .B(n_290), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_276), .Y(n_248) );
OAI21xp5_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_267), .B(n_268), .Y(n_249) );
OAI21xp5_ASAP7_75t_SL g560 ( .A1(n_250), .A2(n_561), .B(n_562), .Y(n_560) );
INVx2_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_L g609 ( .A(n_251), .Y(n_609) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_260), .Y(n_251) );
AND2x2_ASAP7_75t_L g281 ( .A(n_252), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g288 ( .A(n_252), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g325 ( .A(n_252), .B(n_282), .Y(n_325) );
AND2x4_ASAP7_75t_L g359 ( .A(n_252), .B(n_289), .Y(n_359) );
AND2x4_ASAP7_75t_L g366 ( .A(n_252), .B(n_282), .Y(n_366) );
AND2x2_ASAP7_75t_L g381 ( .A(n_252), .B(n_260), .Y(n_381) );
AND2x2_ASAP7_75t_L g414 ( .A(n_252), .B(n_289), .Y(n_414) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_258), .Y(n_252) );
AND2x2_ASAP7_75t_L g271 ( .A(n_253), .B(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
INVx2_ASAP7_75t_L g287 ( .A(n_253), .Y(n_287) );
OAI22x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B1(n_256), .B2(n_257), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g259 ( .A(n_255), .Y(n_259) );
INVx2_ASAP7_75t_L g263 ( .A(n_255), .Y(n_263) );
INVx1_ASAP7_75t_L g266 ( .A(n_255), .Y(n_266) );
INVx2_ASAP7_75t_L g272 ( .A(n_258), .Y(n_272) );
AND2x2_ASAP7_75t_L g286 ( .A(n_258), .B(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_L g295 ( .A(n_258), .Y(n_295) );
AND2x6_ASAP7_75t_L g297 ( .A(n_260), .B(n_286), .Y(n_297) );
AND2x2_ASAP7_75t_L g302 ( .A(n_260), .B(n_271), .Y(n_302) );
AND2x2_ASAP7_75t_L g305 ( .A(n_260), .B(n_299), .Y(n_305) );
AND2x2_ASAP7_75t_L g319 ( .A(n_260), .B(n_271), .Y(n_319) );
AND2x4_ASAP7_75t_L g375 ( .A(n_260), .B(n_271), .Y(n_375) );
AND2x4_ASAP7_75t_L g391 ( .A(n_260), .B(n_299), .Y(n_391) );
AND2x2_ASAP7_75t_L g397 ( .A(n_260), .B(n_286), .Y(n_397) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g270 ( .A(n_262), .B(n_264), .Y(n_270) );
AND2x2_ASAP7_75t_L g275 ( .A(n_262), .B(n_265), .Y(n_275) );
INVx1_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
INVxp67_ASAP7_75t_L g289 ( .A(n_264), .Y(n_289) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g279 ( .A(n_265), .B(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_269), .Y(n_610) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x2_ASAP7_75t_L g285 ( .A(n_270), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g306 ( .A(n_270), .B(n_299), .Y(n_306) );
AND2x4_ASAP7_75t_L g361 ( .A(n_270), .B(n_286), .Y(n_361) );
AND2x2_ASAP7_75t_L g384 ( .A(n_270), .B(n_271), .Y(n_384) );
AND2x4_ASAP7_75t_L g399 ( .A(n_270), .B(n_299), .Y(n_399) );
AND2x2_ASAP7_75t_L g567 ( .A(n_270), .B(n_286), .Y(n_567) );
AND2x4_ASAP7_75t_L g278 ( .A(n_271), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g364 ( .A(n_271), .B(n_279), .Y(n_364) );
AND2x4_ASAP7_75t_L g299 ( .A(n_272), .B(n_287), .Y(n_299) );
AND2x2_ASAP7_75t_SL g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g386 ( .A(n_274), .B(n_275), .Y(n_386) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_274), .B(n_275), .Y(n_412) );
AND2x4_ASAP7_75t_L g294 ( .A(n_275), .B(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g303 ( .A(n_275), .B(n_299), .Y(n_303) );
AND2x4_ASAP7_75t_L g372 ( .A(n_275), .B(n_295), .Y(n_372) );
AND2x4_ASAP7_75t_L g376 ( .A(n_275), .B(n_299), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_284), .Y(n_276) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_279), .B(n_286), .Y(n_293) );
AND2x6_ASAP7_75t_L g298 ( .A(n_279), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g347 ( .A(n_279), .B(n_286), .Y(n_347) );
AND2x2_ASAP7_75t_L g371 ( .A(n_279), .B(n_286), .Y(n_371) );
AND2x4_ASAP7_75t_L g394 ( .A(n_279), .B(n_299), .Y(n_394) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_280), .Y(n_283) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_300), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVx1_ASAP7_75t_L g553 ( .A(n_297), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_313), .Y(n_327) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVxp33_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_322), .Y(n_315) );
NAND4xp25_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .C(n_320), .D(n_321), .Y(n_316) );
NAND3xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .C(n_326), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_329), .Y(n_328) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_591), .B1(n_657), .B2(n_658), .C(n_659), .Y(n_330) );
INVx1_ASAP7_75t_L g658 ( .A(n_331), .Y(n_658) );
XOR2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_465), .Y(n_331) );
XOR2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_402), .Y(n_332) );
AO22x2_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_353), .B1(n_400), .B2(n_401), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
XOR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_352), .Y(n_335) );
XOR2x2_ASAP7_75t_L g401 ( .A(n_336), .B(n_352), .Y(n_401) );
NAND2x1_ASAP7_75t_SL g336 ( .A(n_337), .B(n_344), .Y(n_336) );
NOR2x1_ASAP7_75t_L g337 ( .A(n_338), .B(n_341), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NOR2x1_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx2_ASAP7_75t_L g400 ( .A(n_353), .Y(n_400) );
NAND4xp75_ASAP7_75t_L g354 ( .A(n_355), .B(n_367), .C(n_377), .D(n_387), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_362), .Y(n_355) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g455 ( .A(n_358), .Y(n_455) );
INVx1_ASAP7_75t_L g490 ( .A(n_358), .Y(n_490) );
INVx2_ASAP7_75t_L g517 ( .A(n_358), .Y(n_517) );
INVx2_ASAP7_75t_L g581 ( .A(n_358), .Y(n_581) );
INVx6_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_361), .Y(n_454) );
BUFx3_ASAP7_75t_L g489 ( .A(n_361), .Y(n_489) );
BUFx2_ASAP7_75t_L g580 ( .A(n_361), .Y(n_580) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g487 ( .A(n_364), .Y(n_487) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_364), .Y(n_606) );
BUFx4f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g514 ( .A(n_366), .Y(n_514) );
BUFx6f_ASAP7_75t_SL g565 ( .A(n_366), .Y(n_565) );
BUFx3_ASAP7_75t_L g630 ( .A(n_366), .Y(n_630) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_373), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g523 ( .A(n_370), .Y(n_523) );
INVx1_ASAP7_75t_L g549 ( .A(n_370), .Y(n_549) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g444 ( .A(n_371), .Y(n_444) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_371), .Y(n_479) );
INVx5_ASAP7_75t_SL g446 ( .A(n_372), .Y(n_446) );
BUFx3_ASAP7_75t_L g480 ( .A(n_372), .Y(n_480) );
BUFx2_ASAP7_75t_L g550 ( .A(n_372), .Y(n_550) );
BUFx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx6_ASAP7_75t_L g432 ( .A(n_375), .Y(n_432) );
BUFx3_ASAP7_75t_L g556 ( .A(n_375), .Y(n_556) );
BUFx3_ASAP7_75t_L g430 ( .A(n_376), .Y(n_430) );
INVx2_ASAP7_75t_L g477 ( .A(n_376), .Y(n_477) );
BUFx2_ASAP7_75t_SL g535 ( .A(n_376), .Y(n_535) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_382), .Y(n_377) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_SL g416 ( .A(n_380), .Y(n_416) );
INVx3_ASAP7_75t_L g588 ( .A(n_380), .Y(n_588) );
INVx6_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx3_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx5_ASAP7_75t_L g451 ( .A(n_384), .Y(n_451) );
INVx2_ASAP7_75t_L g504 ( .A(n_384), .Y(n_504) );
BUFx3_ASAP7_75t_L g627 ( .A(n_384), .Y(n_627) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g507 ( .A(n_386), .Y(n_507) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_395), .Y(n_387) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx3_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
INVx3_ASAP7_75t_SL g438 ( .A(n_390), .Y(n_438) );
INVx4_ASAP7_75t_L g528 ( .A(n_390), .Y(n_528) );
INVx2_ASAP7_75t_L g638 ( .A(n_390), .Y(n_638) );
INVx8_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g458 ( .A(n_393), .Y(n_458) );
INVx2_ASAP7_75t_L g473 ( .A(n_393), .Y(n_473) );
INVx2_ASAP7_75t_L g529 ( .A(n_393), .Y(n_529) );
INVx2_ASAP7_75t_L g603 ( .A(n_393), .Y(n_603) );
INVx8_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g460 ( .A(n_396), .Y(n_460) );
BUFx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g573 ( .A(n_397), .Y(n_573) );
BUFx2_ASAP7_75t_L g602 ( .A(n_397), .Y(n_602) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_399), .Y(n_423) );
INVx2_ASAP7_75t_L g483 ( .A(n_399), .Y(n_483) );
BUFx3_ASAP7_75t_L g584 ( .A(n_399), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_425), .B2(n_464), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_417), .Y(n_408) );
NAND4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .C(n_413), .D(n_415), .Y(n_409) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_416), .Y(n_434) );
INVx2_ASAP7_75t_L g500 ( .A(n_416), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_421), .C(n_424), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx2_ASAP7_75t_L g533 ( .A(n_423), .Y(n_533) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_423), .Y(n_636) );
INVx1_ASAP7_75t_L g464 ( .A(n_425), .Y(n_464) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_427), .B(n_447), .Y(n_426) );
A2O1A1Ixp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_433), .B(n_439), .C(n_440), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_428), .B(n_433), .C(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
INVx3_ASAP7_75t_L g575 ( .A(n_432), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_439), .B(n_442), .C(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g524 ( .A(n_446), .Y(n_524) );
INVx3_ASAP7_75t_L g586 ( .A(n_446), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_456), .B(n_461), .Y(n_447) );
INVx1_ASAP7_75t_L g463 ( .A(n_449), .Y(n_463) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_452), .Y(n_449) );
BUFx4f_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g516 ( .A(n_454), .Y(n_516) );
BUFx2_ASAP7_75t_L g624 ( .A(n_454), .Y(n_624) );
INVx1_ASAP7_75t_L g462 ( .A(n_457), .Y(n_462) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_467), .B1(n_540), .B2(n_590), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_493), .B1(n_494), .B2(n_538), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
NOR2xp67_ASAP7_75t_L g470 ( .A(n_471), .B(n_484), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .C(n_478), .D(n_481), .Y(n_471) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_SL g576 ( .A(n_477), .Y(n_576) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g558 ( .A(n_483), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g484 ( .A(n_485), .B(n_488), .C(n_491), .D(n_492), .Y(n_484) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx4_ASAP7_75t_L g512 ( .A(n_487), .Y(n_512) );
INVx1_ASAP7_75t_L g621 ( .A(n_487), .Y(n_621) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AOI22x1_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_536), .B2(n_537), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_518), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_508), .Y(n_498) );
OAI21xp5_ASAP7_75t_SL g499 ( .A1(n_500), .A2(n_501), .B(n_502), .Y(n_499) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NOR2x1_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_525), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .Y(n_530) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g590 ( .A(n_540), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_568), .B2(n_589), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
XNOR2x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_546), .B(n_559), .Y(n_545) );
NOR2x1_ASAP7_75t_L g546 ( .A(n_547), .B(n_554), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx2_ASAP7_75t_L g589 ( .A(n_568), .Y(n_589) );
NAND4xp75_ASAP7_75t_L g569 ( .A(n_570), .B(n_577), .C(n_582), .D(n_587), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g657 ( .A(n_591), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_612), .B1(n_655), .B2(n_656), .Y(n_591) );
INVx1_ASAP7_75t_L g655 ( .A(n_592), .Y(n_655) );
BUFx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g611 ( .A(n_595), .Y(n_611) );
NAND4xp75_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .C(n_604), .D(n_608), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
BUFx3_ASAP7_75t_L g633 ( .A(n_602), .Y(n_633) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g656 ( .A(n_612), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_639), .B1(n_640), .B2(n_654), .Y(n_612) );
INVx2_ASAP7_75t_L g654 ( .A(n_613), .Y(n_654) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
XNOR2x1_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_631), .Y(n_616) );
NAND4xp25_ASAP7_75t_L g617 ( .A(n_618), .B(n_623), .C(n_625), .D(n_628), .Y(n_617) );
OA21x2_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_620), .B(n_622), .Y(n_618) );
INVxp33_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx6f_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
BUFx6f_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .C(n_635), .D(n_637), .Y(n_631) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
XOR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_653), .Y(n_641) );
NAND4xp75_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .C(n_649), .D(n_652), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
endmodule