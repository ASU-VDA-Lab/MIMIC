module fake_jpeg_21766_n_168 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_1),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_3),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_42),
.Y(n_44)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_4),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_48),
.B1(n_38),
.B2(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_18),
.B1(n_17),
.B2(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_55),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_23),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_57),
.C(n_25),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_17),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_35),
.C(n_22),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_5),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_62),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_4),
.Y(n_62)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_38),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_62),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_20),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_71),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_51),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_90),
.Y(n_101)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_5),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_83),
.B(n_91),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_87),
.B(n_8),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_6),
.B1(n_20),
.B2(n_9),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_58),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_50),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_65),
.B1(n_63),
.B2(n_66),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_98),
.B1(n_113),
.B2(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_68),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_66),
.B1(n_53),
.B2(n_49),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_112),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_55),
.B(n_64),
.C(n_6),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_68),
.B1(n_76),
.B2(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_8),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_75),
.B(n_77),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_115),
.C(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_117),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_126),
.B1(n_105),
.B2(n_99),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_89),
.B1(n_81),
.B2(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_84),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_101),
.B(n_95),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_109),
.B(n_96),
.C(n_113),
.D(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_135),
.C(n_115),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_73),
.A3(n_105),
.B1(n_85),
.B2(n_14),
.C1(n_10),
.C2(n_13),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_136),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_137),
.B1(n_118),
.B2(n_124),
.Y(n_141)
);

OA21x2_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_73),
.B(n_72),
.Y(n_136)
);

AND2x4_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_144),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_137),
.B(n_123),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_120),
.C(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_147),
.Y(n_155)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_127),
.C(n_122),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_137),
.B1(n_138),
.B2(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_148),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_152),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_143),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_129),
.B(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_158),
.Y(n_163)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_154),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_129),
.A3(n_119),
.B1(n_117),
.B2(n_107),
.C1(n_14),
.C2(n_12),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_153),
.B1(n_151),
.B2(n_99),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_163),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_166),
.Y(n_168)
);


endmodule