module fake_jpeg_10561_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_3),
.B(n_2),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_10),
.B1(n_8),
.B2(n_12),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_10),
.B1(n_19),
.B2(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_15),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_12),
.C(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_20),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_21),
.B2(n_20),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_7),
.C(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_31),
.C(n_7),
.Y(n_36)
);

A2O1A1O1Ixp25_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_34),
.B(n_17),
.C(n_4),
.D(n_5),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_35),
.B1(n_2),
.B2(n_4),
.Y(n_38)
);

OAI221xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.C(n_17),
.Y(n_39)
);


endmodule