module fake_ariane_785_n_773 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_773);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_773;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_590;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_94),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_28),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_32),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_10),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_107),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_74),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_73),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_14),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_40),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_17),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_0),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_129),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_38),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_20),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_27),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_49),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_13),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_100),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_52),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_51),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_37),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_122),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_41),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_77),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_81),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_21),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_56),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_45),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_75),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_11),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_91),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_30),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_147),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_69),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_13),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_26),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_79),
.Y(n_198)
);

INVxp33_ASAP7_75t_SL g199 ( 
.A(n_140),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_59),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_86),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_60),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_165),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

OAI22x1_ASAP7_75t_R g212 ( 
.A1(n_153),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_154),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

BUFx8_ASAP7_75t_L g222 ( 
.A(n_150),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_173),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_168),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_173),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_158),
.B(n_1),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_178),
.B(n_2),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_196),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_155),
.B(n_3),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_207),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_207),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_R g253 ( 
.A(n_213),
.B(n_148),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_R g263 ( 
.A(n_213),
.B(n_149),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_227),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_176),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_227),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_206),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_233),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_233),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_220),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_190),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_212),
.A2(n_199),
.B1(n_201),
.B2(n_203),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_220),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_211),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_205),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_205),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_210),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_223),
.B(n_202),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_217),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_R g288 ( 
.A(n_245),
.B(n_234),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_217),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_R g291 ( 
.A(n_213),
.B(n_160),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_245),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_234),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_223),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_226),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_226),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_226),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_222),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_222),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_276),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_214),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_256),
.B(n_199),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_222),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_214),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_214),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_247),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_209),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

AOI221xp5_ASAP7_75t_L g315 ( 
.A1(n_274),
.A2(n_238),
.B1(n_248),
.B2(n_219),
.C(n_230),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_256),
.B(n_263),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_256),
.B(n_201),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_236),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_209),
.Y(n_319)
);

BUFx6f_ASAP7_75t_SL g320 ( 
.A(n_251),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_293),
.A2(n_248),
.B1(n_246),
.B2(n_221),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_259),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_257),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_264),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_260),
.B(n_209),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_209),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_266),
.B(n_267),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_209),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_279),
.B(n_231),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_231),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_282),
.B(n_221),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_249),
.B(n_224),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_231),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_250),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_231),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_288),
.B(n_243),
.C(n_241),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_270),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_278),
.B(n_224),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_286),
.B(n_228),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_271),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_281),
.A2(n_228),
.B1(n_246),
.B2(n_232),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_289),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_289),
.B(n_241),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_268),
.B(n_231),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_268),
.B(n_232),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_252),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_258),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_261),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_293),
.A2(n_235),
.B1(n_240),
.B2(n_237),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_288),
.A2(n_193),
.B1(n_172),
.B2(n_174),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_254),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_256),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_294),
.B(n_241),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_294),
.B(n_241),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_249),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_257),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_359),
.B(n_244),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_235),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_241),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_329),
.B(n_157),
.Y(n_367)
);

AO22x1_ASAP7_75t_L g368 ( 
.A1(n_329),
.A2(n_192),
.B1(n_166),
.B2(n_170),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_326),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_243),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_342),
.B(n_243),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_243),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_161),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

AND2x4_ASAP7_75t_SL g376 ( 
.A(n_354),
.B(n_216),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_315),
.A2(n_243),
.B1(n_240),
.B2(n_237),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_318),
.B(n_216),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_305),
.B(n_229),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_313),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_347),
.A2(n_195),
.B1(n_181),
.B2(n_182),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_334),
.Y(n_383)
);

AO22x1_ASAP7_75t_L g384 ( 
.A1(n_346),
.A2(n_197),
.B1(n_188),
.B2(n_189),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_300),
.B(n_179),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_342),
.B(n_194),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_318),
.B(n_216),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_321),
.A2(n_240),
.B1(n_237),
.B2(n_229),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_336),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_303),
.A2(n_198),
.B(n_237),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_353),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_303),
.B(n_216),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_321),
.A2(n_240),
.B1(n_237),
.B2(n_6),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_301),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_342),
.B(n_240),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_360),
.A2(n_83),
.B(n_145),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_320),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_310),
.B(n_4),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_308),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_342),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_302),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_357),
.A2(n_356),
.B1(n_352),
.B2(n_339),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_310),
.B(n_5),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_306),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_300),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_316),
.B(n_7),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_342),
.B(n_298),
.Y(n_416)
);

AND3x1_ASAP7_75t_L g417 ( 
.A(n_311),
.B(n_8),
.C(n_9),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_307),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_361),
.A2(n_88),
.B(n_144),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_322),
.Y(n_420)
);

NAND2x1_ASAP7_75t_SL g421 ( 
.A(n_348),
.B(n_9),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_324),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_349),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_325),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

OR2x2_ASAP7_75t_SL g426 ( 
.A(n_338),
.B(n_10),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_313),
.Y(n_427)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_344),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_429)
);

BUFx6f_ASAP7_75t_SL g430 ( 
.A(n_320),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_327),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_299),
.B(n_12),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_398),
.B(n_369),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_367),
.B(n_350),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_395),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_414),
.B(n_344),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_406),
.B(n_350),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_375),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_383),
.B(n_345),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_390),
.B(n_304),
.Y(n_441)
);

O2A1O1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_413),
.A2(n_317),
.B(n_351),
.C(n_345),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_416),
.A2(n_331),
.B(n_328),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_378),
.B(n_312),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_414),
.B(n_319),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_385),
.A2(n_337),
.B(n_333),
.C(n_332),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_374),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_363),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_407),
.B(n_363),
.Y(n_449)
);

NAND2x1_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_363),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_430),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_400),
.Y(n_452)
);

NOR2x1_ASAP7_75t_L g453 ( 
.A(n_392),
.B(n_15),
.Y(n_453)
);

OR2x6_ASAP7_75t_SL g454 ( 
.A(n_432),
.B(n_430),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_415),
.A2(n_90),
.B(n_142),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_415),
.A2(n_89),
.B(n_141),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_421),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_386),
.B(n_15),
.Y(n_458)
);

OR2x6_ASAP7_75t_SL g459 ( 
.A(n_368),
.B(n_16),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_401),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_426),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_393),
.A2(n_93),
.B(n_139),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_410),
.B(n_18),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_372),
.B(n_19),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_19),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_403),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_373),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_379),
.B(n_388),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_429),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_471)
);

A2O1A1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_25),
.B(n_29),
.C(n_31),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_366),
.B(n_33),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_387),
.A2(n_34),
.B(n_35),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_371),
.A2(n_431),
.B(n_370),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_402),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_381),
.B(n_428),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_377),
.B(n_43),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_405),
.B(n_44),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_377),
.B(n_46),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_396),
.A2(n_47),
.B(n_48),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_394),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_404),
.B(n_55),
.Y(n_485)
);

O2A1O1Ixp33_ASAP7_75t_L g486 ( 
.A1(n_411),
.A2(n_364),
.B(n_409),
.C(n_391),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_408),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_443),
.A2(n_397),
.B(n_419),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_470),
.A2(n_380),
.B(n_427),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_474),
.A2(n_365),
.B(n_380),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_447),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_434),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_434),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_476),
.A2(n_475),
.B(n_462),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_448),
.Y(n_498)
);

AND2x4_ASAP7_75t_SL g499 ( 
.A(n_465),
.B(n_394),
.Y(n_499)
);

AO21x2_ASAP7_75t_L g500 ( 
.A1(n_480),
.A2(n_365),
.B(n_424),
.Y(n_500)
);

CKINVDCx6p67_ASAP7_75t_R g501 ( 
.A(n_451),
.Y(n_501)
);

AO21x2_ASAP7_75t_L g502 ( 
.A1(n_482),
.A2(n_422),
.B(n_420),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_465),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_435),
.B(n_417),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_473),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_433),
.Y(n_506)
);

AO21x2_ASAP7_75t_L g507 ( 
.A1(n_467),
.A2(n_412),
.B(n_418),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_469),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_452),
.Y(n_509)
);

AO21x2_ASAP7_75t_L g510 ( 
.A1(n_463),
.A2(n_389),
.B(n_376),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_455),
.A2(n_428),
.B(n_384),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_457),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_456),
.A2(n_428),
.B(n_382),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_473),
.Y(n_515)
);

BUFx2_ASAP7_75t_SL g516 ( 
.A(n_473),
.Y(n_516)
);

AOI22x1_ASAP7_75t_L g517 ( 
.A1(n_464),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_440),
.B(n_62),
.Y(n_518)
);

AOI22x1_ASAP7_75t_L g519 ( 
.A1(n_483),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_439),
.B(n_66),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_485),
.A2(n_68),
.B(n_70),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_436),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g523 ( 
.A1(n_446),
.A2(n_71),
.B(n_72),
.Y(n_523)
);

BUFx8_ASAP7_75t_L g524 ( 
.A(n_479),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_486),
.A2(n_76),
.B(n_78),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_477),
.A2(n_80),
.B(n_82),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_468),
.Y(n_527)
);

AO21x1_ASAP7_75t_L g528 ( 
.A1(n_442),
.A2(n_84),
.B(n_85),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_438),
.B(n_92),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_439),
.B(n_95),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_479),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_504),
.A2(n_437),
.B1(n_461),
.B2(n_484),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_492),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_511),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_511),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_527),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_522),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_507),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_494),
.B(n_479),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_504),
.A2(n_459),
.B1(n_441),
.B2(n_458),
.Y(n_543)
);

AOI21x1_ASAP7_75t_L g544 ( 
.A1(n_528),
.A2(n_449),
.B(n_450),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_501),
.Y(n_545)
);

INVx6_ASAP7_75t_L g546 ( 
.A(n_524),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_516),
.B(n_444),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_531),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_497),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_522),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_531),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_498),
.B(n_445),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_497),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_506),
.B(n_444),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_499),
.A2(n_481),
.B1(n_453),
.B2(n_454),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_510),
.A2(n_472),
.B1(n_471),
.B2(n_478),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_496),
.A2(n_96),
.B(n_97),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_507),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_510),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_493),
.B(n_102),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_497),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_496),
.A2(n_103),
.B(n_104),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_513),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_497),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_494),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_502),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_520),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_493),
.B(n_146),
.Y(n_569)
);

CKINVDCx11_ASAP7_75t_R g570 ( 
.A(n_501),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_524),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_SL g572 ( 
.A1(n_499),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_508),
.A2(n_110),
.B1(n_111),
.B2(n_113),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_548),
.Y(n_574)
);

AO31x2_ASAP7_75t_L g575 ( 
.A1(n_567),
.A2(n_528),
.A3(n_490),
.B(n_529),
.Y(n_575)
);

OAI222xp33_ASAP7_75t_L g576 ( 
.A1(n_534),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.C1(n_520),
.C2(n_530),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_533),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_534),
.A2(n_525),
.B(n_526),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_543),
.A2(n_517),
.B1(n_510),
.B2(n_523),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_568),
.A2(n_530),
.B1(n_520),
.B2(n_509),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_552),
.B(n_495),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_535),
.B(n_495),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_546),
.B(n_516),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_542),
.B(n_532),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_545),
.B(n_509),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_564),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_536),
.B(n_515),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

AOI221xp5_ASAP7_75t_L g589 ( 
.A1(n_552),
.A2(n_523),
.B1(n_530),
.B2(n_520),
.C(n_532),
.Y(n_589)
);

BUFx6f_ASAP7_75t_SL g590 ( 
.A(n_571),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_R g591 ( 
.A(n_545),
.B(n_524),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_542),
.B(n_532),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_569),
.B(n_515),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_538),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_539),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_546),
.B(n_505),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_547),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_551),
.B(n_497),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_554),
.B(n_546),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_566),
.B(n_505),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_549),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_570),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_540),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_SL g605 ( 
.A(n_570),
.B(n_505),
.C(n_503),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_560),
.B(n_503),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_549),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_503),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_550),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_547),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_547),
.B(n_488),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_555),
.B(n_488),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_549),
.Y(n_613)
);

INVx8_ASAP7_75t_L g614 ( 
.A(n_549),
.Y(n_614)
);

AO31x2_ASAP7_75t_L g615 ( 
.A1(n_567),
.A2(n_500),
.A3(n_502),
.B(n_491),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_550),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_541),
.B(n_488),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_541),
.B(n_502),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_553),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_558),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_SL g621 ( 
.A(n_573),
.B(n_544),
.C(n_563),
.Y(n_621)
);

AND2x4_ASAP7_75t_SL g622 ( 
.A(n_583),
.B(n_553),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_578),
.A2(n_556),
.B1(n_572),
.B2(n_559),
.Y(n_623)
);

OAI211xp5_ASAP7_75t_L g624 ( 
.A1(n_578),
.A2(n_556),
.B(n_559),
.C(n_519),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_620),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_580),
.B(n_562),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_580),
.A2(n_530),
.B1(n_561),
.B2(n_565),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_581),
.B(n_565),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_619),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_600),
.B(n_561),
.Y(n_630)
);

NAND2x1_ASAP7_75t_L g631 ( 
.A(n_583),
.B(n_553),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_589),
.B(n_553),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_588),
.B(n_514),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_523),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_614),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_594),
.B(n_514),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_595),
.B(n_557),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_574),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_599),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_609),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_593),
.B(n_500),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_616),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_617),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_617),
.B(n_512),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_604),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_615),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_598),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_608),
.B(n_521),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_615),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_610),
.A2(n_526),
.B1(n_521),
.B2(n_512),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_611),
.B(n_606),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_598),
.Y(n_653)
);

NOR2x1_ASAP7_75t_SL g654 ( 
.A(n_583),
.B(n_491),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_582),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_644),
.B(n_607),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_632),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_639),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_640),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_643),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_648),
.B(n_587),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_655),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_641),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_652),
.B(n_613),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_648),
.Y(n_665)
);

NAND4xp25_ASAP7_75t_L g666 ( 
.A(n_629),
.B(n_624),
.C(n_623),
.D(n_635),
.Y(n_666)
);

NAND4xp25_ASAP7_75t_SL g667 ( 
.A(n_628),
.B(n_579),
.C(n_612),
.D(n_591),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_641),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_653),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_629),
.B(n_576),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_630),
.B(n_602),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_642),
.B(n_618),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_638),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_646),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_633),
.B(n_602),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_645),
.B(n_575),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_633),
.B(n_601),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_645),
.B(n_575),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_634),
.B(n_637),
.C(n_621),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_645),
.B(n_575),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_649),
.B(n_615),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_676),
.B(n_626),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_668),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_673),
.B(n_634),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_656),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_665),
.B(n_634),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_659),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_673),
.B(n_637),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_660),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_668),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_657),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_669),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_676),
.B(n_626),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_679),
.B(n_637),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_672),
.B(n_626),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_678),
.B(n_638),
.Y(n_696)
);

INVxp33_ASAP7_75t_L g697 ( 
.A(n_695),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_687),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_687),
.B(n_656),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_685),
.B(n_686),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_685),
.B(n_661),
.Y(n_701)
);

NAND4xp25_ASAP7_75t_L g702 ( 
.A(n_691),
.B(n_666),
.C(n_670),
.D(n_677),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_689),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_689),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_692),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_694),
.A2(n_667),
.B1(n_670),
.B2(n_681),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_700),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_698),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_706),
.A2(n_694),
.B1(n_684),
.B2(n_688),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_SL g710 ( 
.A1(n_702),
.A2(n_694),
.B(n_696),
.Y(n_710)
);

OAI221xp5_ASAP7_75t_L g711 ( 
.A1(n_710),
.A2(n_702),
.B1(n_662),
.B2(n_705),
.C(n_699),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_708),
.Y(n_712)
);

AOI21xp33_ASAP7_75t_L g713 ( 
.A1(n_709),
.A2(n_675),
.B(n_697),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_707),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_707),
.B(n_696),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_SL g716 ( 
.A1(n_711),
.A2(n_704),
.B(n_703),
.Y(n_716)
);

NOR3x1_ASAP7_75t_L g717 ( 
.A(n_714),
.B(n_701),
.C(n_603),
.Y(n_717)
);

AOI221xp5_ASAP7_75t_L g718 ( 
.A1(n_713),
.A2(n_678),
.B1(n_680),
.B2(n_658),
.C(n_651),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_715),
.B(n_590),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_718),
.A2(n_716),
.B1(n_719),
.B2(n_712),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_717),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_716),
.A2(n_715),
.B(n_680),
.Y(n_722)
);

OAI211xp5_ASAP7_75t_L g723 ( 
.A1(n_720),
.A2(n_585),
.B(n_605),
.C(n_636),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_722),
.B(n_664),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_721),
.B(n_596),
.C(n_671),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_723),
.B(n_636),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_725),
.B(n_724),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_723),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_723),
.A2(n_590),
.B1(n_693),
.B2(n_682),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_724),
.A2(n_681),
.B1(n_693),
.B2(n_682),
.Y(n_730)
);

CKINVDCx16_ASAP7_75t_R g731 ( 
.A(n_724),
.Y(n_731)
);

INVx3_ASAP7_75t_SL g732 ( 
.A(n_731),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_727),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_728),
.B(n_664),
.Y(n_734)
);

NAND4xp25_ASAP7_75t_L g735 ( 
.A(n_726),
.B(n_627),
.C(n_688),
.D(n_684),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_729),
.B(n_688),
.Y(n_736)
);

INVxp33_ASAP7_75t_SL g737 ( 
.A(n_730),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_731),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_738),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_732),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_733),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_734),
.Y(n_742)
);

AND3x1_ASAP7_75t_L g743 ( 
.A(n_736),
.B(n_690),
.C(n_683),
.Y(n_743)
);

XNOR2x1_ASAP7_75t_L g744 ( 
.A(n_737),
.B(n_695),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_735),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_732),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_746),
.B(n_684),
.Y(n_747)
);

XNOR2xp5_ASAP7_75t_L g748 ( 
.A(n_740),
.B(n_597),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_741),
.A2(n_638),
.B1(n_631),
.B2(n_672),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_740),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_742),
.Y(n_751)
);

XOR2xp5_ASAP7_75t_L g752 ( 
.A(n_744),
.B(n_592),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_739),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_745),
.Y(n_754)
);

XNOR2x1_ASAP7_75t_L g755 ( 
.A(n_743),
.B(n_592),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_750),
.B(n_751),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_755),
.A2(n_651),
.B1(n_663),
.B2(n_674),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_752),
.A2(n_690),
.B1(n_683),
.B2(n_584),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_753),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_754),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_748),
.A2(n_747),
.B1(n_749),
.B2(n_584),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_R g762 ( 
.A1(n_759),
.A2(n_646),
.B1(n_650),
.B2(n_647),
.Y(n_762)
);

OAI22x1_ASAP7_75t_L g763 ( 
.A1(n_760),
.A2(n_614),
.B1(n_622),
.B2(n_647),
.Y(n_763)
);

OAI22x1_ASAP7_75t_L g764 ( 
.A1(n_756),
.A2(n_614),
.B1(n_622),
.B2(n_650),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_757),
.A2(n_489),
.B1(n_625),
.B2(n_654),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_761),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_758),
.B(n_489),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_SL g768 ( 
.A1(n_765),
.A2(n_625),
.B1(n_117),
.B2(n_118),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_763),
.Y(n_769)
);

AOI21xp33_ASAP7_75t_SL g770 ( 
.A1(n_769),
.A2(n_764),
.B(n_762),
.Y(n_770)
);

AOI222xp33_ASAP7_75t_L g771 ( 
.A1(n_770),
.A2(n_767),
.B1(n_768),
.B2(n_121),
.C1(n_123),
.C2(n_125),
.Y(n_771)
);

AOI221xp5_ASAP7_75t_L g772 ( 
.A1(n_771),
.A2(n_116),
.B1(n_120),
.B2(n_126),
.C(n_128),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_SL g773 ( 
.A1(n_772),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_773)
);


endmodule