module fake_netlist_6_167_n_1859 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1859);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1859;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_55),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_84),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_41),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_118),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_16),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_40),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_20),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_48),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_93),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_48),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_54),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_86),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_13),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_91),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_67),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_110),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_63),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_8),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_163),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_127),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_51),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_89),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_87),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_11),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_14),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_45),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_62),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_29),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_67),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_137),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_120),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_143),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_71),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_32),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_18),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_119),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_134),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_53),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_111),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_136),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_70),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_22),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_47),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_152),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_65),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_112),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_32),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_28),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_129),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_79),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_151),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_109),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_166),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_55),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_82),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_5),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_49),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_102),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_75),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_39),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_18),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_47),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_45),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_22),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_2),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_0),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_103),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_40),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_144),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_116),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_36),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_26),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_58),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_56),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_88),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_157),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_28),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_26),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_160),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_168),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_52),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_46),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_41),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_68),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_162),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_132),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_9),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_2),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_72),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_114),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_3),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_138),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_81),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_52),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_153),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_133),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_58),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_23),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_94),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_123),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_12),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_113),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_11),
.Y(n_292)
);

BUFx5_ASAP7_75t_L g293 ( 
.A(n_141),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_53),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_25),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_36),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_16),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_98),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_37),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_21),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_35),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_128),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_35),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_90),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_147),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_46),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_92),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_165),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_164),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_59),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_3),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_66),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_4),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_64),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_77),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_4),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_10),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_69),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_14),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_85),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_5),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_19),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_125),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_121),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_8),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_19),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_39),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g329 ( 
.A(n_159),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_95),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_13),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_161),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_155),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_1),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_1),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_7),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_179),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_251),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_174),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_219),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_188),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_177),
.B(n_0),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_223),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_251),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_251),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_230),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_251),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_239),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_7),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_231),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_177),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_261),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_191),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_194),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_244),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_196),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_199),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_201),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_200),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_205),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_261),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_175),
.B(n_9),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_175),
.B(n_12),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_261),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_261),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_214),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_261),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_216),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_182),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_217),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_182),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_249),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_293),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_249),
.B(n_15),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g378 ( 
.A(n_181),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_263),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_171),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_181),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_190),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_180),
.B(n_15),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_190),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_173),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_220),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_221),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_197),
.B(n_17),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_224),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_301),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_226),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_198),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_198),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_235),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_211),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_211),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_236),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_242),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_178),
.B(n_185),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_252),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_242),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_238),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_256),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_178),
.B(n_17),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_262),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_200),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_243),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_170),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_243),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_185),
.B(n_20),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_186),
.B(n_21),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_231),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_246),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_266),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_246),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_271),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_247),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_247),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_352),
.B(n_329),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_343),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_276),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_365),
.A2(n_240),
.B1(n_218),
.B2(n_209),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_245),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_362),
.B(n_277),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_339),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_343),
.A2(n_376),
.B(n_349),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_349),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_284),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_366),
.B(n_288),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_404),
.A2(n_264),
.B1(n_286),
.B2(n_195),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_316),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_400),
.B(n_329),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_346),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_347),
.B(n_213),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_347),
.A2(n_355),
.B(n_350),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_349),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_376),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_350),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_411),
.B(n_186),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_400),
.B(n_329),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_383),
.B(n_329),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_367),
.B(n_289),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_354),
.B(n_353),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_340),
.B(n_342),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_370),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_383),
.B(n_332),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_370),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_354),
.B(n_298),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_372),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_374),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_374),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_375),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_375),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_381),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_382),
.B(n_183),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_392),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_392),
.B(n_303),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

INVxp33_ASAP7_75t_SL g475 ( 
.A(n_390),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_395),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_395),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_377),
.B(n_213),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_398),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_401),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_407),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_337),
.A2(n_336),
.B1(n_335),
.B2(n_331),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_356),
.B(n_193),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_409),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_413),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_413),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_415),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_353),
.B(n_283),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_357),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_422),
.B(n_359),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_454),
.B(n_447),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_344),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_441),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_454),
.B(n_412),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_422),
.B(n_360),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_447),
.A2(n_377),
.B1(n_344),
.B2(n_283),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_440),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_493),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_440),
.B(n_293),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_493),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_440),
.Y(n_508)
);

BUFx4f_ASAP7_75t_L g509 ( 
.A(n_440),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_461),
.B(n_412),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_439),
.B(n_193),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_421),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_388),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_431),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_427),
.B(n_361),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_419),
.B(n_363),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_427),
.B(n_369),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_L g521 ( 
.A(n_419),
.B(n_371),
.Y(n_521)
);

OAI22xp33_ASAP7_75t_L g522 ( 
.A1(n_435),
.A2(n_436),
.B1(n_434),
.B2(n_423),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_441),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_434),
.B(n_373),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_431),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

OAI22xp33_ASAP7_75t_L g527 ( 
.A1(n_435),
.A2(n_378),
.B1(n_388),
.B2(n_297),
.Y(n_527)
);

INVxp33_ASAP7_75t_SL g528 ( 
.A(n_457),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_431),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_436),
.B(n_387),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_425),
.B(n_389),
.Y(n_531)
);

BUFx8_ASAP7_75t_SL g532 ( 
.A(n_441),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_433),
.B(n_391),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_440),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_442),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_461),
.B(n_487),
.C(n_473),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_442),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g539 ( 
.A(n_457),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_487),
.B(n_183),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_429),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_454),
.A2(n_327),
.B1(n_265),
.B2(n_299),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_203),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_431),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_482),
.B(n_415),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_494),
.B(n_397),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_482),
.A2(n_327),
.B1(n_250),
.B2(n_255),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_494),
.B(n_402),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_431),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_494),
.B(n_215),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_442),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g552 ( 
.A1(n_429),
.A2(n_225),
.B(n_215),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_482),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_442),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_475),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_431),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_462),
.B(n_417),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_433),
.B(n_403),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_475),
.B(n_405),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_431),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_479),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_453),
.B(n_416),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_448),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_424),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_473),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_437),
.B(n_386),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_483),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_483),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_439),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_420),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_462),
.B(n_227),
.C(n_225),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_451),
.A2(n_299),
.B1(n_265),
.B2(n_250),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_420),
.B(n_293),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_439),
.B(n_227),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_426),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_453),
.B(n_305),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_448),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_439),
.B(n_306),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_426),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_451),
.A2(n_255),
.B1(n_315),
.B2(n_336),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_443),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_439),
.A2(n_315),
.B1(n_317),
.B2(n_331),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_448),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_428),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_479),
.B(n_308),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_420),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_479),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_469),
.B(n_417),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_443),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_443),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_469),
.B(n_418),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_444),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_420),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_423),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_444),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_437),
.B(n_394),
.Y(n_600)
);

INVx4_ASAP7_75t_SL g601 ( 
.A(n_471),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_444),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_479),
.Y(n_603)
);

INVxp33_ASAP7_75t_L g604 ( 
.A(n_485),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_444),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_479),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_420),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_472),
.B(n_478),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_449),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_450),
.B(n_414),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_449),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_450),
.B(n_384),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_448),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_449),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_428),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_459),
.B(n_380),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_472),
.B(n_293),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_430),
.Y(n_618)
);

AND2x2_ASAP7_75t_SL g619 ( 
.A(n_483),
.B(n_237),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_430),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_459),
.B(n_203),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_432),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_432),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_448),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_438),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_449),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_438),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_472),
.A2(n_317),
.B1(n_335),
.B2(n_237),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_452),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_445),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_485),
.B(n_232),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_483),
.B(n_385),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_470),
.A2(n_270),
.B1(n_233),
.B2(n_229),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_452),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_470),
.B(n_418),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_474),
.B(n_396),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_471),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_452),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_483),
.B(n_332),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_R g640 ( 
.A(n_472),
.B(n_172),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_472),
.B(n_293),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_452),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_478),
.A2(n_232),
.B1(n_321),
.B2(n_309),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_483),
.B(n_332),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_483),
.B(n_310),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_445),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_558),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_541),
.B(n_241),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_530),
.B(n_345),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_531),
.B(n_348),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_540),
.B(n_478),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_540),
.B(n_537),
.Y(n_652)
);

INVx8_ASAP7_75t_L g653 ( 
.A(n_513),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_541),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_558),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_540),
.B(n_203),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_559),
.B(n_478),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_537),
.B(n_203),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_568),
.B(n_478),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_499),
.B(n_351),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_496),
.B(n_483),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_496),
.B(n_203),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_508),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_522),
.A2(n_471),
.B1(n_484),
.B2(n_486),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_508),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_528),
.B(n_358),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_508),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_572),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_504),
.B(n_293),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_509),
.B(n_204),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_495),
.B(n_484),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_515),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_509),
.B(n_204),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_500),
.B(n_516),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_515),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g676 ( 
.A(n_504),
.B(n_293),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_515),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_520),
.B(n_484),
.Y(n_678)
);

INVxp33_ASAP7_75t_L g679 ( 
.A(n_499),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_566),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_566),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_509),
.B(n_606),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_533),
.B(n_484),
.Y(n_683)
);

OAI221xp5_ASAP7_75t_L g684 ( 
.A1(n_501),
.A2(n_384),
.B1(n_396),
.B2(n_489),
.C(n_488),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_524),
.B(n_379),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_563),
.B(n_176),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_592),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_606),
.A2(n_480),
.B(n_476),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_503),
.A2(n_319),
.B1(n_324),
.B2(n_325),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_603),
.B(n_484),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_612),
.B(n_184),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_523),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_592),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_612),
.B(n_187),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_580),
.B(n_484),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_509),
.B(n_204),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g697 ( 
.A(n_569),
.B(n_192),
.C(n_189),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_572),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_498),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_615),
.B(n_484),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_615),
.B(n_484),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_567),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_615),
.B(n_486),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_503),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_560),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_622),
.B(n_486),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_595),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_619),
.B(n_504),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_579),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_619),
.A2(n_471),
.B1(n_486),
.B2(n_253),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_595),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_622),
.B(n_486),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_622),
.B(n_486),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_625),
.B(n_486),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_625),
.B(n_486),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_635),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_572),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_625),
.B(n_446),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_553),
.B(n_446),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_635),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_619),
.B(n_204),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_553),
.B(n_456),
.Y(n_722)
);

INVx8_ASAP7_75t_L g723 ( 
.A(n_513),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_600),
.B(n_259),
.C(n_254),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_498),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_554),
.B(n_456),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_554),
.B(n_458),
.Y(n_727)
);

AND2x6_ASAP7_75t_SL g728 ( 
.A(n_631),
.B(n_241),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_579),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_583),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_504),
.B(n_204),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_507),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_610),
.B(n_260),
.C(n_248),
.Y(n_733)
);

BUFx6f_ASAP7_75t_SL g734 ( 
.A(n_631),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_504),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_583),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_510),
.B(n_202),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_507),
.B(n_253),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_535),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_504),
.B(n_330),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_588),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_588),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_510),
.B(n_268),
.C(n_228),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_562),
.B(n_333),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_562),
.B(n_458),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_573),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_591),
.B(n_464),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_591),
.B(n_464),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_618),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_618),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_502),
.B(n_463),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_502),
.B(n_464),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_535),
.B(n_206),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_534),
.B(n_464),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_534),
.B(n_257),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_620),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_620),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_497),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_511),
.A2(n_471),
.B1(n_321),
.B2(n_309),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_623),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_636),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_511),
.B(n_463),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_556),
.B(n_474),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_623),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_545),
.B(n_464),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_616),
.B(n_207),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_546),
.B(n_210),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_636),
.B(n_477),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_627),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_556),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_545),
.B(n_468),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_511),
.B(n_468),
.Y(n_772)
);

INVx8_ASAP7_75t_L g773 ( 
.A(n_513),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_511),
.B(n_468),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_578),
.B(n_468),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_578),
.B(n_468),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_627),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_630),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_630),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_578),
.B(n_646),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_539),
.B(n_477),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_578),
.B(n_463),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_646),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_573),
.B(n_476),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_550),
.B(n_481),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_608),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_573),
.B(n_476),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_573),
.B(n_463),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_L g789 ( 
.A(n_548),
.B(n_481),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_590),
.B(n_597),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_590),
.B(n_463),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_608),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_590),
.Y(n_793)
);

AO221x1_ASAP7_75t_L g794 ( 
.A1(n_527),
.A2(n_272),
.B1(n_273),
.B2(n_291),
.C(n_285),
.Y(n_794)
);

NAND3xp33_ASAP7_75t_L g795 ( 
.A(n_542),
.B(n_294),
.C(n_222),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_633),
.B(n_295),
.C(n_234),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_497),
.A2(n_257),
.B1(n_291),
.B2(n_285),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_590),
.B(n_476),
.Y(n_798)
);

AND2x6_ASAP7_75t_SL g799 ( 
.A(n_631),
.B(n_267),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_505),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_597),
.B(n_480),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_597),
.B(n_463),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_632),
.B(n_212),
.C(n_258),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_497),
.A2(n_267),
.B1(n_281),
.B2(n_280),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_497),
.B(n_488),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_505),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_505),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_497),
.B(n_517),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_597),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_604),
.A2(n_282),
.B(n_281),
.C(n_280),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_589),
.B(n_480),
.Y(n_811)
);

NOR2xp67_ASAP7_75t_L g812 ( 
.A(n_574),
.B(n_489),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_521),
.B(n_269),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_582),
.B(n_480),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_512),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_514),
.B(n_491),
.Y(n_816)
);

OR2x6_ASAP7_75t_L g817 ( 
.A(n_513),
.B(n_272),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_674),
.B(n_550),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_735),
.B(n_514),
.Y(n_819)
);

OAI22x1_ASAP7_75t_L g820 ( 
.A1(n_699),
.A2(n_598),
.B1(n_633),
.B2(n_631),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_659),
.B(n_550),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_761),
.B(n_631),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_735),
.B(n_506),
.Y(n_823)
);

NOR2x1_ASAP7_75t_L g824 ( 
.A(n_763),
.B(n_513),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_766),
.A2(n_506),
.B(n_575),
.C(n_584),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_725),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_680),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_678),
.A2(n_683),
.B(n_708),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_708),
.A2(n_624),
.B(n_549),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_652),
.A2(n_550),
.B1(n_640),
.B2(n_645),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_663),
.B(n_514),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_681),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_681),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_660),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_770),
.B(n_574),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_695),
.A2(n_624),
.B(n_549),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_652),
.A2(n_550),
.B1(n_639),
.B2(n_644),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_679),
.B(n_514),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_761),
.B(n_601),
.Y(n_839)
);

AO21x1_ASAP7_75t_L g840 ( 
.A1(n_656),
.A2(n_641),
.B(n_617),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_671),
.A2(n_624),
.B(n_549),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_811),
.A2(n_557),
.B(n_544),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_670),
.A2(n_529),
.B(n_525),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_679),
.B(n_525),
.Y(n_844)
);

NOR2x1_ASAP7_75t_R g845 ( 
.A(n_781),
.B(n_274),
.Y(n_845)
);

NOR3xp33_ASAP7_75t_L g846 ( 
.A(n_649),
.B(n_621),
.C(n_490),
.Y(n_846)
);

AOI21x1_ASAP7_75t_L g847 ( 
.A1(n_670),
.A2(n_696),
.B(n_673),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_702),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_663),
.B(n_525),
.Y(n_849)
);

AND2x2_ASAP7_75t_SL g850 ( 
.A(n_808),
.B(n_273),
.Y(n_850)
);

INVx5_ASAP7_75t_L g851 ( 
.A(n_653),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_786),
.B(n_552),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_704),
.B(n_601),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_814),
.A2(n_557),
.B(n_544),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_792),
.B(n_552),
.Y(n_855)
);

AOI21x1_ASAP7_75t_L g856 ( 
.A1(n_673),
.A2(n_641),
.B(n_518),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_682),
.A2(n_544),
.B(n_557),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_686),
.B(n_552),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_696),
.A2(n_751),
.B(n_731),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_753),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_704),
.B(n_552),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_682),
.A2(n_557),
.B(n_544),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_668),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_732),
.B(n_525),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_702),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_768),
.B(n_586),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_661),
.A2(n_587),
.B(n_564),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_657),
.A2(n_780),
.B(n_731),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_729),
.B(n_529),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_690),
.A2(n_587),
.B(n_564),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_665),
.B(n_529),
.Y(n_871)
);

AOI21xp33_ASAP7_75t_L g872 ( 
.A1(n_813),
.A2(n_547),
.B(n_282),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_651),
.A2(n_577),
.B(n_538),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_691),
.A2(n_576),
.B(n_643),
.C(n_628),
.Y(n_874)
);

INVx1_ASAP7_75t_SL g875 ( 
.A(n_692),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_665),
.B(n_570),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_765),
.A2(n_564),
.B(n_565),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_692),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_741),
.B(n_512),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_737),
.B(n_208),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_751),
.A2(n_577),
.B(n_512),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_771),
.A2(n_565),
.B(n_564),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_747),
.A2(n_565),
.B(n_581),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_656),
.A2(n_576),
.B(n_490),
.C(n_518),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_667),
.A2(n_607),
.B1(n_613),
.B2(n_570),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_756),
.B(n_518),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_805),
.A2(n_543),
.B1(n_607),
.B2(n_613),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_694),
.A2(n_607),
.B(n_613),
.C(n_536),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_667),
.A2(n_613),
.B1(n_570),
.B2(n_571),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_668),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_739),
.B(n_650),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_685),
.B(n_705),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_672),
.B(n_570),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_777),
.B(n_526),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_748),
.A2(n_581),
.B(n_587),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_709),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_752),
.A2(n_581),
.B(n_587),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_754),
.A2(n_581),
.B(n_565),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_672),
.B(n_570),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_675),
.B(n_570),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_778),
.B(n_526),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_790),
.A2(n_561),
.B(n_519),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_705),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_772),
.A2(n_775),
.B(n_774),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_662),
.A2(n_577),
.B(n_526),
.C(n_536),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_705),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_709),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_779),
.B(n_536),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_743),
.B(n_675),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_767),
.B(n_73),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_658),
.A2(n_593),
.B(n_538),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_783),
.B(n_538),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_730),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_653),
.B(n_543),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_677),
.B(n_571),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_658),
.A2(n_593),
.B(n_551),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_776),
.A2(n_519),
.B(n_561),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_666),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_785),
.A2(n_543),
.B1(n_571),
.B2(n_585),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_677),
.A2(n_571),
.B1(n_551),
.B2(n_599),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_736),
.B(n_551),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_762),
.A2(n_519),
.B(n_561),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_742),
.B(n_749),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_762),
.A2(n_519),
.B(n_561),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_668),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_647),
.B(n_208),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_655),
.B(n_275),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_668),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_782),
.A2(n_519),
.B(n_561),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_687),
.B(n_278),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_742),
.B(n_555),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_662),
.A2(n_594),
.B(n_555),
.C(n_585),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_782),
.A2(n_519),
.B(n_561),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_SL g934 ( 
.A(n_734),
.B(n_532),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_669),
.A2(n_596),
.B(n_555),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_700),
.A2(n_571),
.B(n_594),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_749),
.B(n_585),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_693),
.B(n_208),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_701),
.A2(n_571),
.B(n_596),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_750),
.B(n_593),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_707),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_703),
.A2(n_599),
.B(n_594),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_706),
.A2(n_596),
.B(n_599),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_717),
.B(n_602),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_711),
.B(n_252),
.Y(n_945)
);

NAND2xp33_ASAP7_75t_SL g946 ( 
.A(n_734),
.B(n_279),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_750),
.B(n_602),
.Y(n_947)
);

NOR2xp67_ASAP7_75t_L g948 ( 
.A(n_796),
.B(n_74),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_712),
.A2(n_602),
.B(n_605),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_795),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_757),
.B(n_605),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_716),
.B(n_601),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_757),
.B(n_605),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_760),
.B(n_609),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_717),
.B(n_601),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_760),
.B(n_609),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_717),
.B(n_601),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_810),
.A2(n_720),
.B(n_764),
.C(n_769),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_764),
.B(n_609),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_SL g960 ( 
.A1(n_721),
.A2(n_642),
.B(n_638),
.C(n_634),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_789),
.A2(n_642),
.B(n_638),
.C(n_611),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_810),
.A2(n_642),
.B(n_638),
.C(n_634),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_713),
.A2(n_637),
.B(n_634),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_769),
.B(n_611),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_745),
.B(n_611),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_755),
.A2(n_721),
.B(n_684),
.C(n_797),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_738),
.B(n_287),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_738),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_669),
.A2(n_676),
.B(n_740),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_793),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_809),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_717),
.B(n_637),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_698),
.A2(n_614),
.B1(n_629),
.B2(n_626),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_654),
.A2(n_755),
.B(n_812),
.C(n_803),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_785),
.A2(n_543),
.B1(n_471),
.B2(n_491),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_738),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_714),
.A2(n_637),
.B(n_629),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_653),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_698),
.B(n_614),
.Y(n_979)
);

NOR2x2_ASAP7_75t_L g980 ( 
.A(n_738),
.B(n_252),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_744),
.B(n_290),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_698),
.B(n_637),
.Y(n_982)
);

NOR2x1_ASAP7_75t_L g983 ( 
.A(n_817),
.B(n_614),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_715),
.A2(n_637),
.B(n_629),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_746),
.B(n_626),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_785),
.A2(n_746),
.B(n_740),
.C(n_784),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_648),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_697),
.B(n_724),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_758),
.B(n_491),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_746),
.B(n_626),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_676),
.A2(n_543),
.B(n_637),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_654),
.A2(n_323),
.B1(n_296),
.B2(n_300),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_718),
.B(n_543),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_800),
.B(n_543),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_800),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_SL g996 ( 
.A(n_734),
.B(n_252),
.Y(n_996)
);

AO21x1_ASAP7_75t_L g997 ( 
.A1(n_804),
.A2(n_492),
.B(n_491),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_688),
.A2(n_816),
.B(n_801),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_664),
.B(n_463),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_787),
.A2(n_492),
.B(n_465),
.C(n_466),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_806),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_806),
.B(n_543),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_826),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_850),
.A2(n_723),
.B1(n_653),
.B2(n_773),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_866),
.B(n_744),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_860),
.B(n_689),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_823),
.A2(n_723),
.B(n_773),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_875),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_918),
.B(n_728),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_SL g1010 ( 
.A1(n_825),
.A2(n_788),
.B(n_791),
.C(n_802),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_995),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_850),
.B(n_733),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_891),
.B(n_799),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_880),
.B(n_719),
.Y(n_1014)
);

OA22x2_ASAP7_75t_L g1015 ( 
.A1(n_820),
.A2(n_794),
.B1(n_817),
.B2(n_326),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_818),
.B(n_722),
.Y(n_1016)
);

INVx3_ASAP7_75t_SL g1017 ( 
.A(n_980),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_872),
.A2(n_726),
.B(n_727),
.C(n_798),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_950),
.B(n_76),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_981),
.A2(n_817),
.B(n_788),
.C(n_802),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_1001),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_838),
.B(n_723),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_827),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_891),
.B(n_817),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_966),
.A2(n_773),
.B(n_723),
.C(n_815),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_978),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_830),
.A2(n_773),
.B1(n_710),
.B2(n_759),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_823),
.A2(n_791),
.B(n_807),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_838),
.B(n_648),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_826),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_844),
.B(n_648),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_892),
.B(n_807),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_844),
.B(n_648),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_832),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_892),
.B(n_815),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_858),
.A2(n_648),
.B(n_455),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_981),
.B(n_648),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_941),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_834),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_828),
.A2(n_492),
.B(n_455),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_822),
.B(n_292),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_SL g1042 ( 
.A(n_878),
.B(n_322),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_958),
.A2(n_466),
.B(n_465),
.C(n_460),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_978),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_903),
.B(n_906),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_863),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_837),
.A2(n_302),
.B1(n_304),
.B2(n_307),
.Y(n_1047)
);

AO21x2_ASAP7_75t_L g1048 ( 
.A1(n_868),
.A2(n_460),
.B(n_455),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_958),
.A2(n_466),
.B(n_465),
.C(n_460),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_841),
.A2(n_448),
.B(n_467),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_865),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_988),
.A2(n_471),
.B1(n_320),
.B2(n_318),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_836),
.A2(n_448),
.B(n_467),
.Y(n_1053)
);

AND2x4_ASAP7_75t_SL g1054 ( 
.A(n_978),
.B(n_463),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_967),
.B(n_311),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_974),
.A2(n_312),
.B(n_313),
.C(n_314),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_909),
.B(n_467),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_978),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_854),
.A2(n_467),
.B(n_78),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_946),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_842),
.A2(n_986),
.B(n_867),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_863),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_967),
.A2(n_328),
.B(n_467),
.C(n_25),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_835),
.B(n_23),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_968),
.B(n_24),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_974),
.A2(n_24),
.B(n_27),
.C(n_29),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_927),
.B(n_467),
.Y(n_1067)
);

O2A1O1Ixp5_ASAP7_75t_L g1068 ( 
.A1(n_997),
.A2(n_471),
.B(n_97),
.C(n_99),
.Y(n_1068)
);

BUFx8_ASAP7_75t_L g1069 ( 
.A(n_926),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_989),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_824),
.B(n_467),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_863),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_852),
.A2(n_467),
.B1(n_83),
.B2(n_169),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_927),
.B(n_471),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_851),
.B(n_863),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_976),
.B(n_154),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_910),
.A2(n_27),
.B(n_30),
.C(n_31),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_833),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_874),
.A2(n_30),
.B(n_31),
.C(n_33),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_848),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_989),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_896),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_930),
.B(n_33),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_925),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_930),
.B(n_471),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_970),
.B(n_34),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_907),
.A2(n_471),
.B1(n_37),
.B2(n_38),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_925),
.B(n_100),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_965),
.B(n_34),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_829),
.A2(n_106),
.B(n_149),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_L g1091 ( 
.A(n_845),
.B(n_992),
.C(n_846),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_925),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_913),
.B(n_38),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_925),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_923),
.B(n_42),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_938),
.A2(n_42),
.B(n_43),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_928),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_904),
.A2(n_115),
.B(n_148),
.Y(n_1098)
);

AO32x2_ASAP7_75t_L g1099 ( 
.A1(n_973),
.A2(n_43),
.A3(n_44),
.B1(n_50),
.B2(n_56),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_928),
.B(n_117),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_971),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_821),
.A2(n_44),
.B(n_50),
.C(n_57),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_855),
.B(n_57),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_934),
.B(n_130),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_928),
.B(n_839),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_888),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_890),
.B(n_60),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_890),
.B(n_61),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_883),
.A2(n_139),
.B(n_146),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_861),
.B(n_64),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_R g1111 ( 
.A(n_928),
.B(n_122),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_996),
.B(n_66),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_945),
.B(n_131),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_960),
.A2(n_140),
.B(n_142),
.C(n_150),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_SL g1115 ( 
.A(n_955),
.B(n_957),
.C(n_864),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_960),
.A2(n_961),
.B(n_884),
.C(n_999),
.Y(n_1116)
);

O2A1O1Ixp5_ASAP7_75t_L g1117 ( 
.A1(n_847),
.A2(n_840),
.B(n_999),
.C(n_859),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_921),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_895),
.A2(n_862),
.B(n_857),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_853),
.B(n_839),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_853),
.B(n_851),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_952),
.B(n_879),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_870),
.A2(n_914),
.B(n_877),
.Y(n_1123)
);

AOI22x1_ASAP7_75t_L g1124 ( 
.A1(n_998),
.A2(n_936),
.B1(n_939),
.B2(n_977),
.Y(n_1124)
);

NOR2x1_ASAP7_75t_L g1125 ( 
.A(n_948),
.B(n_952),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_983),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_851),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_882),
.A2(n_898),
.B(n_897),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_856),
.A2(n_949),
.B(n_943),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_851),
.B(n_987),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_993),
.A2(n_962),
.B(n_887),
.C(n_843),
.Y(n_1131)
);

NOR2x1_ASAP7_75t_R g1132 ( 
.A(n_955),
.B(n_957),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_919),
.B(n_975),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_869),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_886),
.B(n_908),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_979),
.A2(n_991),
.B(n_900),
.Y(n_1136)
);

BUFx4f_ASAP7_75t_L g1137 ( 
.A(n_819),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_905),
.A2(n_932),
.B(n_984),
.C(n_963),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_SL g1139 ( 
.A1(n_982),
.A2(n_972),
.B(n_915),
.C(n_900),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_819),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_894),
.B(n_912),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_889),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_SL g1143 ( 
.A(n_901),
.B(n_954),
.C(n_956),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1000),
.A2(n_915),
.B(n_899),
.C(n_893),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_959),
.B(n_964),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_931),
.B(n_947),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_937),
.B(n_940),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_935),
.A2(n_942),
.B(n_873),
.C(n_990),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_985),
.A2(n_1002),
.B(n_994),
.C(n_953),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_944),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_951),
.B(n_831),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_831),
.B(n_849),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1123),
.A2(n_876),
.B(n_944),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1039),
.B(n_972),
.Y(n_1154)
);

AOI221x1_ASAP7_75t_L g1155 ( 
.A1(n_1083),
.A2(n_911),
.B1(n_916),
.B2(n_885),
.C(n_920),
.Y(n_1155)
);

BUFx10_ASAP7_75t_L g1156 ( 
.A(n_1009),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1101),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1025),
.A2(n_902),
.A3(n_917),
.B(n_922),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1061),
.A2(n_924),
.A3(n_929),
.B(n_933),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1003),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1038),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1055),
.A2(n_871),
.B1(n_881),
.B2(n_1064),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_SL g1163 ( 
.A1(n_1037),
.A2(n_1012),
.B(n_1029),
.Y(n_1163)
);

AO32x2_ASAP7_75t_L g1164 ( 
.A1(n_1073),
.A2(n_1047),
.A3(n_1027),
.B1(n_1004),
.B2(n_1099),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1055),
.A2(n_1056),
.B(n_1020),
.C(n_1024),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1050),
.A2(n_1053),
.B(n_1129),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1119),
.A2(n_1128),
.B(n_1016),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1148),
.A2(n_1141),
.B(n_1036),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1038),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1023),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1067),
.A2(n_1018),
.B(n_1146),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1040),
.A2(n_1124),
.B(n_1028),
.Y(n_1172)
);

O2A1O1Ixp5_ASAP7_75t_SL g1173 ( 
.A1(n_1035),
.A2(n_1071),
.B(n_1110),
.C(n_1103),
.Y(n_1173)
);

AO21x1_ASAP7_75t_L g1174 ( 
.A1(n_1066),
.A2(n_1106),
.B(n_1114),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1087),
.A2(n_1005),
.B1(n_1014),
.B2(n_1142),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1092),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1041),
.B(n_1070),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_1138),
.A2(n_1131),
.A3(n_1079),
.B(n_1059),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1007),
.A2(n_1136),
.B(n_1117),
.Y(n_1179)
);

NOR4xp25_ASAP7_75t_L g1180 ( 
.A(n_1102),
.B(n_1096),
.C(n_1063),
.D(n_1077),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1081),
.B(n_1026),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1043),
.A2(n_1049),
.B(n_1144),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1134),
.B(n_1041),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1116),
.A2(n_1090),
.B(n_1151),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1109),
.A2(n_1145),
.B(n_1033),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1147),
.A2(n_1022),
.B(n_1010),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1031),
.A2(n_1135),
.B(n_1137),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1149),
.A2(n_1152),
.A3(n_1032),
.B(n_1074),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1127),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1069),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1098),
.A2(n_1075),
.B(n_1068),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_SL g1192 ( 
.A1(n_1133),
.A2(n_1076),
.B(n_1088),
.C(n_1100),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1137),
.A2(n_1143),
.B(n_1139),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1026),
.B(n_1091),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1013),
.A2(n_1042),
.B1(n_1009),
.B2(n_1112),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1085),
.A2(n_1089),
.A3(n_1095),
.B(n_1107),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_1142),
.A2(n_1115),
.B(n_1093),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_1008),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1108),
.A2(n_1019),
.B(n_1130),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1122),
.A2(n_1118),
.B(n_1125),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1013),
.A2(n_1091),
.B(n_1006),
.C(n_1113),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1121),
.A2(n_1105),
.B(n_1048),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1030),
.B(n_1069),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1087),
.A2(n_1052),
.B(n_1065),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1086),
.A2(n_1115),
.B(n_1126),
.C(n_1051),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1086),
.B(n_1120),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_1045),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1127),
.B(n_1060),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1017),
.A2(n_1045),
.B(n_1080),
.C(n_1082),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1046),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1015),
.A2(n_1078),
.B1(n_1034),
.B2(n_1021),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_L g1212 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1140),
.A2(n_1150),
.B1(n_1011),
.B2(n_1044),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1046),
.A2(n_1094),
.B(n_1072),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1017),
.A2(n_1072),
.B1(n_1044),
.B2(n_1058),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1084),
.A2(n_1097),
.B(n_1132),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1140),
.A2(n_1044),
.B1(n_1058),
.B2(n_1062),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1104),
.A2(n_1111),
.B(n_1054),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1140),
.A2(n_1062),
.B(n_1058),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1140),
.A2(n_1058),
.B1(n_1062),
.B2(n_1099),
.Y(n_1220)
);

NOR2xp67_ASAP7_75t_SL g1221 ( 
.A(n_1062),
.B(n_1099),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1099),
.A2(n_1083),
.B(n_1055),
.C(n_766),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1127),
.B(n_851),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1092),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1101),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1057),
.A2(n_1123),
.B(n_828),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1134),
.B(n_891),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1123),
.A2(n_1053),
.B(n_1050),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1008),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_1079),
.A2(n_652),
.B(n_656),
.C(n_1077),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1014),
.B(n_496),
.Y(n_1234)
);

AOI211x1_ASAP7_75t_L g1235 ( 
.A1(n_1006),
.A2(n_522),
.B(n_1096),
.C(n_652),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_1009),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1117),
.A2(n_1025),
.B(n_1036),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1083),
.A2(n_522),
.B(n_766),
.C(n_530),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1025),
.A2(n_997),
.A3(n_1061),
.B(n_1138),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1101),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1014),
.B(n_496),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1025),
.A2(n_997),
.A3(n_1061),
.B(n_1138),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1134),
.B(n_891),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_1083),
.A2(n_652),
.B(n_1056),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1083),
.A2(n_850),
.B1(n_540),
.B2(n_652),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1011),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1014),
.B(n_496),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1025),
.A2(n_997),
.A3(n_1061),
.B(n_1138),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1249)
);

AOI21xp33_ASAP7_75t_L g1250 ( 
.A1(n_1083),
.A2(n_766),
.B(n_850),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1003),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1127),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1003),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1079),
.A2(n_652),
.B(n_656),
.C(n_1077),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1014),
.B(n_496),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1123),
.A2(n_1053),
.B(n_1050),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1003),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1123),
.A2(n_1053),
.B(n_1050),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1039),
.B(n_875),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1057),
.A2(n_1123),
.B(n_828),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1014),
.B(n_496),
.Y(n_1263)
);

NOR4xp25_ASAP7_75t_L g1264 ( 
.A(n_1102),
.B(n_1083),
.C(n_1066),
.D(n_1079),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1123),
.A2(n_1053),
.B(n_1050),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1003),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1005),
.B(n_674),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1083),
.A2(n_850),
.B1(n_540),
.B2(n_652),
.Y(n_1268)
);

AOI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1057),
.A2(n_1123),
.B(n_828),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1014),
.B(n_496),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1101),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1083),
.A2(n_1055),
.B(n_766),
.C(n_530),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1092),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1117),
.A2(n_1025),
.B(n_1036),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1070),
.B(n_1081),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1131),
.A2(n_858),
.B(n_868),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1123),
.A2(n_1053),
.B(n_1050),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1123),
.A2(n_1053),
.B(n_1050),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1003),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1123),
.A2(n_1053),
.B(n_1050),
.Y(n_1281)
);

NAND2x1p5_ASAP7_75t_L g1282 ( 
.A(n_1127),
.B(n_851),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_SL g1283 ( 
.A(n_1044),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1083),
.A2(n_522),
.B1(n_850),
.B2(n_1055),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1083),
.A2(n_850),
.B1(n_540),
.B2(n_652),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1101),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1014),
.B(n_496),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1003),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1055),
.A2(n_649),
.B1(n_650),
.B2(n_528),
.Y(n_1290)
);

NAND3x1_ASAP7_75t_L g1291 ( 
.A(n_1112),
.B(n_423),
.C(n_1013),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1123),
.A2(n_735),
.B(n_969),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1005),
.B(n_674),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1011),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1011),
.Y(n_1295)
);

OAI22x1_ASAP7_75t_L g1296 ( 
.A1(n_1083),
.A2(n_1013),
.B1(n_1055),
.B2(n_1024),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1083),
.A2(n_1055),
.B(n_766),
.C(n_530),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1005),
.B(n_674),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1041),
.B(n_660),
.Y(n_1299)
);

AOI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1083),
.A2(n_522),
.B1(n_527),
.B2(n_604),
.C(n_1055),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1101),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1101),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1267),
.B(n_1293),
.Y(n_1303)
);

INVx4_ASAP7_75t_L g1304 ( 
.A(n_1283),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1284),
.A2(n_1300),
.B1(n_1250),
.B2(n_1290),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1160),
.Y(n_1306)
);

INVx6_ASAP7_75t_L g1307 ( 
.A(n_1176),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1194),
.Y(n_1308)
);

BUFx8_ASAP7_75t_SL g1309 ( 
.A(n_1198),
.Y(n_1309)
);

INVx6_ASAP7_75t_L g1310 ( 
.A(n_1176),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1284),
.A2(n_1250),
.B1(n_1296),
.B2(n_1245),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1245),
.A2(n_1268),
.B1(n_1285),
.B2(n_1183),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1176),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1156),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1157),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1231),
.Y(n_1316)
);

CKINVDCx11_ASAP7_75t_R g1317 ( 
.A(n_1156),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1207),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1299),
.B(n_1177),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1225),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1261),
.Y(n_1321)
);

BUFx8_ASAP7_75t_L g1322 ( 
.A(n_1283),
.Y(n_1322)
);

BUFx10_ASAP7_75t_L g1323 ( 
.A(n_1224),
.Y(n_1323)
);

AOI21xp33_ASAP7_75t_L g1324 ( 
.A1(n_1238),
.A2(n_1297),
.B(n_1273),
.Y(n_1324)
);

BUFx10_ASAP7_75t_L g1325 ( 
.A(n_1224),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1224),
.Y(n_1326)
);

CKINVDCx14_ASAP7_75t_R g1327 ( 
.A(n_1190),
.Y(n_1327)
);

BUFx8_ASAP7_75t_L g1328 ( 
.A(n_1274),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1252),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1240),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1274),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1267),
.B(n_1293),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1280),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1268),
.A2(n_1285),
.B1(n_1195),
.B2(n_1298),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1298),
.B(n_1234),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1204),
.A2(n_1243),
.B1(n_1229),
.B2(n_1206),
.Y(n_1336)
);

CKINVDCx11_ASAP7_75t_R g1337 ( 
.A(n_1236),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1241),
.A2(n_1247),
.B1(n_1287),
.B2(n_1271),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1256),
.B(n_1263),
.Y(n_1339)
);

BUFx4f_ASAP7_75t_SL g1340 ( 
.A(n_1274),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1161),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1272),
.Y(n_1342)
);

INVx4_ASAP7_75t_L g1343 ( 
.A(n_1181),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1175),
.A2(n_1174),
.B1(n_1244),
.B2(n_1194),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1236),
.Y(n_1345)
);

BUFx12f_ASAP7_75t_L g1346 ( 
.A(n_1207),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1201),
.A2(n_1291),
.B1(n_1222),
.B2(n_1165),
.Y(n_1347)
);

BUFx12f_ASAP7_75t_L g1348 ( 
.A(n_1259),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1266),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1175),
.A2(n_1277),
.B1(n_1162),
.B2(n_1168),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1235),
.B(n_1276),
.Y(n_1351)
);

INVx6_ASAP7_75t_L g1352 ( 
.A(n_1181),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1288),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1254),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1276),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1154),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1169),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1218),
.A2(n_1205),
.B1(n_1204),
.B2(n_1162),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1210),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1208),
.A2(n_1218),
.B1(n_1203),
.B2(n_1215),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1286),
.Y(n_1361)
);

BUFx8_ASAP7_75t_SL g1362 ( 
.A(n_1246),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1214),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1215),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1216),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1277),
.A2(n_1221),
.B1(n_1197),
.B2(n_1301),
.Y(n_1366)
);

BUFx10_ASAP7_75t_L g1367 ( 
.A(n_1302),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1216),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1197),
.A2(n_1170),
.B1(n_1211),
.B2(n_1171),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1294),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1295),
.Y(n_1371)
);

CKINVDCx11_ASAP7_75t_R g1372 ( 
.A(n_1217),
.Y(n_1372)
);

CKINVDCx11_ASAP7_75t_R g1373 ( 
.A(n_1217),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1187),
.A2(n_1200),
.B1(n_1208),
.B2(n_1186),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1193),
.A2(n_1213),
.B1(n_1199),
.B2(n_1220),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1213),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1220),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1212),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1264),
.A2(n_1182),
.B1(n_1184),
.B2(n_1180),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1264),
.A2(n_1180),
.B1(n_1275),
.B2(n_1237),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1209),
.A2(n_1292),
.B1(n_1289),
.B2(n_1226),
.Y(n_1381)
);

CKINVDCx14_ASAP7_75t_R g1382 ( 
.A(n_1189),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1212),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1223),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1237),
.A2(n_1275),
.B1(n_1249),
.B2(n_1270),
.Y(n_1385)
);

CKINVDCx8_ASAP7_75t_R g1386 ( 
.A(n_1163),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1155),
.A2(n_1253),
.B1(n_1257),
.B2(n_1233),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1219),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1228),
.A2(n_1251),
.B1(n_1164),
.B2(n_1191),
.Y(n_1389)
);

BUFx10_ASAP7_75t_L g1390 ( 
.A(n_1282),
.Y(n_1390)
);

BUFx4f_ASAP7_75t_SL g1391 ( 
.A(n_1192),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1164),
.A2(n_1255),
.B1(n_1232),
.B2(n_1185),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1188),
.B(n_1196),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1202),
.A2(n_1167),
.B1(n_1153),
.B2(n_1227),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1188),
.B(n_1196),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1173),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1196),
.Y(n_1397)
);

BUFx4f_ASAP7_75t_SL g1398 ( 
.A(n_1178),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1164),
.A2(n_1179),
.B1(n_1279),
.B2(n_1278),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1188),
.Y(n_1400)
);

AOI22x1_ASAP7_75t_L g1401 ( 
.A1(n_1178),
.A2(n_1242),
.B1(n_1248),
.B2(n_1239),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1172),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1230),
.A2(n_1281),
.B1(n_1265),
.B2(n_1260),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1258),
.A2(n_1166),
.B1(n_1178),
.B2(n_1239),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1242),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1262),
.A2(n_1269),
.B1(n_1242),
.B2(n_1248),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1158),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1158),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1159),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1159),
.A2(n_1284),
.B1(n_1300),
.B2(n_1083),
.Y(n_1410)
);

AOI22x1_ASAP7_75t_L g1411 ( 
.A1(n_1159),
.A2(n_1296),
.B1(n_880),
.B2(n_1193),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1284),
.A2(n_1297),
.B1(n_1273),
.B2(n_1290),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1160),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1284),
.A2(n_1300),
.B1(n_1083),
.B2(n_1250),
.Y(n_1414)
);

BUFx10_ASAP7_75t_L g1415 ( 
.A(n_1231),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1194),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1284),
.A2(n_1300),
.B1(n_1083),
.B2(n_1250),
.Y(n_1417)
);

INVx8_ASAP7_75t_L g1418 ( 
.A(n_1283),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1231),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1284),
.A2(n_1300),
.B1(n_1083),
.B2(n_1250),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1198),
.Y(n_1421)
);

INVx8_ASAP7_75t_L g1422 ( 
.A(n_1283),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1284),
.A2(n_1296),
.B1(n_1183),
.B2(n_1300),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1198),
.Y(n_1424)
);

CKINVDCx11_ASAP7_75t_R g1425 ( 
.A(n_1198),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1284),
.A2(n_1297),
.B1(n_1273),
.B2(n_1290),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1381),
.B(n_1363),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1393),
.B(n_1395),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1398),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1371),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1359),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1319),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1312),
.B(n_1311),
.Y(n_1433)
);

AO21x1_ASAP7_75t_L g1434 ( 
.A1(n_1347),
.A2(n_1426),
.B(n_1412),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1377),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1333),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1363),
.B(n_1408),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1400),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1311),
.B(n_1410),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1410),
.B(n_1334),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1391),
.A2(n_1358),
.B1(n_1365),
.B2(n_1368),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1335),
.B(n_1303),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1308),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1403),
.A2(n_1385),
.B(n_1401),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1403),
.A2(n_1385),
.B(n_1404),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1354),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1405),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1329),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1414),
.A2(n_1417),
.B1(n_1420),
.B2(n_1305),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1409),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1397),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1356),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1363),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1376),
.A2(n_1351),
.B(n_1332),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1407),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1402),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1407),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1367),
.Y(n_1458)
);

AOI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1339),
.A2(n_1378),
.B(n_1383),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1342),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1341),
.Y(n_1461)
);

OAI21xp33_ASAP7_75t_SL g1462 ( 
.A1(n_1414),
.A2(n_1420),
.B(n_1417),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1407),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1411),
.A2(n_1374),
.B(n_1379),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1315),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1320),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1330),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1416),
.B(n_1344),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1374),
.A2(n_1379),
.B(n_1350),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1406),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1375),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1370),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1366),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1350),
.A2(n_1380),
.B(n_1366),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1380),
.Y(n_1475)
);

BUFx10_ASAP7_75t_L g1476 ( 
.A(n_1318),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1392),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1399),
.Y(n_1478)
);

AO31x2_ASAP7_75t_L g1479 ( 
.A1(n_1389),
.A2(n_1324),
.A3(n_1387),
.B(n_1394),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1336),
.B(n_1338),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1386),
.Y(n_1481)
);

INVx5_ASAP7_75t_SL g1482 ( 
.A(n_1372),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1305),
.B(n_1369),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1369),
.B(n_1364),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1361),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1396),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1367),
.Y(n_1487)
);

CKINVDCx11_ASAP7_75t_R g1488 ( 
.A(n_1424),
.Y(n_1488)
);

BUFx2_ASAP7_75t_SL g1489 ( 
.A(n_1388),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1423),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1338),
.B(n_1321),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1372),
.A2(n_1373),
.B1(n_1355),
.B2(n_1360),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1390),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1309),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1390),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1341),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1384),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1373),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1329),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1499),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1478),
.B(n_1357),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1478),
.B(n_1467),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1496),
.B(n_1306),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1496),
.B(n_1306),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1449),
.A2(n_1327),
.B1(n_1382),
.B2(n_1304),
.Y(n_1505)
);

AND2x4_ASAP7_75t_SL g1506 ( 
.A(n_1461),
.B(n_1415),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1460),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1430),
.B(n_1419),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1462),
.A2(n_1413),
.B(n_1382),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1480),
.A2(n_1304),
.B(n_1421),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1453),
.Y(n_1511)
);

AO32x2_ASAP7_75t_L g1512 ( 
.A1(n_1458),
.A2(n_1343),
.A3(n_1326),
.B1(n_1362),
.B2(n_1345),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1433),
.A2(n_1422),
.B(n_1418),
.C(n_1327),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1467),
.B(n_1352),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1473),
.B(n_1346),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1489),
.B(n_1309),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1460),
.Y(n_1517)
);

OR2x6_ASAP7_75t_L g1518 ( 
.A(n_1427),
.B(n_1422),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1473),
.B(n_1346),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1465),
.B(n_1345),
.Y(n_1520)
);

O2A1O1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1434),
.A2(n_1316),
.B(n_1362),
.C(n_1317),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1463),
.B(n_1326),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1491),
.B(n_1418),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1466),
.B(n_1314),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1489),
.B(n_1425),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1432),
.B(n_1425),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1460),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1442),
.B(n_1422),
.Y(n_1528)
);

OR2x6_ASAP7_75t_L g1529 ( 
.A(n_1427),
.B(n_1418),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1436),
.B(n_1424),
.Y(n_1530)
);

AO32x2_ASAP7_75t_L g1531 ( 
.A1(n_1458),
.A2(n_1443),
.A3(n_1435),
.B1(n_1428),
.B2(n_1454),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1492),
.A2(n_1307),
.B1(n_1310),
.B2(n_1313),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1452),
.B(n_1322),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1428),
.B(n_1317),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1441),
.A2(n_1337),
.B(n_1314),
.Y(n_1535)
);

AOI221xp5_ASAP7_75t_L g1536 ( 
.A1(n_1434),
.A2(n_1433),
.B1(n_1490),
.B2(n_1439),
.C(n_1486),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1446),
.B(n_1322),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1490),
.B(n_1322),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1427),
.A2(n_1384),
.B(n_1337),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1431),
.Y(n_1540)
);

BUFx8_ASAP7_75t_SL g1541 ( 
.A(n_1494),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1448),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1427),
.B(n_1353),
.Y(n_1543)
);

INVx5_ASAP7_75t_L g1544 ( 
.A(n_1437),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1469),
.A2(n_1328),
.B(n_1340),
.C(n_1313),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1488),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1481),
.A2(n_1307),
.B1(n_1310),
.B2(n_1313),
.Y(n_1547)
);

A2O1A1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1469),
.A2(n_1328),
.B(n_1331),
.C(n_1310),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1463),
.B(n_1457),
.Y(n_1549)
);

INVx6_ASAP7_75t_SL g1550 ( 
.A(n_1476),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1484),
.B(n_1348),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1481),
.B(n_1348),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1482),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1440),
.A2(n_1349),
.B1(n_1353),
.B2(n_1331),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1483),
.A2(n_1323),
.B(n_1325),
.Y(n_1555)
);

A2O1A1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1483),
.A2(n_1440),
.B(n_1439),
.C(n_1474),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_SL g1557 ( 
.A(n_1459),
.B(n_1437),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1475),
.B(n_1484),
.Y(n_1558)
);

AOI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1459),
.A2(n_1454),
.B(n_1451),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1475),
.B(n_1470),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1485),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1486),
.B(n_1472),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_SL g1563 ( 
.A1(n_1485),
.A2(n_1477),
.B(n_1487),
.Y(n_1563)
);

AO21x2_ASAP7_75t_L g1564 ( 
.A1(n_1444),
.A2(n_1445),
.B(n_1464),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1470),
.B(n_1456),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1536),
.A2(n_1471),
.B1(n_1535),
.B2(n_1509),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1565),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1507),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1558),
.B(n_1435),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1515),
.B(n_1487),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1511),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1544),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1517),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1517),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1527),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1565),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1527),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1564),
.B(n_1450),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1502),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_L g1582 ( 
.A(n_1543),
.B(n_1451),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1561),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1559),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1518),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1560),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1514),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1515),
.B(n_1519),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1510),
.A2(n_1477),
.B1(n_1482),
.B2(n_1474),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1549),
.B(n_1518),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1514),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1557),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1556),
.B(n_1438),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1500),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1556),
.B(n_1450),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1575),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1573),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1568),
.B(n_1540),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1596),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1575),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1573),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1521),
.C(n_1519),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1590),
.B(n_1520),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1596),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1590),
.B(n_1520),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1576),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1576),
.Y(n_1610)
);

AOI221xp5_ASAP7_75t_L g1611 ( 
.A1(n_1567),
.A2(n_1505),
.B1(n_1538),
.B2(n_1498),
.C(n_1501),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1574),
.B(n_1593),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1569),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1594),
.B(n_1524),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1577),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1592),
.B(n_1525),
.C(n_1516),
.D(n_1534),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1594),
.B(n_1524),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1566),
.B(n_1571),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1595),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1578),
.B(n_1479),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1592),
.A2(n_1545),
.B(n_1548),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1578),
.B(n_1518),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1597),
.B(n_1518),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1589),
.B(n_1447),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1570),
.B(n_1479),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1595),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1598),
.A2(n_1482),
.B1(n_1501),
.B2(n_1468),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1579),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1591),
.B(n_1553),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1572),
.A2(n_1468),
.B1(n_1482),
.B2(n_1498),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1573),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1598),
.A2(n_1482),
.B1(n_1468),
.B2(n_1551),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1597),
.B(n_1529),
.Y(n_1634)
);

OR2x6_ASAP7_75t_SL g1635 ( 
.A(n_1595),
.B(n_1523),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1597),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1579),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1593),
.B(n_1529),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1612),
.B(n_1574),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1599),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1599),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1612),
.B(n_1600),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1585),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1603),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1603),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1635),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1619),
.B(n_1566),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1602),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1609),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1619),
.B(n_1566),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1602),
.B(n_1571),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1609),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1610),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1571),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1635),
.B(n_1583),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1610),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1615),
.Y(n_1658)
);

NAND2x1p5_ASAP7_75t_L g1659 ( 
.A(n_1621),
.B(n_1582),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1607),
.B(n_1585),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1604),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1615),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1622),
.A2(n_1584),
.B(n_1583),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1620),
.B(n_1627),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1620),
.B(n_1583),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1626),
.B(n_1588),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1616),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1616),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1629),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1629),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1612),
.B(n_1574),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1613),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1621),
.B(n_1580),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1625),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1627),
.B(n_1584),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1637),
.Y(n_1676)
);

AND2x2_ASAP7_75t_SL g1677 ( 
.A(n_1611),
.B(n_1584),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1626),
.B(n_1581),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1640),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1640),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1669),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1669),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1646),
.B(n_1655),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1643),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1641),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1677),
.A2(n_1605),
.B1(n_1611),
.B2(n_1622),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1646),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1641),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1644),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1677),
.A2(n_1605),
.B1(n_1546),
.B2(n_1553),
.Y(n_1690)
);

NAND2xp33_ASAP7_75t_SL g1691 ( 
.A(n_1655),
.B(n_1546),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1655),
.B(n_1612),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1677),
.B(n_1606),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1664),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1643),
.B(n_1606),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1644),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1660),
.B(n_1608),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1666),
.B(n_1601),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1645),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1639),
.B(n_1541),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1645),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1649),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1660),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1674),
.B(n_1608),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1649),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1664),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1656),
.B(n_1638),
.Y(n_1707)
);

AND2x2_ASAP7_75t_SL g1708 ( 
.A(n_1639),
.B(n_1506),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1663),
.A2(n_1617),
.B1(n_1630),
.B2(n_1636),
.C(n_1633),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1674),
.B(n_1614),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1652),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1652),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1664),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1653),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1666),
.B(n_1601),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1639),
.B(n_1617),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1663),
.B(n_1614),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1639),
.B(n_1638),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1656),
.B(n_1618),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1653),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1656),
.A2(n_1572),
.B1(n_1591),
.B2(n_1618),
.C(n_1542),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1685),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1685),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1688),
.Y(n_1724)
);

INVxp67_ASAP7_75t_SL g1725 ( 
.A(n_1716),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1688),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1687),
.B(n_1673),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1683),
.B(n_1639),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1689),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1700),
.B(n_1541),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1693),
.B(n_1698),
.Y(n_1731)
);

OAI21xp33_ASAP7_75t_L g1732 ( 
.A1(n_1686),
.A2(n_1628),
.B(n_1633),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1703),
.B(n_1709),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_SL g1734 ( 
.A(n_1690),
.B(n_1587),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1689),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1684),
.B(n_1648),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1683),
.B(n_1708),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1721),
.B(n_1648),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1708),
.B(n_1671),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1692),
.B(n_1671),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1696),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1695),
.B(n_1648),
.Y(n_1742)
);

AND2x2_ASAP7_75t_SL g1743 ( 
.A(n_1717),
.B(n_1506),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1707),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1697),
.B(n_1651),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1707),
.B(n_1704),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1692),
.B(n_1671),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1691),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1691),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1718),
.B(n_1671),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1710),
.B(n_1651),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1698),
.B(n_1673),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1718),
.A2(n_1671),
.B1(n_1631),
.B2(n_1587),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1696),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1715),
.B(n_1673),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_L g1756 ( 
.A(n_1679),
.B(n_1530),
.C(n_1533),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1680),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1737),
.B(n_1718),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1722),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1722),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1744),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_SL g1762 ( 
.A1(n_1725),
.A2(n_1651),
.B1(n_1659),
.B2(n_1719),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1733),
.B(n_1719),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1732),
.A2(n_1682),
.B(n_1681),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1748),
.A2(n_1631),
.B1(n_1628),
.B2(n_1659),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1728),
.Y(n_1766)
);

NAND4xp25_ASAP7_75t_L g1767 ( 
.A(n_1749),
.B(n_1513),
.C(n_1554),
.D(n_1526),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1723),
.Y(n_1768)
);

AOI21xp33_ASAP7_75t_L g1769 ( 
.A1(n_1734),
.A2(n_1706),
.B(n_1694),
.Y(n_1769)
);

INVxp67_ASAP7_75t_SL g1770 ( 
.A(n_1737),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1738),
.A2(n_1659),
.B(n_1699),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1723),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1726),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1726),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1743),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1743),
.A2(n_1694),
.B1(n_1713),
.B2(n_1706),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1728),
.B(n_1740),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1757),
.B(n_1713),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1739),
.A2(n_1587),
.B1(n_1543),
.B2(n_1529),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1756),
.B(n_1715),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1744),
.B(n_1701),
.Y(n_1781)
);

AOI21xp33_ASAP7_75t_L g1782 ( 
.A1(n_1731),
.A2(n_1720),
.B(n_1711),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1735),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1758),
.B(n_1739),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1761),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1777),
.Y(n_1786)
);

AOI21xp33_ASAP7_75t_L g1787 ( 
.A1(n_1770),
.A2(n_1727),
.B(n_1731),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1759),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1763),
.B(n_1746),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1764),
.B(n_1727),
.Y(n_1790)
);

AOI21xp33_ASAP7_75t_L g1791 ( 
.A1(n_1775),
.A2(n_1736),
.B(n_1729),
.Y(n_1791)
);

NAND4xp25_ASAP7_75t_L g1792 ( 
.A(n_1780),
.B(n_1753),
.C(n_1730),
.D(n_1750),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1766),
.B(n_1740),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1758),
.B(n_1750),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1766),
.B(n_1747),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1776),
.A2(n_1747),
.B(n_1513),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1762),
.A2(n_1659),
.B1(n_1742),
.B2(n_1751),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1777),
.B(n_1745),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1771),
.A2(n_1741),
.B1(n_1724),
.B2(n_1735),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1759),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1782),
.A2(n_1754),
.B1(n_1755),
.B2(n_1752),
.C(n_1702),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1773),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_SL g1803 ( 
.A1(n_1778),
.A2(n_1755),
.B1(n_1752),
.B2(n_1754),
.C(n_1545),
.Y(n_1803)
);

AOI322xp5_ASAP7_75t_L g1804 ( 
.A1(n_1790),
.A2(n_1769),
.A3(n_1774),
.B1(n_1760),
.B2(n_1772),
.C1(n_1768),
.C2(n_1783),
.Y(n_1804)
);

NAND2xp67_ASAP7_75t_SL g1805 ( 
.A(n_1801),
.B(n_1665),
.Y(n_1805)
);

OAI322xp33_ASAP7_75t_L g1806 ( 
.A1(n_1802),
.A2(n_1783),
.A3(n_1760),
.B1(n_1768),
.B2(n_1772),
.C1(n_1781),
.C2(n_1765),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1792),
.B(n_1767),
.Y(n_1807)
);

AOI33xp33_ASAP7_75t_L g1808 ( 
.A1(n_1799),
.A2(n_1785),
.A3(n_1786),
.B1(n_1784),
.B2(n_1794),
.B3(n_1798),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1789),
.B(n_1779),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1788),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1784),
.Y(n_1811)
);

XOR2xp5_ASAP7_75t_L g1812 ( 
.A(n_1797),
.B(n_1532),
.Y(n_1812)
);

INVxp67_ASAP7_75t_L g1813 ( 
.A(n_1793),
.Y(n_1813)
);

OAI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1791),
.A2(n_1543),
.B1(n_1550),
.B2(n_1636),
.Y(n_1814)
);

NOR4xp25_ASAP7_75t_L g1815 ( 
.A(n_1802),
.B(n_1720),
.C(n_1711),
.D(n_1537),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1787),
.B(n_1796),
.Y(n_1816)
);

OAI321xp33_ASAP7_75t_L g1817 ( 
.A1(n_1807),
.A2(n_1803),
.A3(n_1799),
.B1(n_1795),
.B2(n_1800),
.C(n_1547),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1811),
.B(n_1705),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1810),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1816),
.A2(n_1809),
.B1(n_1805),
.B2(n_1813),
.Y(n_1820)
);

NAND3xp33_ASAP7_75t_L g1821 ( 
.A(n_1804),
.B(n_1803),
.C(n_1714),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_SL g1822 ( 
.A(n_1808),
.B(n_1815),
.C(n_1812),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_L g1823 ( 
.A(n_1806),
.B(n_1552),
.C(n_1508),
.Y(n_1823)
);

AOI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1814),
.A2(n_1539),
.B(n_1548),
.C(n_1528),
.Y(n_1824)
);

NAND5xp2_ASAP7_75t_L g1825 ( 
.A(n_1814),
.B(n_1555),
.C(n_1455),
.D(n_1634),
.E(n_1624),
.Y(n_1825)
);

OAI211xp5_ASAP7_75t_L g1826 ( 
.A1(n_1804),
.A2(n_1582),
.B(n_1712),
.C(n_1497),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1811),
.B(n_1665),
.Y(n_1827)
);

O2A1O1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1822),
.A2(n_1661),
.B(n_1672),
.C(n_1654),
.Y(n_1828)
);

O2A1O1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1817),
.A2(n_1661),
.B(n_1672),
.C(n_1654),
.Y(n_1829)
);

NAND5xp2_ASAP7_75t_L g1830 ( 
.A(n_1820),
.B(n_1826),
.C(n_1823),
.D(n_1827),
.E(n_1818),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1821),
.A2(n_1586),
.B1(n_1665),
.B2(n_1675),
.C(n_1672),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_SL g1832 ( 
.A(n_1824),
.B(n_1476),
.C(n_1624),
.Y(n_1832)
);

AOI321xp33_ASAP7_75t_L g1833 ( 
.A1(n_1828),
.A2(n_1819),
.A3(n_1825),
.B1(n_1586),
.B2(n_1642),
.C(n_1493),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1830),
.A2(n_1642),
.B1(n_1675),
.B2(n_1654),
.C(n_1670),
.Y(n_1834)
);

O2A1O1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1831),
.A2(n_1661),
.B(n_1675),
.C(n_1642),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1829),
.B(n_1642),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1832),
.A2(n_1642),
.B1(n_1676),
.B2(n_1670),
.C(n_1668),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1831),
.B(n_1657),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1836),
.B(n_1678),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1834),
.A2(n_1476),
.B1(n_1497),
.B2(n_1634),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1835),
.A2(n_1497),
.B(n_1661),
.Y(n_1841)
);

NAND4xp75_ASAP7_75t_L g1842 ( 
.A(n_1837),
.B(n_1838),
.C(n_1833),
.D(n_1493),
.Y(n_1842)
);

OAI211xp5_ASAP7_75t_L g1843 ( 
.A1(n_1833),
.A2(n_1497),
.B(n_1476),
.C(n_1495),
.Y(n_1843)
);

AOI322xp5_ASAP7_75t_L g1844 ( 
.A1(n_1840),
.A2(n_1650),
.A3(n_1647),
.B1(n_1623),
.B2(n_1667),
.C1(n_1657),
.C2(n_1668),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1843),
.A2(n_1495),
.B(n_1676),
.C(n_1667),
.Y(n_1845)
);

NAND4xp75_ASAP7_75t_L g1846 ( 
.A(n_1841),
.B(n_1647),
.C(n_1650),
.D(n_1662),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1845),
.A2(n_1839),
.B(n_1842),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1847),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1848),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1848),
.A2(n_1846),
.B1(n_1844),
.B2(n_1550),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1849),
.A2(n_1550),
.B1(n_1543),
.B2(n_1512),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1850),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1852),
.A2(n_1662),
.B1(n_1658),
.B2(n_1600),
.C(n_1632),
.Y(n_1853)
);

OA21x2_ASAP7_75t_L g1854 ( 
.A1(n_1851),
.A2(n_1658),
.B(n_1650),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1854),
.A2(n_1504),
.B(n_1503),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1855),
.B(n_1853),
.Y(n_1856)
);

OAI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1678),
.B1(n_1600),
.B2(n_1632),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1637),
.B1(n_1563),
.B2(n_1522),
.C(n_1632),
.Y(n_1858)
);

AOI211xp5_ASAP7_75t_L g1859 ( 
.A1(n_1858),
.A2(n_1429),
.B(n_1522),
.C(n_1455),
.Y(n_1859)
);


endmodule