module fake_jpeg_14239_n_63 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_21),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_17),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_0),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_28),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_26),
.B1(n_29),
.B2(n_33),
.Y(n_36)
);

OAI22x1_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_40),
.B1(n_20),
.B2(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_1),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_1),
.B(n_2),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_26),
.B1(n_28),
.B2(n_11),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_24),
.C(n_23),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_47),
.C(n_49),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_40),
.B1(n_4),
.B2(n_5),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_2),
.B(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_53),
.C(n_43),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_3),
.B(n_4),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.C(n_58),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_7),
.B(n_8),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_9),
.C(n_10),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_51),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_53),
.B(n_52),
.Y(n_62)
);

OAI321xp33_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_50),
.A3(n_14),
.B1(n_15),
.B2(n_8),
.C(n_7),
.Y(n_63)
);


endmodule