module fake_jpeg_3204_n_473 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_473);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_473;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx8_ASAP7_75t_SL g39 ( 
.A(n_6),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_41),
.B(n_77),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_51),
.Y(n_101)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_47),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_50),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_27),
.B(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_64),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_70),
.Y(n_132)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_13),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_36),
.Y(n_81)
);

INVx2_ASAP7_75t_R g136 ( 
.A(n_81),
.Y(n_136)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_84),
.Y(n_149)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_20),
.B(n_13),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_20),
.Y(n_111)
);

INVx8_ASAP7_75t_SL g87 ( 
.A(n_26),
.Y(n_87)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_103),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_142),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_111),
.A2(n_18),
.B(n_17),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_29),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_146),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_75),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_42),
.A2(n_16),
.B1(n_20),
.B2(n_37),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_37),
.B1(n_30),
.B2(n_16),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_80),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_74),
.B(n_78),
.C(n_89),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_82),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_69),
.B(n_22),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_22),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_158),
.B(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_168),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_116),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_120),
.B(n_30),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_171),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_182),
.Y(n_221)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_179),
.Y(n_210)
);

CKINVDCx12_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_174),
.Y(n_206)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_178),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_109),
.B(n_31),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_177),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_101),
.B(n_18),
.Y(n_178)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_181),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g182 ( 
.A(n_102),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_184),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_186),
.Y(n_212)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_188),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_126),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_101),
.B(n_91),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_104),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_102),
.A2(n_47),
.B(n_71),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_149),
.B(n_126),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_193),
.B1(n_139),
.B2(n_125),
.Y(n_195)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_195),
.A2(n_166),
.B1(n_179),
.B2(n_185),
.Y(n_244)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_132),
.A3(n_117),
.B1(n_141),
.B2(n_122),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_224),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_133),
.C(n_127),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_131),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_153),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_169),
.B(n_161),
.Y(n_242)
);

NOR2x1p5_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_149),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_108),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_220),
.A2(n_163),
.B(n_181),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_231),
.B(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_177),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_229),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_228),
.Y(n_264)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_176),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_212),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_219),
.B(n_225),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_156),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_241),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_154),
.B1(n_155),
.B2(n_186),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_202),
.B1(n_212),
.B2(n_223),
.Y(n_258)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_212),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_119),
.B1(n_118),
.B2(n_145),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_240),
.A2(n_192),
.B1(n_160),
.B2(n_165),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_193),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_164),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_250),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_244),
.A2(n_247),
.B1(n_83),
.B2(n_84),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_204),
.B(n_199),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_223),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_202),
.A2(n_104),
.B1(n_95),
.B2(n_173),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

AND2x6_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_180),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_213),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_255),
.A2(n_271),
.B(n_254),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_272),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_203),
.C(n_206),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_268),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_261),
.A2(n_237),
.B1(n_216),
.B2(n_232),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_246),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_241),
.B(n_223),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_270),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_215),
.C(n_208),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_207),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_243),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_210),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_210),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_210),
.B1(n_196),
.B2(n_214),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_240),
.B1(n_238),
.B2(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_279),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_252),
.A2(n_245),
.B1(n_250),
.B2(n_242),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_280),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_282),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_298),
.B1(n_301),
.B2(n_270),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_250),
.B1(n_231),
.B2(n_229),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_287),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_285),
.B(n_290),
.Y(n_322)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_255),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_288),
.A2(n_264),
.B1(n_256),
.B2(n_213),
.Y(n_318)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_214),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_293),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_L g294 ( 
.A1(n_259),
.A2(n_229),
.B(n_235),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_272),
.Y(n_315)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_201),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_296),
.B(n_264),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_299),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_259),
.A2(n_267),
.B1(n_257),
.B2(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_300),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_267),
.A2(n_249),
.B1(n_194),
.B2(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_276),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_280),
.A2(n_257),
.B1(n_254),
.B2(n_265),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_306),
.A2(n_283),
.B1(n_292),
.B2(n_284),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_255),
.B(n_264),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_291),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_310),
.A2(n_318),
.B1(n_321),
.B2(n_297),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_311),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_315),
.A2(n_327),
.B(n_328),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_299),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_148),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_268),
.C(n_274),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_292),
.C(n_284),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_301),
.A2(n_261),
.B1(n_256),
.B2(n_276),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_287),
.Y(n_329)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_215),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_180),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_201),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_278),
.B(n_249),
.Y(n_328)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_329),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_310),
.A2(n_281),
.B1(n_278),
.B2(n_298),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_322),
.B(n_281),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_332),
.B(n_338),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_333),
.A2(n_335),
.B1(n_339),
.B2(n_345),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_326),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_336),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_328),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_304),
.A2(n_284),
.B1(n_279),
.B2(n_295),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_340),
.A2(n_325),
.B(n_317),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g341 ( 
.A(n_306),
.B(n_289),
.CI(n_300),
.CON(n_341),
.SN(n_341)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_347),
.Y(n_359)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_305),
.Y(n_342)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_322),
.B(n_307),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_344),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_319),
.A2(n_302),
.B1(n_188),
.B2(n_184),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_228),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_319),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_316),
.A2(n_228),
.B1(n_135),
.B2(n_125),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_228),
.C(n_134),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_350),
.C(n_308),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_228),
.C(n_183),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_351),
.B(n_312),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_324),
.Y(n_352)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_353),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_355),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_363),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_333),
.A2(n_304),
.B1(n_321),
.B2(n_311),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_362),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_309),
.Y(n_360)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_309),
.C(n_307),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_339),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_349),
.C(n_351),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_365),
.C(n_362),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_346),
.B(n_303),
.C(n_323),
.Y(n_365)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_368),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_303),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_372),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_373),
.A2(n_303),
.B1(n_325),
.B2(n_317),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_330),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_209),
.B(n_135),
.Y(n_390)
);

AO22x1_ASAP7_75t_L g378 ( 
.A1(n_367),
.A2(n_358),
.B1(n_370),
.B2(n_368),
.Y(n_378)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_364),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_397),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_314),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_385),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_369),
.B(n_345),
.C(n_314),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_347),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_388),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_341),
.C(n_145),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_341),
.Y(n_389)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_390),
.A2(n_137),
.B1(n_123),
.B2(n_62),
.Y(n_412)
);

AOI321xp33_ASAP7_75t_L g391 ( 
.A1(n_361),
.A2(n_209),
.A3(n_90),
.B1(n_76),
.B2(n_119),
.C(n_115),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_391),
.A2(n_49),
.B1(n_66),
.B2(n_60),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_128),
.C(n_45),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_393),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_128),
.C(n_44),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_373),
.A2(n_43),
.B(n_73),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_395),
.A2(n_379),
.B(n_386),
.Y(n_410)
);

FAx1_ASAP7_75t_SL g397 ( 
.A(n_365),
.B(n_137),
.CI(n_123),
.CON(n_397),
.SN(n_397)
);

BUFx24_ASAP7_75t_SL g398 ( 
.A(n_375),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_377),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_399),
.B(n_403),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_394),
.B(n_357),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g424 ( 
.A(n_402),
.B(n_392),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_355),
.C(n_366),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_359),
.C(n_360),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_408),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_359),
.C(n_372),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_409),
.B(n_414),
.Y(n_428)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_410),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_413),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_72),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_58),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_415),
.B(n_379),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_400),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_417),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_385),
.Y(n_417)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_404),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_419),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_380),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_420),
.B(n_422),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_407),
.B(n_388),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_408),
.B(n_411),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_423),
.B(n_50),
.Y(n_434)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_424),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_393),
.Y(n_426)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_426),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_400),
.A2(n_378),
.B(n_397),
.Y(n_430)
);

AOI21xp33_ASAP7_75t_L g435 ( 
.A1(n_430),
.A2(n_0),
.B(n_1),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_421),
.A2(n_402),
.B1(n_401),
.B2(n_53),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_434),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_439),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_48),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_436),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_32),
.C(n_2),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_0),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_441),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_2),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_442),
.B(n_440),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_427),
.C(n_430),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_445),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_433),
.B(n_429),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_450),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_437),
.B(n_2),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_448),
.B(n_453),
.Y(n_456)
);

AOI322xp5_ASAP7_75t_L g450 ( 
.A1(n_443),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_3),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_432),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_457),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_444),
.B(n_431),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_446),
.A2(n_436),
.B(n_439),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_459),
.A2(n_460),
.B(n_7),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_451),
.A2(n_3),
.B(n_4),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_458),
.A2(n_452),
.B(n_451),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_461),
.A2(n_7),
.B(n_9),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_11),
.C(n_8),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_463),
.C(n_11),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

NOR3xp33_ASAP7_75t_L g468 ( 
.A(n_465),
.B(n_464),
.C(n_10),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_466),
.B(n_467),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_9),
.C(n_10),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_469),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_470),
.C(n_9),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_472),
.B(n_11),
.Y(n_473)
);


endmodule