module real_jpeg_16242_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_432),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_0),
.B(n_433),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_1),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_1),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_1),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_1),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_1),
.B(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_2),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_3),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_3),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_3),
.Y(n_309)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_4),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_4),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_4),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_4),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_4),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_5),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_5),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_5),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_5),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_5),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_5),
.B(n_157),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_117),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_6),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_6),
.B(n_183),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_6),
.B(n_45),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_7),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_7),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_7),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_7),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_7),
.B(n_377),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_7),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_8),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_9),
.Y(n_168)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_9),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_10),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_11),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_12),
.B(n_39),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_12),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_12),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_12),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_12),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_12),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_12),
.B(n_302),
.Y(n_301)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_13),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_13),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_15),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_16),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_16),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_16),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_16),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_16),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g307 ( 
.A(n_16),
.B(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_17),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_392),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_345),
.B(n_390),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_194),
.B(n_342),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21x1_ASAP7_75t_L g342 ( 
.A1(n_23),
.A2(n_343),
.B(n_344),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_148),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_24),
.B(n_148),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_104),
.C(n_134),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_25),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_67),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_48),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_27),
.B(n_48),
.C(n_67),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_47),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_28),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_28),
.B(n_34),
.C(n_41),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_28),
.A2(n_47),
.B1(n_425),
.B2(n_428),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_35),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_35),
.B(n_117),
.Y(n_125)
);

NAND2x1_ASAP7_75t_L g182 ( 
.A(n_35),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_35),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_35),
.B(n_368),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_35),
.B(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_40),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_40),
.Y(n_223)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_49),
.B(n_60),
.C(n_65),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.C(n_56),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_56),
.B(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_64),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_82),
.C(n_93),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_68),
.B(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_77),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

MAJx3_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_74),
.C(n_77),
.Y(n_147)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_73),
.Y(n_240)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_79),
.Y(n_427)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_80),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_81),
.B(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_84),
.A2(n_125),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_161),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_84),
.A2(n_125),
.B(n_155),
.Y(n_373)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_85),
.Y(n_285)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_85),
.Y(n_300)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_91),
.Y(n_322)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.C(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_94),
.A2(n_100),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_94),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_95),
.B(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_99),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_100),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_100),
.A2(n_209),
.B1(n_239),
.B2(n_370),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_101),
.Y(n_316)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_104),
.B(n_135),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_122),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_105),
.B(n_109),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_107),
.B(n_381),
.C(n_384),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_115),
.B(n_121),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_117),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_129),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_123),
.A2(n_124),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_124),
.B(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_125),
.B(n_247),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_125),
.A2(n_162),
.B1(n_239),
.B2(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_125),
.B(n_367),
.C(n_370),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_126),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_144),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_145),
.C(n_147),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_140),
.C(n_143),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_143),
.B(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_149),
.B(n_151),
.C(n_389),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_176),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_163),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_153),
.B(n_154),
.C(n_164),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_162),
.B(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_165),
.B(n_170),
.C(n_361),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_168),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_168),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_174),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_176),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_177),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_180),
.B(n_182),
.C(n_186),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_190),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_191),
.B(n_348),
.C(n_349),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_192),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_226),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_224),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_197),
.B(n_224),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.C(n_205),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_198),
.A2(n_199),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_201),
.A2(n_202),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_211),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.C(n_222),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_212),
.A2(n_213),
.B1(n_222),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_215),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI21x1_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_333),
.B(n_341),
.Y(n_227)
);

AOI21x1_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_278),
.B(n_332),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_254),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_230),
.B(n_254),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_252),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_232),
.B(n_236),
.C(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.C(n_246),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_239),
.Y(n_370)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_256),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_252),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_275),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_275),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.C(n_271),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_267),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_294),
.B(n_331),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_292),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_292),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.C(n_290),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_283),
.A2(n_290),
.B1(n_291),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_286),
.Y(n_304)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_325),
.B(n_330),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_313),
.B(n_324),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_303),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_297),
.B(n_303),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_301),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_307),
.C(n_310),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_318),
.B(n_323),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_317),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_317),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_339),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_339),
.Y(n_341)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_388),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_346),
.B(n_388),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.Y(n_346)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_365),
.B1(n_386),
.B2(n_387),
.Y(n_350)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_362),
.C(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_353)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_354),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_354),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_360),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_356),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_359),
.C(n_360),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_357),
.A2(n_358),
.B1(n_406),
.B2(n_410),
.Y(n_405)
);

INVx3_ASAP7_75t_SL g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_365),
.B(n_386),
.C(n_430),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_371),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_372),
.C(n_374),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_381),
.B1(n_384),
.B2(n_385),
.Y(n_375)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_376),
.Y(n_384)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_381),
.Y(n_385)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_R g392 ( 
.A(n_393),
.B(n_431),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_429),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_429),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_411),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_406),
.Y(n_410)
);

INVx3_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx8_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2x2_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_420),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_419),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_422),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_425),
.Y(n_428)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);


endmodule