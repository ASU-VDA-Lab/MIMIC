module fake_jpeg_18342_n_304 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx2_ASAP7_75t_SL g74 ( 
.A(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_51),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_21),
.B1(n_22),
.B2(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_28),
.B1(n_33),
.B2(n_16),
.Y(n_92)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_26),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_22),
.B1(n_41),
.B2(n_19),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_65),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_90),
.B1(n_81),
.B2(n_83),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_32),
.B1(n_31),
.B2(n_19),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_75),
.B1(n_85),
.B2(n_65),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_19),
.B1(n_32),
.B2(n_30),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_17),
.C(n_42),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_17),
.C(n_90),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_30),
.B1(n_33),
.B2(n_27),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_40),
.B1(n_29),
.B2(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_52),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_17),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_60),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_28),
.B1(n_49),
.B2(n_55),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_61),
.B(n_64),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_107),
.B(n_108),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_45),
.B1(n_62),
.B2(n_55),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_45),
.B1(n_62),
.B2(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_105),
.B1(n_71),
.B2(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_101),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_45),
.B1(n_62),
.B2(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_53),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_43),
.B1(n_53),
.B2(n_59),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_90),
.C(n_70),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_50),
.B(n_59),
.C(n_44),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_60),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_24),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_24),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_85),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_25),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_116),
.C(n_118),
.Y(n_154)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_140),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_95),
.B1(n_102),
.B2(n_107),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_126),
.B(n_139),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_77),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_90),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_84),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_135),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_89),
.B1(n_74),
.B2(n_44),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_138),
.B(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_80),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_83),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_89),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_83),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_104),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_89),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_50),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_25),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_152),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_175),
.C(n_24),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_127),
.B1(n_129),
.B2(n_135),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_94),
.B1(n_116),
.B2(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_168),
.B1(n_144),
.B2(n_124),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_158),
.A2(n_169),
.B(n_171),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_118),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_123),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_97),
.B(n_119),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_166),
.B(n_174),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_95),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_167),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_165),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_97),
.B(n_119),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_128),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_94),
.B1(n_105),
.B2(n_96),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_109),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_66),
.B(n_109),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_121),
.A2(n_88),
.B(n_79),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_100),
.C(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_100),
.B(n_16),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_29),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_132),
.B(n_122),
.C(n_137),
.D(n_131),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_170),
.B(n_177),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_137),
.B1(n_144),
.B2(n_132),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_159),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_191),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_122),
.B1(n_145),
.B2(n_141),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_161),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_203),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_192),
.C(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_143),
.B1(n_29),
.B2(n_24),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_170),
.B(n_8),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_195),
.B(n_13),
.Y(n_217)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_8),
.C(n_15),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_12),
.B(n_14),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_0),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_167),
.B1(n_152),
.B2(n_173),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_206),
.A2(n_224),
.B1(n_204),
.B2(n_199),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_151),
.C(n_154),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_192),
.C(n_180),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_215),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_212),
.B(n_218),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_195),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_158),
.B(n_153),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_227),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_166),
.B(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_171),
.B(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_169),
.B(n_151),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_228),
.B1(n_200),
.B2(n_1),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_155),
.B(n_173),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_188),
.A2(n_169),
.B(n_150),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_229),
.B1(n_182),
.B2(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_159),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_238),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_234),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_186),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_207),
.B(n_160),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_191),
.C(n_183),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_237),
.A2(n_209),
.B1(n_216),
.B2(n_213),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_181),
.C(n_201),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_193),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_245),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_200),
.C(n_7),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_216),
.C(n_217),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_213),
.B1(n_224),
.B2(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_253),
.B1(n_252),
.B2(n_258),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_256),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_220),
.B1(n_221),
.B2(n_226),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_212),
.C(n_225),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_SL g257 ( 
.A1(n_240),
.A2(n_218),
.B(n_206),
.C(n_228),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_229),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_260),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_235),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_222),
.C(n_221),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_244),
.C(n_238),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_239),
.C(n_247),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_222),
.C(n_248),
.Y(n_269)
);

OAI221xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_232),
.B1(n_209),
.B2(n_246),
.C(n_9),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_12),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_6),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_267),
.A2(n_251),
.B1(n_254),
.B2(n_3),
.Y(n_275)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_275),
.Y(n_287)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_254),
.B(n_6),
.C(n_9),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_14),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_269),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_281),
.Y(n_292)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_11),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_0),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_11),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_0),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_286),
.Y(n_293)
);

OAI322xp33_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_268),
.A3(n_271),
.B1(n_274),
.B2(n_6),
.C1(n_11),
.C2(n_4),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_292),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_291),
.A2(n_277),
.B(n_281),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_280),
.C(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.C(n_280),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_299),
.Y(n_301)
);

OAI311xp33_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_276),
.A3(n_288),
.B1(n_291),
.C1(n_2),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_298),
.C(n_300),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_297),
.Y(n_304)
);


endmodule