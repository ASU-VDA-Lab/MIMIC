module fake_jpeg_13569_n_206 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_206);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_90),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_70),
.Y(n_93)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_79),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_104),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_62),
.B1(n_67),
.B2(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_64),
.B1(n_60),
.B2(n_2),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_62),
.B1(n_55),
.B2(n_72),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_102),
.B1(n_64),
.B2(n_71),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_55),
.B1(n_72),
.B2(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_61),
.B1(n_82),
.B2(n_80),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_61),
.B1(n_99),
.B2(n_98),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_78),
.C(n_65),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_73),
.B(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_64),
.Y(n_115)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_123),
.B(n_111),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_57),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_116),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_73),
.B(n_70),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_95),
.B(n_60),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_59),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_0),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_7),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_68),
.B1(n_72),
.B2(n_71),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_135),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_136),
.B(n_7),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_25),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_15),
.C(n_16),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_110),
.B(n_118),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_1),
.B(n_3),
.C(n_5),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_13),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_11),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_164)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_6),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_29),
.B1(n_54),
.B2(n_53),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_33),
.B(n_49),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_11),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_26),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_168),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_156),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_164),
.B1(n_137),
.B2(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_31),
.B1(n_37),
.B2(n_42),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_160),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_8),
.B(n_10),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_18),
.B(n_22),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_145),
.B1(n_131),
.B2(n_136),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_153),
.B1(n_163),
.B2(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_163),
.Y(n_175)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_38),
.C(n_47),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_148),
.C(n_168),
.Y(n_172)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_170),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_173),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_134),
.B1(n_17),
.B2(n_16),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_183),
.B1(n_176),
.B2(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_179),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_158),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_23),
.C(n_27),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_186),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_191),
.B1(n_175),
.B2(n_172),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_167),
.B(n_155),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_184),
.Y(n_194)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_175),
.A2(n_162),
.B1(n_157),
.B2(n_46),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_162),
.B1(n_177),
.B2(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_199),
.A2(n_195),
.B(n_185),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_200),
.A2(n_193),
.B(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_192),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_196),
.C(n_194),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_198),
.B(n_188),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_204),
.A2(n_190),
.B1(n_171),
.B2(n_184),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_205),
.B(n_43),
.Y(n_206)
);


endmodule