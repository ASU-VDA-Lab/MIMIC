module fake_jpeg_25793_n_91 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_91);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_4),
.B(n_10),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_49),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_58),
.B1(n_59),
.B2(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_23),
.B(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_6),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_42),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_60),
.C(n_61),
.Y(n_64)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_15),
.B1(n_7),
.B2(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_42),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_27),
.C(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_66),
.B(n_45),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_33),
.B1(n_30),
.B2(n_45),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_61),
.B1(n_45),
.B2(n_38),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_73),
.B1(n_69),
.B2(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_57),
.B(n_53),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_51),
.B1(n_44),
.B2(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_60),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_78),
.C(n_76),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_64),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_80),
.B1(n_68),
.B2(n_75),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_66),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_84),
.B(n_79),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_80),
.B(n_81),
.C(n_82),
.Y(n_87)
);

AOI322xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_88),
.A3(n_85),
.B1(n_67),
.B2(n_46),
.C1(n_35),
.C2(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_74),
.B1(n_33),
.B2(n_56),
.Y(n_88)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_28),
.A3(n_35),
.B1(n_39),
.B2(n_37),
.C1(n_29),
.C2(n_55),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_68),
.B1(n_28),
.B2(n_13),
.Y(n_91)
);


endmodule