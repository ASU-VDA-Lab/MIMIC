module real_aes_16197_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1044;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1768;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_1712;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_1749;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1691;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
XNOR2xp5_ASAP7_75t_L g936 ( .A(n_0), .B(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1446 ( .A1(n_0), .A2(n_92), .B1(n_1413), .B2(n_1418), .Y(n_1446) );
INVx1_ASAP7_75t_L g665 ( .A(n_1), .Y(n_665) );
INVx1_ASAP7_75t_L g557 ( .A(n_2), .Y(n_557) );
INVx1_ASAP7_75t_L g360 ( .A(n_3), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_3), .B(n_370), .Y(n_567) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_3), .B(n_244), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_3), .B(n_385), .Y(n_1691) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_4), .A2(n_249), .B1(n_445), .B2(n_449), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_4), .A2(n_190), .B1(n_516), .B2(n_519), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g1336 ( .A(n_5), .Y(n_1336) );
INVx1_ASAP7_75t_L g1379 ( .A(n_6), .Y(n_1379) );
OAI22xp5_ASAP7_75t_SL g1393 ( .A1(n_7), .A2(n_216), .B1(n_926), .B2(n_1175), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_7), .A2(n_216), .B1(n_645), .B2(n_985), .Y(n_1396) );
INVx1_ASAP7_75t_L g1309 ( .A(n_8), .Y(n_1309) );
OAI22xp33_ASAP7_75t_SL g1348 ( .A1(n_9), .A2(n_331), .B1(n_614), .B2(n_1349), .Y(n_1348) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_9), .A2(n_174), .B1(n_491), .B2(n_586), .Y(n_1361) );
INVx1_ASAP7_75t_L g1260 ( .A(n_10), .Y(n_1260) );
INVx1_ASAP7_75t_L g1368 ( .A(n_11), .Y(n_1368) );
INVx1_ASAP7_75t_L g428 ( .A(n_12), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_12), .A2(n_249), .B1(n_519), .B2(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g1310 ( .A1(n_13), .A2(n_143), .B1(n_362), .B2(n_641), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1312 ( .A1(n_13), .A2(n_143), .B1(n_586), .B2(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g681 ( .A(n_14), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_15), .Y(n_1217) );
OAI22xp33_ASAP7_75t_L g1394 ( .A1(n_16), .A2(n_142), .B1(n_362), .B2(n_641), .Y(n_1394) );
OAI22xp33_ASAP7_75t_L g1402 ( .A1(n_16), .A2(n_142), .B1(n_659), .B2(n_1202), .Y(n_1402) );
AOI22xp33_ASAP7_75t_SL g1668 ( .A1(n_17), .A2(n_213), .B1(n_1669), .B2(n_1670), .Y(n_1668) );
INVxp67_ASAP7_75t_SL g1717 ( .A(n_17), .Y(n_1717) );
CKINVDCx5p33_ASAP7_75t_R g1742 ( .A(n_18), .Y(n_1742) );
OAI22xp5_ASAP7_75t_L g1192 ( .A1(n_19), .A2(n_305), .B1(n_771), .B2(n_1175), .Y(n_1192) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_19), .A2(n_305), .B1(n_760), .B2(n_1136), .Y(n_1195) );
INVx2_ASAP7_75t_L g471 ( .A(n_20), .Y(n_471) );
INVx1_ASAP7_75t_L g1014 ( .A(n_21), .Y(n_1014) );
INVx1_ASAP7_75t_L g1010 ( .A(n_22), .Y(n_1010) );
INVx1_ASAP7_75t_L g1102 ( .A(n_23), .Y(n_1102) );
INVx1_ASAP7_75t_L g1073 ( .A(n_24), .Y(n_1073) );
INVx1_ASAP7_75t_L g1255 ( .A(n_25), .Y(n_1255) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_26), .A2(n_88), .B1(n_702), .B2(n_993), .C(n_995), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_26), .A2(n_43), .B1(n_1043), .B2(n_1045), .Y(n_1042) );
INVx1_ASAP7_75t_L g735 ( .A(n_27), .Y(n_735) );
AOI22xp33_ASAP7_75t_SL g1284 ( .A1(n_28), .A2(n_160), .B1(n_449), .B2(n_1285), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_28), .A2(n_199), .B1(n_723), .B2(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g890 ( .A(n_29), .Y(n_890) );
INVx1_ASAP7_75t_L g1097 ( .A(n_30), .Y(n_1097) );
OAI211xp5_ASAP7_75t_L g1123 ( .A1(n_31), .A2(n_625), .B(n_1124), .C(n_1127), .Y(n_1123) );
INVx1_ASAP7_75t_L g1134 ( .A(n_31), .Y(n_1134) );
INVx1_ASAP7_75t_L g781 ( .A(n_32), .Y(n_781) );
OAI221xp5_ASAP7_75t_L g585 ( .A1(n_33), .A2(n_87), .B1(n_477), .B2(n_586), .C(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g610 ( .A(n_33), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_34), .A2(n_309), .B1(n_612), .B2(n_865), .Y(n_1238) );
OAI22xp33_ASAP7_75t_L g1248 ( .A1(n_34), .A2(n_309), .B1(n_477), .B2(n_483), .Y(n_1248) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_35), .Y(n_355) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_35), .B(n_353), .Y(n_1414) );
CKINVDCx5p33_ASAP7_75t_R g1630 ( .A(n_36), .Y(n_1630) );
INVx1_ASAP7_75t_L g949 ( .A(n_37), .Y(n_949) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_38), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g1445 ( .A1(n_39), .A2(n_67), .B1(n_1421), .B2(n_1430), .Y(n_1445) );
INVx1_ASAP7_75t_L g1391 ( .A(n_40), .Y(n_1391) );
INVx1_ASAP7_75t_L g1156 ( .A(n_41), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_42), .A2(n_180), .B1(n_749), .B2(n_750), .Y(n_748) );
OAI22xp33_ASAP7_75t_L g765 ( .A1(n_42), .A2(n_180), .B1(n_362), .B2(n_382), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g998 ( .A1(n_43), .A2(n_72), .B1(n_702), .B2(n_993), .C(n_999), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1666 ( .A1(n_44), .A2(n_277), .B1(n_514), .B2(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1712 ( .A(n_44), .Y(n_1712) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_45), .A2(n_263), .B1(n_614), .B2(n_615), .Y(n_1239) );
OAI22xp33_ASAP7_75t_SL g1241 ( .A1(n_45), .A2(n_263), .B1(n_491), .B2(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g914 ( .A(n_46), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_46), .A2(n_337), .B1(n_636), .B2(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g758 ( .A(n_47), .Y(n_758) );
OAI211xp5_ASAP7_75t_L g766 ( .A1(n_47), .A2(n_625), .B(n_767), .C(n_768), .Y(n_766) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_48), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_49), .Y(n_419) );
INVx1_ASAP7_75t_L g952 ( .A(n_50), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g1276 ( .A1(n_51), .A2(n_199), .B1(n_391), .B2(n_1277), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_51), .A2(n_160), .B1(n_1289), .B2(n_1290), .Y(n_1288) );
INVx1_ASAP7_75t_L g1004 ( .A(n_52), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_52), .A2(n_254), .B1(n_449), .B2(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g561 ( .A(n_53), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g1429 ( .A1(n_54), .A2(n_116), .B1(n_1421), .B2(n_1430), .Y(n_1429) );
AOI22xp5_ASAP7_75t_L g1437 ( .A1(n_55), .A2(n_255), .B1(n_1421), .B2(n_1430), .Y(n_1437) );
INVx1_ASAP7_75t_L g1654 ( .A(n_56), .Y(n_1654) );
INVx1_ASAP7_75t_L g882 ( .A(n_57), .Y(n_882) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_58), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g1080 ( .A(n_59), .Y(n_1080) );
INVx1_ASAP7_75t_L g1378 ( .A(n_60), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_61), .B(n_470), .Y(n_589) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_61), .Y(n_604) );
OAI211xp5_ASAP7_75t_L g1344 ( .A1(n_62), .A2(n_573), .B(n_598), .C(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1360 ( .A(n_62), .Y(n_1360) );
INVx1_ASAP7_75t_L g733 ( .A(n_63), .Y(n_733) );
INVx1_ASAP7_75t_L g1376 ( .A(n_64), .Y(n_1376) );
CKINVDCx5p33_ASAP7_75t_R g1328 ( .A(n_65), .Y(n_1328) );
OAI222xp33_ASAP7_75t_L g394 ( .A1(n_66), .A2(n_177), .B1(n_395), .B2(n_399), .C1(n_403), .C2(n_404), .Y(n_394) );
OAI222xp33_ASAP7_75t_L g458 ( .A1(n_66), .A2(n_177), .B1(n_217), .B2(n_459), .C1(n_467), .C2(n_473), .Y(n_458) );
INVx1_ASAP7_75t_L g1259 ( .A(n_68), .Y(n_1259) );
OAI22xp33_ASAP7_75t_L g1176 ( .A1(n_69), .A2(n_291), .B1(n_362), .B2(n_641), .Y(n_1176) );
OAI22xp33_ASAP7_75t_L g1178 ( .A1(n_69), .A2(n_291), .B1(n_659), .B2(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1126 ( .A(n_70), .Y(n_1126) );
OAI211xp5_ASAP7_75t_L g1132 ( .A1(n_70), .A2(n_648), .B(n_649), .C(n_1133), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_71), .A2(n_181), .B1(n_491), .B2(n_593), .Y(n_592) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_71), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_72), .A2(n_88), .B1(n_440), .B2(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g1304 ( .A(n_73), .Y(n_1304) );
AOI22xp33_ASAP7_75t_SL g1663 ( .A1(n_74), .A2(n_170), .B1(n_1011), .B2(n_1664), .Y(n_1663) );
INVxp67_ASAP7_75t_SL g1715 ( .A(n_74), .Y(n_1715) );
CKINVDCx5p33_ASAP7_75t_R g1751 ( .A(n_75), .Y(n_1751) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_76), .A2(n_167), .B1(n_760), .B2(n_761), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_76), .A2(n_167), .B1(n_636), .B2(n_771), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_77), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g1452 ( .A1(n_78), .A2(n_235), .B1(n_1421), .B2(n_1430), .Y(n_1452) );
OAI211xp5_ASAP7_75t_L g1233 ( .A1(n_79), .A2(n_598), .B(n_1234), .C(n_1235), .Y(n_1233) );
INVx1_ASAP7_75t_L g1245 ( .A(n_79), .Y(n_1245) );
AOI22xp5_ASAP7_75t_L g1412 ( .A1(n_80), .A2(n_243), .B1(n_1413), .B2(n_1418), .Y(n_1412) );
INVx1_ASAP7_75t_L g634 ( .A(n_81), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_81), .A2(n_648), .B(n_649), .C(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g559 ( .A(n_82), .Y(n_559) );
INVx1_ASAP7_75t_L g947 ( .A(n_83), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g1420 ( .A1(n_84), .A2(n_104), .B1(n_1421), .B2(n_1423), .Y(n_1420) );
INVx1_ASAP7_75t_L g1724 ( .A(n_84), .Y(n_1724) );
AOI22xp33_ASAP7_75t_L g1728 ( .A1(n_84), .A2(n_1729), .B1(n_1732), .B2(n_1771), .Y(n_1728) );
AO22x1_ASAP7_75t_L g1443 ( .A1(n_85), .A2(n_256), .B1(n_1413), .B2(n_1418), .Y(n_1443) );
XNOR2xp5_ASAP7_75t_L g835 ( .A(n_86), .B(n_836), .Y(n_835) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_87), .A2(n_181), .B1(n_614), .B2(n_615), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_89), .A2(n_188), .B1(n_477), .B2(n_491), .Y(n_1007) );
INVx1_ASAP7_75t_L g1020 ( .A(n_89), .Y(n_1020) );
INVx1_ASAP7_75t_L g1104 ( .A(n_90), .Y(n_1104) );
INVx1_ASAP7_75t_L g823 ( .A(n_91), .Y(n_823) );
OAI211xp5_ASAP7_75t_L g828 ( .A1(n_91), .A2(n_829), .B(n_831), .C(n_832), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g1758 ( .A1(n_93), .A2(n_261), .B1(n_612), .B2(n_614), .Y(n_1758) );
OAI22xp5_ASAP7_75t_SL g1766 ( .A1(n_93), .A2(n_128), .B1(n_483), .B2(n_491), .Y(n_1766) );
INVx1_ASAP7_75t_L g591 ( .A(n_94), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g1761 ( .A(n_95), .Y(n_1761) );
INVx1_ASAP7_75t_L g1263 ( .A(n_96), .Y(n_1263) );
CKINVDCx5p33_ASAP7_75t_R g1741 ( .A(n_97), .Y(n_1741) );
OAI22xp33_ASAP7_75t_L g1122 ( .A1(n_98), .A2(n_156), .B1(n_362), .B2(n_615), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_98), .A2(n_156), .B1(n_657), .B2(n_750), .Y(n_1131) );
CKINVDCx5p33_ASAP7_75t_R g1327 ( .A(n_99), .Y(n_1327) );
INVx1_ASAP7_75t_L g1015 ( .A(n_100), .Y(n_1015) );
AOI22xp33_ASAP7_75t_SL g1286 ( .A1(n_101), .A2(n_341), .B1(n_391), .B2(n_1277), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_101), .A2(n_102), .B1(n_1292), .B2(n_1295), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_102), .A2(n_311), .B1(n_449), .B2(n_1281), .Y(n_1280) );
XOR2xp5_ASAP7_75t_L g1322 ( .A(n_103), .B(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g950 ( .A(n_105), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_106), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g1748 ( .A(n_107), .Y(n_1748) );
OAI22xp33_ASAP7_75t_L g976 ( .A1(n_108), .A2(n_138), .B1(n_614), .B2(n_641), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_108), .A2(n_125), .B1(n_491), .B2(n_760), .Y(n_978) );
INVx1_ASAP7_75t_L g943 ( .A(n_109), .Y(n_943) );
INVx1_ASAP7_75t_L g1237 ( .A(n_110), .Y(n_1237) );
INVx1_ASAP7_75t_L g954 ( .A(n_111), .Y(n_954) );
INVx1_ASAP7_75t_L g1162 ( .A(n_112), .Y(n_1162) );
OAI211xp5_ASAP7_75t_L g818 ( .A1(n_113), .A2(n_598), .B(n_819), .C(n_820), .Y(n_818) );
INVx1_ASAP7_75t_L g833 ( .A(n_113), .Y(n_833) );
INVx1_ASAP7_75t_L g353 ( .A(n_114), .Y(n_353) );
INVx1_ASAP7_75t_L g1371 ( .A(n_115), .Y(n_1371) );
AO221x2_ASAP7_75t_L g1530 ( .A1(n_117), .A2(n_322), .B1(n_1413), .B2(n_1418), .C(n_1531), .Y(n_1530) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_118), .A2(n_288), .B1(n_637), .B2(n_641), .Y(n_825) );
OAI22xp33_ASAP7_75t_L g834 ( .A1(n_118), .A2(n_152), .B1(n_477), .B2(n_483), .Y(n_834) );
XOR2xp5_ASAP7_75t_L g378 ( .A(n_119), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g670 ( .A(n_120), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g1665 ( .A1(n_121), .A2(n_175), .B1(n_514), .B2(n_993), .Y(n_1665) );
INVx1_ASAP7_75t_L g1713 ( .A(n_121), .Y(n_1713) );
CKINVDCx5p33_ASAP7_75t_R g972 ( .A(n_122), .Y(n_972) );
INVx1_ASAP7_75t_L g1150 ( .A(n_123), .Y(n_1150) );
INVx1_ASAP7_75t_L g1076 ( .A(n_124), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_125), .A2(n_212), .B1(n_636), .B2(n_975), .Y(n_974) );
OAI22xp33_ASAP7_75t_SL g1763 ( .A1(n_126), .A2(n_128), .B1(n_615), .B2(n_865), .Y(n_1763) );
OAI22xp5_ASAP7_75t_L g1770 ( .A1(n_126), .A2(n_132), .B1(n_1358), .B2(n_1359), .Y(n_1770) );
INVx1_ASAP7_75t_L g1643 ( .A(n_127), .Y(n_1643) );
OAI222xp33_ASAP7_75t_L g1706 ( .A1(n_127), .A2(n_200), .B1(n_1707), .B2(n_1711), .C1(n_1714), .C2(n_1718), .Y(n_1706) );
INVx1_ASAP7_75t_L g1079 ( .A(n_129), .Y(n_1079) );
CKINVDCx5p33_ASAP7_75t_R g1213 ( .A(n_130), .Y(n_1213) );
INVx1_ASAP7_75t_L g731 ( .A(n_131), .Y(n_731) );
INVx1_ASAP7_75t_L g1762 ( .A(n_132), .Y(n_1762) );
INVx1_ASAP7_75t_L g1077 ( .A(n_133), .Y(n_1077) );
AOI31xp33_ASAP7_75t_L g989 ( .A1(n_134), .A2(n_990), .A3(n_1006), .B(n_1018), .Y(n_989) );
NAND2xp33_ASAP7_75t_SL g1035 ( .A(n_134), .B(n_1036), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g1048 ( .A(n_134), .Y(n_1048) );
AO22x1_ASAP7_75t_L g1434 ( .A1(n_134), .A2(n_326), .B1(n_1413), .B2(n_1418), .Y(n_1434) );
INVx1_ASAP7_75t_L g1099 ( .A(n_135), .Y(n_1099) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_136), .A2(n_182), .B1(n_641), .B2(n_865), .Y(n_864) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_136), .A2(n_173), .B1(n_477), .B2(n_483), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_137), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_138), .A2(n_212), .B1(n_659), .B2(n_985), .Y(n_984) );
CKINVDCx5p33_ASAP7_75t_R g1216 ( .A(n_139), .Y(n_1216) );
CKINVDCx5p33_ASAP7_75t_R g840 ( .A(n_140), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g1745 ( .A(n_141), .Y(n_1745) );
INVx1_ASAP7_75t_L g1106 ( .A(n_144), .Y(n_1106) );
CKINVDCx5p33_ASAP7_75t_R g1330 ( .A(n_145), .Y(n_1330) );
INVx1_ASAP7_75t_L g1683 ( .A(n_146), .Y(n_1683) );
OAI211xp5_ASAP7_75t_L g1169 ( .A1(n_147), .A2(n_767), .B(n_1170), .C(n_1171), .Y(n_1169) );
INVx1_ASAP7_75t_L g1182 ( .A(n_147), .Y(n_1182) );
INVx1_ASAP7_75t_L g945 ( .A(n_148), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_149), .Y(n_693) );
INVx1_ASAP7_75t_L g1172 ( .A(n_150), .Y(n_1172) );
INVx1_ASAP7_75t_L g1308 ( .A(n_151), .Y(n_1308) );
OAI22xp33_ASAP7_75t_L g824 ( .A1(n_152), .A2(n_265), .B1(n_614), .B2(n_639), .Y(n_824) );
INVx1_ASAP7_75t_L g862 ( .A(n_153), .Y(n_862) );
OAI211xp5_ASAP7_75t_L g868 ( .A1(n_153), .A2(n_829), .B(n_831), .C(n_869), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_154), .Y(n_787) );
AO22x1_ASAP7_75t_L g1441 ( .A1(n_155), .A2(n_327), .B1(n_1421), .B2(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g555 ( .A(n_157), .Y(n_555) );
CKINVDCx16_ASAP7_75t_R g1532 ( .A(n_158), .Y(n_1532) );
OAI211xp5_ASAP7_75t_SL g1389 ( .A1(n_159), .A2(n_625), .B(n_767), .C(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1401 ( .A(n_159), .Y(n_1401) );
INVx1_ASAP7_75t_L g1074 ( .A(n_161), .Y(n_1074) );
INVx1_ASAP7_75t_L g633 ( .A(n_162), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g1733 ( .A1(n_163), .A2(n_1734), .B1(n_1735), .B2(n_1736), .Y(n_1733) );
CKINVDCx5p33_ASAP7_75t_R g1734 ( .A(n_163), .Y(n_1734) );
OAI22xp5_ASAP7_75t_L g1174 ( .A1(n_164), .A2(n_284), .B1(n_771), .B2(n_1175), .Y(n_1174) );
OAI22xp33_ASAP7_75t_L g1183 ( .A1(n_164), .A2(n_284), .B1(n_760), .B2(n_761), .Y(n_1183) );
OAI211xp5_ASAP7_75t_L g859 ( .A1(n_165), .A2(n_598), .B(n_819), .C(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g870 ( .A(n_165), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g1333 ( .A(n_166), .Y(n_1333) );
INVx1_ASAP7_75t_L g1161 ( .A(n_168), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_169), .A2(n_245), .B1(n_636), .B2(n_638), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_169), .A2(n_245), .B1(n_645), .B2(n_646), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g1694 ( .A1(n_170), .A2(n_213), .B1(n_1695), .B2(n_1697), .C(n_1698), .Y(n_1694) );
OAI22xp33_ASAP7_75t_L g863 ( .A1(n_171), .A2(n_173), .B1(n_614), .B2(n_639), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g867 ( .A1(n_171), .A2(n_182), .B1(n_491), .B2(n_586), .Y(n_867) );
INVx1_ASAP7_75t_L g690 ( .A(n_172), .Y(n_690) );
OAI22xp33_ASAP7_75t_SL g1350 ( .A1(n_174), .A2(n_294), .B1(n_637), .B2(n_641), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1699 ( .A1(n_175), .A2(n_277), .B1(n_445), .B2(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g1145 ( .A(n_176), .Y(n_1145) );
INVx1_ASAP7_75t_L g1070 ( .A(n_178), .Y(n_1070) );
INVx2_ASAP7_75t_L g1416 ( .A(n_179), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_179), .B(n_1417), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_179), .B(n_290), .Y(n_1424) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_183), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g1747 ( .A(n_184), .Y(n_1747) );
INVx1_ASAP7_75t_L g680 ( .A(n_185), .Y(n_680) );
INVx1_ASAP7_75t_L g720 ( .A(n_186), .Y(n_720) );
XNOR2xp5_ASAP7_75t_L g1362 ( .A(n_187), .B(n_1363), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_188), .A2(n_271), .B1(n_612), .B2(n_865), .Y(n_1024) );
INVx1_ASAP7_75t_L g973 ( .A(n_189), .Y(n_973) );
OAI211xp5_ASAP7_75t_L g979 ( .A1(n_189), .A2(n_831), .B(n_980), .C(n_981), .Y(n_979) );
INVx1_ASAP7_75t_L g434 ( .A(n_190), .Y(n_434) );
XOR2xp5_ASAP7_75t_L g539 ( .A(n_191), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g917 ( .A(n_192), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g932 ( .A1(n_192), .A2(n_225), .B1(n_614), .B2(n_641), .Y(n_932) );
XNOR2x2_ASAP7_75t_L g1091 ( .A(n_193), .B(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g546 ( .A(n_194), .Y(n_546) );
INVx1_ASAP7_75t_L g1679 ( .A(n_195), .Y(n_1679) );
INVx1_ASAP7_75t_L g1057 ( .A(n_196), .Y(n_1057) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_197), .Y(n_796) );
INVx1_ASAP7_75t_L g1236 ( .A(n_198), .Y(n_1236) );
INVx1_ASAP7_75t_L g1648 ( .A(n_200), .Y(n_1648) );
XOR2x2_ASAP7_75t_L g1230 ( .A(n_201), .B(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1375 ( .A(n_202), .Y(n_1375) );
INVx1_ASAP7_75t_L g717 ( .A(n_203), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_204), .A2(n_382), .B(n_388), .C(n_408), .Y(n_381) );
INVx1_ASAP7_75t_L g492 ( .A(n_204), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g1189 ( .A(n_205), .Y(n_1189) );
INVx1_ASAP7_75t_L g1151 ( .A(n_206), .Y(n_1151) );
INVx1_ASAP7_75t_L g549 ( .A(n_207), .Y(n_549) );
INVx2_ASAP7_75t_L g501 ( .A(n_208), .Y(n_501) );
INVx1_ASAP7_75t_L g529 ( .A(n_208), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g1635 ( .A(n_208), .B(n_471), .Y(n_1635) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_209), .Y(n_788) );
XOR2xp5_ASAP7_75t_L g711 ( .A(n_210), .B(n_712), .Y(n_711) );
OAI22xp33_ASAP7_75t_L g1053 ( .A1(n_211), .A2(n_269), .B1(n_612), .B2(n_865), .Y(n_1053) );
OAI22xp5_ASAP7_75t_SL g1060 ( .A1(n_211), .A2(n_238), .B1(n_477), .B2(n_491), .Y(n_1060) );
INVx1_ASAP7_75t_L g892 ( .A(n_214), .Y(n_892) );
INVx1_ASAP7_75t_L g402 ( .A(n_215), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_215), .A2(n_242), .B1(n_477), .B2(n_483), .Y(n_476) );
INVx1_ASAP7_75t_L g390 ( .A(n_217), .Y(n_390) );
INVx1_ASAP7_75t_L g909 ( .A(n_218), .Y(n_909) );
OA211x2_ASAP7_75t_L g927 ( .A1(n_218), .A2(n_628), .B(n_673), .C(n_928), .Y(n_927) );
BUFx3_ASAP7_75t_L g466 ( .A(n_219), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_220), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_221), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g1214 ( .A(n_222), .Y(n_1214) );
OAI22xp5_ASAP7_75t_SL g875 ( .A1(n_223), .A2(n_876), .B1(n_923), .B2(n_934), .Y(n_875) );
NAND4xp25_ASAP7_75t_L g876 ( .A(n_223), .B(n_877), .C(n_894), .D(n_903), .Y(n_876) );
XOR2xp5_ASAP7_75t_L g1140 ( .A(n_224), .B(n_1141), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_224), .A2(n_226), .B1(n_1413), .B2(n_1418), .Y(n_1453) );
INVx1_ASAP7_75t_L g913 ( .A(n_225), .Y(n_913) );
INVx1_ASAP7_75t_L g1191 ( .A(n_227), .Y(n_1191) );
OAI211xp5_ASAP7_75t_L g1196 ( .A1(n_227), .A2(n_831), .B(n_1197), .C(n_1199), .Y(n_1196) );
INVx1_ASAP7_75t_L g1307 ( .A(n_228), .Y(n_1307) );
INVx1_ASAP7_75t_L g417 ( .A(n_229), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_229), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g1147 ( .A(n_230), .Y(n_1147) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_231), .Y(n_844) );
INVx1_ASAP7_75t_L g885 ( .A(n_232), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_233), .Y(n_792) );
INVx1_ASAP7_75t_L g729 ( .A(n_234), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_236), .A2(n_307), .B1(n_362), .B2(n_641), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_236), .A2(n_307), .B1(n_657), .B2(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g1056 ( .A(n_237), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_238), .A2(n_275), .B1(n_614), .B2(n_615), .Y(n_1058) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_239), .Y(n_1211) );
INVx1_ASAP7_75t_L g672 ( .A(n_240), .Y(n_672) );
INVx1_ASAP7_75t_L g1256 ( .A(n_241), .Y(n_1256) );
INVx1_ASAP7_75t_L g414 ( .A(n_242), .Y(n_414) );
BUFx3_ASAP7_75t_L g370 ( .A(n_244), .Y(n_370) );
INVx1_ASAP7_75t_L g385 ( .A(n_244), .Y(n_385) );
INVx1_ASAP7_75t_L g1125 ( .A(n_246), .Y(n_1125) );
CKINVDCx20_ASAP7_75t_R g1534 ( .A(n_247), .Y(n_1534) );
AOI22xp5_ASAP7_75t_L g1436 ( .A1(n_248), .A2(n_262), .B1(n_1413), .B2(n_1418), .Y(n_1436) );
INVx1_ASAP7_75t_L g545 ( .A(n_250), .Y(n_545) );
INVx1_ASAP7_75t_L g908 ( .A(n_251), .Y(n_908) );
INVx1_ASAP7_75t_L g893 ( .A(n_252), .Y(n_893) );
INVx1_ASAP7_75t_L g1252 ( .A(n_253), .Y(n_1252) );
AOI22xp5_ASAP7_75t_L g991 ( .A1(n_254), .A2(n_280), .B1(n_537), .B2(n_911), .Y(n_991) );
INVx1_ASAP7_75t_L g1109 ( .A(n_257), .Y(n_1109) );
INVx1_ASAP7_75t_L g716 ( .A(n_258), .Y(n_716) );
OAI211xp5_ASAP7_75t_L g1054 ( .A1(n_259), .A2(n_598), .B(n_673), .C(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1065 ( .A(n_259), .Y(n_1065) );
CKINVDCx5p33_ASAP7_75t_R g1331 ( .A(n_260), .Y(n_1331) );
NOR2xp33_ASAP7_75t_L g1765 ( .A(n_261), .B(n_477), .Y(n_1765) );
CKINVDCx5p33_ASAP7_75t_R g1750 ( .A(n_264), .Y(n_1750) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_265), .A2(n_288), .B1(n_491), .B2(n_586), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g1334 ( .A(n_266), .Y(n_1334) );
INVx1_ASAP7_75t_L g889 ( .A(n_267), .Y(n_889) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_268), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g1066 ( .A1(n_269), .A2(n_275), .B1(n_483), .B2(n_586), .Y(n_1066) );
XOR2x2_ASAP7_75t_L g1272 ( .A(n_270), .B(n_1273), .Y(n_1272) );
AOI22xp5_ASAP7_75t_L g1428 ( .A1(n_270), .A2(n_335), .B1(n_1413), .B2(n_1418), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g1016 ( .A1(n_271), .A2(n_310), .B1(n_483), .B2(n_586), .Y(n_1016) );
INVx1_ASAP7_75t_L g1305 ( .A(n_272), .Y(n_1305) );
AO22x1_ASAP7_75t_L g1433 ( .A1(n_273), .A2(n_279), .B1(n_1421), .B2(n_1430), .Y(n_1433) );
INVx1_ASAP7_75t_L g464 ( .A(n_274), .Y(n_464) );
INVx1_ASAP7_75t_L g482 ( .A(n_274), .Y(n_482) );
INVx1_ASAP7_75t_L g1108 ( .A(n_276), .Y(n_1108) );
INVx1_ASAP7_75t_L g1101 ( .A(n_278), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_280), .A2(n_313), .B1(n_440), .B2(n_1040), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1128 ( .A1(n_281), .A2(n_325), .B1(n_636), .B2(n_926), .Y(n_1128) );
OAI22xp33_ASAP7_75t_L g1135 ( .A1(n_281), .A2(n_325), .B1(n_760), .B2(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g886 ( .A(n_282), .Y(n_886) );
OAI211xp5_ASAP7_75t_L g751 ( .A1(n_283), .A2(n_649), .B(n_752), .C(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g769 ( .A(n_283), .Y(n_769) );
INVx1_ASAP7_75t_L g1346 ( .A(n_285), .Y(n_1346) );
OAI211xp5_ASAP7_75t_SL g1353 ( .A1(n_285), .A2(n_649), .B(n_1354), .C(n_1355), .Y(n_1353) );
OAI22xp33_ASAP7_75t_L g1193 ( .A1(n_286), .A2(n_287), .B1(n_362), .B2(n_641), .Y(n_1193) );
OAI22xp33_ASAP7_75t_L g1201 ( .A1(n_286), .A2(n_287), .B1(n_659), .B2(n_1202), .Y(n_1201) );
INVx1_ASAP7_75t_L g548 ( .A(n_289), .Y(n_548) );
INVx1_ASAP7_75t_L g1417 ( .A(n_290), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_290), .B(n_1416), .Y(n_1422) );
INVx1_ASAP7_75t_L g1253 ( .A(n_292), .Y(n_1253) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_293), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_294), .A2(n_331), .B1(n_477), .B2(n_483), .Y(n_1352) );
CKINVDCx5p33_ASAP7_75t_R g1206 ( .A(n_295), .Y(n_1206) );
INVx1_ASAP7_75t_L g1262 ( .A(n_296), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_297), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_298), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g1759 ( .A1(n_299), .A2(n_573), .B(n_598), .C(n_1760), .Y(n_1759) );
OAI211xp5_ASAP7_75t_SL g1767 ( .A1(n_299), .A2(n_649), .B(n_1768), .C(n_1769), .Y(n_1767) );
INVx1_ASAP7_75t_L g1071 ( .A(n_300), .Y(n_1071) );
OAI21xp33_ASAP7_75t_L g1673 ( .A1(n_301), .A2(n_1674), .B(n_1678), .Y(n_1673) );
INVx1_ASAP7_75t_L g1392 ( .A(n_302), .Y(n_1392) );
OAI211xp5_ASAP7_75t_SL g1397 ( .A1(n_302), .A2(n_649), .B(n_1398), .C(n_1400), .Y(n_1397) );
INVx1_ASAP7_75t_L g590 ( .A(n_303), .Y(n_590) );
XOR2x2_ASAP7_75t_L g1050 ( .A(n_304), .B(n_1051), .Y(n_1050) );
OAI211xp5_ASAP7_75t_L g1187 ( .A1(n_306), .A2(n_628), .B(n_1170), .C(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1200 ( .A(n_306), .Y(n_1200) );
OAI211xp5_ASAP7_75t_L g969 ( .A1(n_308), .A2(n_628), .B(n_970), .C(n_971), .Y(n_969) );
INVx1_ASAP7_75t_L g983 ( .A(n_308), .Y(n_983) );
INVxp67_ASAP7_75t_SL g1022 ( .A(n_310), .Y(n_1022) );
AOI22xp33_ASAP7_75t_SL g1291 ( .A1(n_311), .A2(n_341), .B1(n_1292), .B2(n_1295), .Y(n_1291) );
INVx1_ASAP7_75t_L g1173 ( .A(n_312), .Y(n_1173) );
OAI211xp5_ASAP7_75t_L g1180 ( .A1(n_312), .A2(n_831), .B(n_960), .C(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1002 ( .A(n_313), .Y(n_1002) );
OAI211xp5_ASAP7_75t_SL g624 ( .A1(n_314), .A2(n_625), .B(n_628), .C(n_630), .Y(n_624) );
INVx1_ASAP7_75t_L g653 ( .A(n_314), .Y(n_653) );
INVx1_ASAP7_75t_L g667 ( .A(n_315), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g1337 ( .A(n_316), .Y(n_1337) );
CKINVDCx5p33_ASAP7_75t_R g1207 ( .A(n_317), .Y(n_1207) );
INVx1_ASAP7_75t_L g881 ( .A(n_318), .Y(n_881) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_319), .Y(n_366) );
INVx1_ASAP7_75t_L g1155 ( .A(n_320), .Y(n_1155) );
CKINVDCx5p33_ASAP7_75t_R g1210 ( .A(n_321), .Y(n_1210) );
INVx1_ASAP7_75t_L g724 ( .A(n_323), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_324), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g1347 ( .A(n_328), .Y(n_1347) );
CKINVDCx5p33_ASAP7_75t_R g1744 ( .A(n_329), .Y(n_1744) );
XOR2x2_ASAP7_75t_L g1184 ( .A(n_330), .B(n_1185), .Y(n_1184) );
INVx2_ASAP7_75t_L g454 ( .A(n_332), .Y(n_454) );
INVx1_ASAP7_75t_L g506 ( .A(n_332), .Y(n_506) );
INVx1_ASAP7_75t_L g528 ( .A(n_332), .Y(n_528) );
INVx1_ASAP7_75t_L g757 ( .A(n_333), .Y(n_757) );
INVx1_ASAP7_75t_L g941 ( .A(n_334), .Y(n_941) );
INVx1_ASAP7_75t_L g1367 ( .A(n_336), .Y(n_1367) );
INVx1_ASAP7_75t_L g919 ( .A(n_337), .Y(n_919) );
INVx1_ASAP7_75t_L g1370 ( .A(n_338), .Y(n_1370) );
AOI21xp33_ASAP7_75t_L g439 ( .A1(n_339), .A2(n_440), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g512 ( .A(n_339), .Y(n_512) );
INVx1_ASAP7_75t_L g910 ( .A(n_340), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_342), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_343), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_371), .B(n_1404), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx4f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_356), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g1727 ( .A(n_350), .B(n_359), .Y(n_1727) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g1731 ( .A(n_352), .B(n_355), .Y(n_1731) );
INVx1_ASAP7_75t_L g1773 ( .A(n_352), .Y(n_1773) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g1775 ( .A(n_355), .B(n_1773), .Y(n_1775) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AOI21xp5_ASAP7_75t_SL g380 ( .A1(n_359), .A2(n_381), .B(n_415), .Y(n_380) );
AND2x4_ASAP7_75t_L g616 ( .A(n_359), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g435 ( .A(n_360), .B(n_370), .Y(n_435) );
AND2x4_ASAP7_75t_L g443 ( .A(n_360), .B(n_369), .Y(n_443) );
AND2x4_ASAP7_75t_SL g1726 ( .A(n_361), .B(n_1727), .Y(n_1726) );
INVx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_363), .B(n_368), .Y(n_362) );
BUFx4f_ASAP7_75t_L g418 ( .A(n_363), .Y(n_418) );
OR2x6_ASAP7_75t_L g637 ( .A(n_363), .B(n_384), .Y(n_637) );
OR2x2_ASAP7_75t_L g865 ( .A(n_363), .B(n_384), .Y(n_865) );
INVx1_ASAP7_75t_L g1271 ( .A(n_363), .Y(n_1271) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g403 ( .A(n_364), .Y(n_403) );
BUFx4f_ASAP7_75t_L g689 ( .A(n_364), .Y(n_689) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x2_ASAP7_75t_L g386 ( .A(n_366), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g393 ( .A(n_366), .B(n_367), .Y(n_393) );
INVx1_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
INVx2_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
NAND2x1_ASAP7_75t_L g427 ( .A(n_366), .B(n_367), .Y(n_427) );
INVx2_ASAP7_75t_L g433 ( .A(n_366), .Y(n_433) );
INVx2_ASAP7_75t_L g387 ( .A(n_367), .Y(n_387) );
BUFx2_ASAP7_75t_L g398 ( .A(n_367), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_367), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g432 ( .A(n_367), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g448 ( .A(n_367), .Y(n_448) );
AND2x2_ASAP7_75t_L g450 ( .A(n_367), .B(n_413), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_368), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_399) );
OR2x6_ASAP7_75t_L g614 ( .A(n_368), .B(n_403), .Y(n_614) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g397 ( .A(n_369), .Y(n_397) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g389 ( .A(n_370), .Y(n_389) );
AND2x4_ASAP7_75t_L g405 ( .A(n_370), .B(n_406), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_1226), .B2(n_1227), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
XNOR2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_775), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_619), .B2(n_774), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
XOR2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_539), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_451), .B(n_455), .Y(n_379) );
INVx3_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx4_ASAP7_75t_L g615 ( .A(n_383), .Y(n_615) );
CKINVDCx16_ASAP7_75t_R g641 ( .A(n_383), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g1019 ( .A1(n_383), .A2(n_1020), .B1(n_1021), .B2(n_1022), .Y(n_1019) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_386), .Y(n_441) );
BUFx3_ASAP7_75t_L g1279 ( .A(n_386), .Y(n_1279) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B(n_391), .C(n_394), .Y(n_388) );
INVx1_ASAP7_75t_L g401 ( .A(n_389), .Y(n_401) );
OR2x2_ASAP7_75t_L g410 ( .A(n_389), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g603 ( .A(n_389), .B(n_398), .Y(n_603) );
AND2x2_ASAP7_75t_L g608 ( .A(n_389), .B(n_609), .Y(n_608) );
AND2x4_ASAP7_75t_L g632 ( .A(n_389), .B(n_398), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g602 ( .A1(n_391), .A2(n_590), .B1(n_591), .B2(n_603), .C1(n_604), .C2(n_605), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g1306 ( .A1(n_391), .A2(n_605), .B1(n_632), .B2(n_1307), .C1(n_1308), .C2(n_1309), .Y(n_1306) );
BUFx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g629 ( .A(n_392), .B(n_397), .Y(n_629) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_392), .Y(n_1040) );
AND2x6_ASAP7_75t_L g1702 ( .A(n_392), .B(n_1639), .Y(n_1702) );
AND2x4_ASAP7_75t_SL g1710 ( .A(n_392), .B(n_1691), .Y(n_1710) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g601 ( .A(n_393), .Y(n_601) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_396), .A2(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_396), .A2(n_605), .B1(n_861), .B2(n_862), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_396), .A2(n_405), .B1(n_1010), .B2(n_1014), .Y(n_1026) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g599 ( .A(n_397), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g612 ( .A(n_397), .B(n_411), .Y(n_612) );
INVx1_ASAP7_75t_L g1721 ( .A(n_398), .Y(n_1721) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_400), .A2(n_490), .B1(n_492), .B2(n_493), .Y(n_489) );
BUFx3_ASAP7_75t_L g569 ( .A(n_403), .Y(n_569) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_403), .Y(n_579) );
BUFx3_ASAP7_75t_L g666 ( .A(n_403), .Y(n_666) );
INVx2_ASAP7_75t_L g822 ( .A(n_404), .Y(n_822) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g605 ( .A(n_405), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_405), .A2(n_632), .B1(n_757), .B2(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g930 ( .A(n_405), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_406), .B(n_1639), .Y(n_1676) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_409), .B(n_414), .Y(n_408) );
INVx2_ASAP7_75t_L g1349 ( .A(n_409), .Y(n_1349) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_L g639 ( .A(n_410), .Y(n_639) );
INVx2_ASAP7_75t_L g772 ( .A(n_410), .Y(n_772) );
INVx8_ASAP7_75t_L g422 ( .A(n_411), .Y(n_422) );
BUFx2_ASAP7_75t_L g899 ( .A(n_411), .Y(n_899) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_423), .B(n_436), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g898 ( .A1(n_418), .A2(n_881), .B1(n_892), .B2(n_899), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_418), .A2(n_841), .B1(n_886), .B2(n_890), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g1164 ( .A1(n_418), .A2(n_420), .B1(n_1145), .B2(n_1161), .Y(n_1164) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_419), .A2(n_437), .B1(n_531), .B2(n_533), .C(n_536), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g1167 ( .A1(n_420), .A2(n_740), .B1(n_1151), .B2(n_1156), .Y(n_1167) );
OAI22xp5_ASAP7_75t_L g1714 ( .A1(n_420), .A2(n_1715), .B1(n_1716), .B2(n_1717), .Y(n_1714) );
INVx5_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx6_ASAP7_75t_L g668 ( .A(n_421), .Y(n_668) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx4_ASAP7_75t_L g570 ( .A(n_422), .Y(n_570) );
INVx2_ASAP7_75t_L g581 ( .A(n_422), .Y(n_581) );
INVx1_ASAP7_75t_L g692 ( .A(n_422), .Y(n_692) );
INVx1_ASAP7_75t_L g741 ( .A(n_422), .Y(n_741) );
INVx2_ASAP7_75t_SL g841 ( .A(n_422), .Y(n_841) );
INVx2_ASAP7_75t_L g953 ( .A(n_422), .Y(n_953) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_428), .B1(n_429), .B2(n_434), .C(n_435), .Y(n_423) );
OAI22xp5_ASAP7_75t_SL g900 ( .A1(n_424), .A2(n_814), .B1(n_885), .B2(n_889), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_424), .A2(n_429), .B1(n_882), .B2(n_893), .Y(n_901) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g812 ( .A(n_425), .Y(n_812) );
INVx1_ASAP7_75t_L g819 ( .A(n_425), .Y(n_819) );
INVx2_ASAP7_75t_L g970 ( .A(n_425), .Y(n_970) );
INVx4_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx4f_ASAP7_75t_L g438 ( .A(n_426), .Y(n_438) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_426), .Y(n_573) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_426), .Y(n_577) );
BUFx4f_ASAP7_75t_L g627 ( .A(n_426), .Y(n_627) );
BUFx4f_ASAP7_75t_L g744 ( .A(n_426), .Y(n_744) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g675 ( .A(n_427), .Y(n_675) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g671 ( .A(n_431), .Y(n_671) );
INVx2_ASAP7_75t_L g811 ( .A(n_431), .Y(n_811) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx3_ASAP7_75t_L g572 ( .A(n_432), .Y(n_572) );
INVx1_ASAP7_75t_L g576 ( .A(n_432), .Y(n_576) );
BUFx2_ASAP7_75t_L g679 ( .A(n_432), .Y(n_679) );
BUFx2_ASAP7_75t_L g814 ( .A(n_432), .Y(n_814) );
AND2x2_ASAP7_75t_L g447 ( .A(n_433), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_SL g583 ( .A(n_435), .B(n_504), .Y(n_583) );
AND2x4_ASAP7_75t_L g683 ( .A(n_435), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g1698 ( .A(n_435), .Y(n_1698) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_438), .B(n_439), .C(n_444), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_438), .A2(n_743), .B1(n_1147), .B2(n_1162), .Y(n_1166) );
BUFx3_ASAP7_75t_L g1697 ( .A(n_440), .Y(n_1697) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g1692 ( .A(n_441), .B(n_1691), .Y(n_1692) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g1711 ( .A1(n_443), .A2(n_573), .B1(n_946), .B2(n_1712), .C(n_1713), .Y(n_1711) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g1038 ( .A(n_446), .Y(n_1038) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_447), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g1638 ( .A(n_447), .B(n_1639), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_447), .B(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_SL g1701 ( .A(n_449), .Y(n_1701) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g1046 ( .A(n_450), .Y(n_1046) );
BUFx6f_ASAP7_75t_L g1705 ( .A(n_450), .Y(n_1705) );
INVx2_ASAP7_75t_L g1723 ( .A(n_451), .Y(n_1723) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR2x6_ASAP7_75t_L g562 ( .A(n_453), .B(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g566 ( .A(n_453), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g806 ( .A(n_453), .B(n_563), .Y(n_806) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g997 ( .A(n_454), .Y(n_997) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_498), .B(n_507), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_457), .B(n_489), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_476), .C(n_486), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g543 ( .A1(n_459), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_543) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g648 ( .A(n_460), .Y(n_648) );
INVx1_ASAP7_75t_L g734 ( .A(n_460), .Y(n_734) );
INVx1_ASAP7_75t_L g960 ( .A(n_460), .Y(n_960) );
INVx1_ASAP7_75t_L g980 ( .A(n_460), .Y(n_980) );
INVx4_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_461), .Y(n_560) );
INVx3_ASAP7_75t_L g790 ( .A(n_461), .Y(n_790) );
HB1xp67_ASAP7_75t_L g1382 ( .A(n_461), .Y(n_1382) );
OR2x2_ASAP7_75t_L g1677 ( .A(n_461), .B(n_1634), .Y(n_1677) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g699 ( .A(n_462), .Y(n_699) );
BUFx2_ASAP7_75t_L g754 ( .A(n_462), .Y(n_754) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .Y(n_462) );
BUFx2_ASAP7_75t_L g475 ( .A(n_463), .Y(n_475) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_464), .B(n_466), .Y(n_485) );
INVx2_ASAP7_75t_L g488 ( .A(n_464), .Y(n_488) );
BUFx2_ASAP7_75t_L g472 ( .A(n_465), .Y(n_472) );
AND2x4_ASAP7_75t_L g522 ( .A(n_465), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g1359 ( .A(n_465), .Y(n_1359) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g480 ( .A(n_466), .B(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g487 ( .A(n_466), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g497 ( .A(n_466), .Y(n_497) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_468), .A2(n_474), .B1(n_588), .B2(n_589), .C1(n_590), .C2(n_591), .Y(n_587) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_468), .A2(n_474), .B1(n_821), .B2(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_468), .A2(n_474), .B1(n_861), .B2(n_870), .Y(n_869) );
AOI222xp33_ASAP7_75t_L g907 ( .A1(n_468), .A2(n_655), .B1(n_908), .B2(n_909), .C1(n_910), .C2(n_911), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_468), .A2(n_474), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_468), .A2(n_474), .B1(n_1056), .B2(n_1065), .Y(n_1064) );
AOI22xp5_ASAP7_75t_L g1769 ( .A1(n_468), .A2(n_1356), .B1(n_1761), .B2(n_1770), .Y(n_1769) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_472), .Y(n_468) );
AND2x2_ASAP7_75t_L g474 ( .A(n_469), .B(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g652 ( .A(n_469), .B(n_472), .Y(n_652) );
AND2x4_ASAP7_75t_L g655 ( .A(n_469), .B(n_475), .Y(n_655) );
AND2x4_ASAP7_75t_L g982 ( .A(n_469), .B(n_472), .Y(n_982) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND3x4_ASAP7_75t_L g996 ( .A(n_470), .B(n_501), .C(n_997), .Y(n_996) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_470), .B(n_1357), .Y(n_1356) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g479 ( .A(n_471), .Y(n_479) );
NAND2xp33_ASAP7_75t_SL g510 ( .A(n_471), .B(n_501), .Y(n_510) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_474), .A2(n_982), .B1(n_1236), .B2(n_1245), .Y(n_1244) );
AOI32xp33_ASAP7_75t_L g1355 ( .A1(n_474), .A2(n_1347), .A3(n_1356), .B1(n_1358), .B2(n_1360), .Y(n_1355) );
INVxp67_ASAP7_75t_L g1768 ( .A(n_474), .Y(n_1768) );
BUFx2_ASAP7_75t_L g645 ( .A(n_477), .Y(n_645) );
BUFx3_ASAP7_75t_L g760 ( .A(n_477), .Y(n_760) );
INVx2_ASAP7_75t_SL g920 ( .A(n_477), .Y(n_920) );
OR2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
AND2x2_ASAP7_75t_L g493 ( .A(n_478), .B(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g660 ( .A(n_478), .B(n_494), .Y(n_660) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR2x6_ASAP7_75t_L g483 ( .A(n_479), .B(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_L g486 ( .A(n_479), .B(n_487), .Y(n_486) );
OR2x4_ASAP7_75t_L g491 ( .A(n_479), .B(n_480), .Y(n_491) );
NAND3x1_ASAP7_75t_L g526 ( .A(n_479), .B(n_527), .C(n_529), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_479), .B(n_529), .Y(n_563) );
AND2x4_ASAP7_75t_L g1646 ( .A(n_479), .B(n_1647), .Y(n_1646) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_480), .Y(n_544) );
BUFx3_ASAP7_75t_L g697 ( .A(n_480), .Y(n_697) );
BUFx3_ASAP7_75t_L g709 ( .A(n_480), .Y(n_709) );
INVx2_ASAP7_75t_L g803 ( .A(n_480), .Y(n_803) );
INVx1_ASAP7_75t_L g518 ( .A(n_481), .Y(n_518) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVxp67_ASAP7_75t_L g496 ( .A(n_482), .Y(n_496) );
INVx2_ASAP7_75t_L g594 ( .A(n_483), .Y(n_594) );
INVx1_ASAP7_75t_L g762 ( .A(n_483), .Y(n_762) );
INVx1_ASAP7_75t_L g915 ( .A(n_483), .Y(n_915) );
BUFx3_ASAP7_75t_L g985 ( .A(n_483), .Y(n_985) );
BUFx3_ASAP7_75t_L g703 ( .A(n_484), .Y(n_703) );
INVx1_ASAP7_75t_L g727 ( .A(n_484), .Y(n_727) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g535 ( .A(n_485), .Y(n_535) );
CKINVDCx8_ASAP7_75t_R g649 ( .A(n_486), .Y(n_649) );
CKINVDCx8_ASAP7_75t_R g831 ( .A(n_486), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_486), .B(n_906), .Y(n_905) );
BUFx2_ASAP7_75t_L g519 ( .A(n_487), .Y(n_519) );
BUFx2_ASAP7_75t_L g588 ( .A(n_487), .Y(n_588) );
BUFx2_ASAP7_75t_L g911 ( .A(n_487), .Y(n_911) );
BUFx3_ASAP7_75t_L g1001 ( .A(n_487), .Y(n_1001) );
INVx2_ASAP7_75t_L g1012 ( .A(n_487), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1063 ( .A(n_487), .Y(n_1063) );
BUFx2_ASAP7_75t_L g1672 ( .A(n_487), .Y(n_1672) );
INVx1_ASAP7_75t_L g523 ( .A(n_488), .Y(n_523) );
INVx1_ASAP7_75t_L g1202 ( .A(n_490), .Y(n_1202) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_SL g658 ( .A(n_491), .Y(n_658) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_491), .Y(n_749) );
INVx1_ASAP7_75t_L g918 ( .A(n_491), .Y(n_918) );
INVx2_ASAP7_75t_SL g1314 ( .A(n_491), .Y(n_1314) );
INVx2_ASAP7_75t_L g586 ( .A(n_493), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_493), .A2(n_913), .B1(n_914), .B2(n_915), .Y(n_912) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_494), .Y(n_514) );
BUFx6f_ASAP7_75t_L g702 ( .A(n_494), .Y(n_702) );
INVx2_ASAP7_75t_L g705 ( .A(n_494), .Y(n_705) );
INVx1_ASAP7_75t_L g730 ( .A(n_494), .Y(n_730) );
INVx2_ASAP7_75t_L g964 ( .A(n_494), .Y(n_964) );
INVx2_ASAP7_75t_L g1386 ( .A(n_494), .Y(n_1386) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g532 ( .A(n_495), .Y(n_532) );
BUFx8_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_495), .Y(n_723) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
AND2x4_ASAP7_75t_L g517 ( .A(n_497), .B(n_518), .Y(n_517) );
OAI31xp33_ASAP7_75t_L g643 ( .A1(n_498), .A2(n_644), .A3(n_647), .B(n_656), .Y(n_643) );
BUFx2_ASAP7_75t_L g1137 ( .A(n_498), .Y(n_1137) );
AND2x2_ASAP7_75t_SL g498 ( .A(n_499), .B(n_502), .Y(n_498) );
AND2x2_ASAP7_75t_L g595 ( .A(n_499), .B(n_502), .Y(n_595) );
AND2x2_ASAP7_75t_L g763 ( .A(n_499), .B(n_502), .Y(n_763) );
AND2x4_ASAP7_75t_L g922 ( .A(n_499), .B(n_502), .Y(n_922) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_499), .B(n_502), .Y(n_1017) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g1647 ( .A(n_501), .Y(n_1647) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g509 ( .A(n_504), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g685 ( .A(n_504), .Y(n_685) );
OR2x2_ASAP7_75t_L g1634 ( .A(n_504), .B(n_1635), .Y(n_1634) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g618 ( .A(n_505), .Y(n_618) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_511), .B1(n_524), .B2(n_530), .Y(n_507) );
OAI33xp33_ASAP7_75t_L g542 ( .A1(n_508), .A2(n_543), .A3(n_547), .B1(n_552), .B2(n_558), .B3(n_562), .Y(n_542) );
OAI33xp33_ASAP7_75t_L g878 ( .A1(n_508), .A2(n_562), .A3(n_879), .B1(n_883), .B2(n_887), .B3(n_891), .Y(n_878) );
OAI33xp33_ASAP7_75t_L g1380 ( .A1(n_508), .A2(n_524), .A3(n_1381), .B1(n_1383), .B2(n_1385), .B3(n_1387), .Y(n_1380) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx8_ASAP7_75t_L g695 ( .A(n_509), .Y(n_695) );
BUFx4f_ASAP7_75t_L g785 ( .A(n_509), .Y(n_785) );
BUFx4f_ASAP7_75t_L g1111 ( .A(n_509), .Y(n_1111) );
OAI211xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_515), .C(n_520), .Y(n_511) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_SL g1003 ( .A(n_516), .Y(n_1003) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx8_ASAP7_75t_L g538 ( .A(n_517), .Y(n_538) );
BUFx3_ASAP7_75t_L g1294 ( .A(n_517), .Y(n_1294) );
NAND2x1p5_ASAP7_75t_L g1657 ( .A(n_517), .B(n_1646), .Y(n_1657) );
AND2x4_ASAP7_75t_L g1660 ( .A(n_519), .B(n_1645), .Y(n_1660) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx5_ASAP7_75t_L g994 ( .A(n_522), .Y(n_994) );
BUFx3_ASAP7_75t_L g1290 ( .A(n_522), .Y(n_1290) );
BUFx12f_ASAP7_75t_L g1298 ( .A(n_522), .Y(n_1298) );
INVx1_ASAP7_75t_L g1357 ( .A(n_523), .Y(n_1357) );
OAI33xp33_ASAP7_75t_L g694 ( .A1(n_524), .A2(n_695), .A3(n_696), .B1(n_700), .B2(n_704), .B3(n_706), .Y(n_694) );
OAI33xp33_ASAP7_75t_L g714 ( .A1(n_524), .A2(n_695), .A3(n_715), .B1(n_719), .B2(n_728), .B3(n_732), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g965 ( .A(n_525), .Y(n_965) );
INVx2_ASAP7_75t_L g1119 ( .A(n_525), .Y(n_1119) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx3_ASAP7_75t_L g1159 ( .A(n_526), .Y(n_1159) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g1637 ( .A(n_528), .Y(n_1637) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_531), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_547) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx3_ASAP7_75t_L g798 ( .A(n_532), .Y(n_798) );
BUFx2_ASAP7_75t_L g884 ( .A(n_532), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_533), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
OAI22xp33_ASAP7_75t_SL g963 ( .A1(n_533), .A2(n_947), .B1(n_954), .B2(n_964), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_533), .A2(n_722), .B1(n_1101), .B2(n_1108), .Y(n_1117) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_533), .A2(n_1153), .B1(n_1155), .B2(n_1156), .Y(n_1152) );
CKINVDCx8_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g556 ( .A(n_534), .Y(n_556) );
INVx3_ASAP7_75t_L g794 ( .A(n_534), .Y(n_794) );
INVx3_ASAP7_75t_L g1086 ( .A(n_534), .Y(n_1086) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g551 ( .A(n_535), .Y(n_551) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g1669 ( .A(n_538), .Y(n_1669) );
INVx2_ASAP7_75t_L g1681 ( .A(n_538), .Y(n_1681) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_584), .C(n_596), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_564), .Y(n_541) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_544), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_544), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g1087 ( .A1(n_544), .A2(n_734), .B1(n_1071), .B2(n_1077), .Y(n_1087) );
OAI22xp33_ASAP7_75t_L g1251 ( .A1(n_544), .A2(n_560), .B1(n_1252), .B2(n_1253), .Y(n_1251) );
OAI22xp33_ASAP7_75t_L g1261 ( .A1(n_544), .A2(n_699), .B1(n_1262), .B2(n_1263), .Y(n_1261) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_544), .A2(n_560), .B1(n_1327), .B2(n_1328), .Y(n_1326) );
OAI22xp33_ASAP7_75t_L g1335 ( .A1(n_544), .A2(n_699), .B1(n_1336), .B2(n_1337), .Y(n_1335) );
OAI22xp5_ASAP7_75t_L g1740 ( .A1(n_544), .A2(n_789), .B1(n_1741), .B2(n_1742), .Y(n_1740) );
OAI22xp5_ASAP7_75t_L g1749 ( .A1(n_544), .A2(n_699), .B1(n_1750), .B2(n_1751), .Y(n_1749) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_545), .A2(n_559), .B1(n_569), .B2(n_570), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_546), .A2(n_561), .B1(n_575), .B2(n_577), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_548), .A2(n_555), .B1(n_572), .B2(n_573), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_549), .A2(n_557), .B1(n_579), .B2(n_580), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_550), .A2(n_884), .B1(n_885), .B2(n_886), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_550), .A2(n_888), .B1(n_889), .B2(n_890), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_550), .A2(n_1258), .B1(n_1259), .B2(n_1260), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_550), .A2(n_1084), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g1633 ( .A(n_551), .B(n_1634), .Y(n_1633) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_555), .B1(n_556), .B2(n_557), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g1254 ( .A1(n_553), .A2(n_800), .B1(n_1255), .B2(n_1256), .Y(n_1254) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g888 ( .A(n_554), .Y(n_888) );
INVx2_ASAP7_75t_SL g1258 ( .A(n_554), .Y(n_1258) );
AND2x4_ASAP7_75t_L g1684 ( .A(n_554), .B(n_1682), .Y(n_1684) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_556), .A2(n_845), .B1(n_851), .B2(n_856), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_560), .A2(n_802), .B1(n_840), .B2(n_847), .Y(n_853) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_560), .A2(n_697), .B1(n_892), .B2(n_893), .Y(n_891) );
INVx1_ASAP7_75t_L g1198 ( .A(n_560), .Y(n_1198) );
INVx1_ASAP7_75t_L g1005 ( .A(n_562), .Y(n_1005) );
OAI33xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .A3(n_571), .B1(n_574), .B2(n_578), .B3(n_582), .Y(n_564) );
OAI33xp33_ASAP7_75t_L g807 ( .A1(n_565), .A2(n_808), .A3(n_810), .B1(n_813), .B2(n_815), .B3(n_816), .Y(n_807) );
OAI33xp33_ASAP7_75t_L g1264 ( .A1(n_565), .A2(n_582), .A3(n_1265), .B1(n_1266), .B2(n_1268), .B3(n_1269), .Y(n_1264) );
OAI33xp33_ASAP7_75t_L g1338 ( .A1(n_565), .A2(n_582), .A3(n_1339), .B1(n_1340), .B2(n_1341), .B3(n_1342), .Y(n_1338) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx4_ASAP7_75t_L g663 ( .A(n_566), .Y(n_663) );
INVx2_ASAP7_75t_L g738 ( .A(n_566), .Y(n_738) );
INVx2_ASAP7_75t_L g1095 ( .A(n_566), .Y(n_1095) );
INVx1_ASAP7_75t_L g1208 ( .A(n_566), .Y(n_1208) );
OAI22xp5_ASAP7_75t_L g1753 ( .A1(n_569), .A2(n_580), .B1(n_1741), .B2(n_1750), .Y(n_1753) );
OAI22xp5_ASAP7_75t_L g1756 ( .A1(n_569), .A2(n_570), .B1(n_1745), .B2(n_1748), .Y(n_1756) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_570), .A2(n_793), .B1(n_799), .B2(n_809), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_570), .A2(n_1256), .B1(n_1260), .B2(n_1270), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_570), .A2(n_809), .B1(n_1327), .B2(n_1336), .Y(n_1339) );
OAI22xp5_ASAP7_75t_L g1342 ( .A1(n_570), .A2(n_1270), .B1(n_1331), .B2(n_1334), .Y(n_1342) );
OAI22xp5_ASAP7_75t_L g1755 ( .A1(n_572), .A2(n_970), .B1(n_1742), .B2(n_1751), .Y(n_1755) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_575), .A2(n_673), .B1(n_949), .B2(n_950), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g1209 ( .A1(n_575), .A2(n_819), .B1(n_1210), .B2(n_1211), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_575), .A2(n_627), .B1(n_1213), .B2(n_1214), .Y(n_1212) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g1267 ( .A(n_576), .Y(n_1267) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_577), .A2(n_811), .B1(n_847), .B2(n_848), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_577), .A2(n_811), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_577), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_580), .A2(n_787), .B1(n_804), .B2(n_809), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_580), .A2(n_809), .B1(n_850), .B2(n_851), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g1069 ( .A1(n_580), .A2(n_809), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI33xp33_ASAP7_75t_L g1752 ( .A1(n_582), .A2(n_738), .A3(n_1753), .B1(n_1754), .B2(n_1755), .B3(n_1756), .Y(n_1752) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g816 ( .A(n_583), .Y(n_816) );
AOI33xp33_ASAP7_75t_L g1036 ( .A1(n_583), .A2(n_897), .A3(n_1037), .B1(n_1039), .B2(n_1041), .B3(n_1042), .Y(n_1036) );
NAND3xp33_ASAP7_75t_L g1283 ( .A(n_583), .B(n_1284), .C(n_1286), .Y(n_1283) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_592), .B(n_595), .Y(n_584) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g646 ( .A(n_594), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_594), .A2(n_920), .B1(n_1304), .B2(n_1305), .Y(n_1317) );
OAI31xp33_ASAP7_75t_SL g826 ( .A1(n_595), .A2(n_827), .A3(n_828), .B(n_834), .Y(n_826) );
OAI31xp33_ASAP7_75t_SL g866 ( .A1(n_595), .A2(n_867), .A3(n_868), .B(n_871), .Y(n_866) );
OAI31xp33_ASAP7_75t_L g1240 ( .A1(n_595), .A2(n_1241), .A3(n_1243), .B(n_1248), .Y(n_1240) );
OAI21xp5_ASAP7_75t_L g1311 ( .A1(n_595), .A2(n_1312), .B(n_1315), .Y(n_1311) );
OAI31xp33_ASAP7_75t_SL g1351 ( .A1(n_595), .A2(n_1352), .A3(n_1353), .B(n_1361), .Y(n_1351) );
OAI31xp33_ASAP7_75t_SL g1764 ( .A1(n_595), .A2(n_1765), .A3(n_1766), .B(n_1767), .Y(n_1764) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_613), .B(n_616), .Y(n_596) );
NAND3xp33_ASAP7_75t_SL g597 ( .A(n_598), .B(n_602), .C(n_606), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g1302 ( .A(n_598), .B(n_1303), .C(n_1306), .Y(n_1302) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g1030 ( .A(n_599), .Y(n_1030) );
INVx1_ASAP7_75t_L g1029 ( .A(n_600), .Y(n_1029) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx2_ASAP7_75t_L g1696 ( .A(n_601), .Y(n_1696) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_603), .A2(n_1189), .B1(n_1190), .B2(n_1191), .Y(n_1188) );
AOI22xp5_ASAP7_75t_L g1345 ( .A1(n_603), .A2(n_822), .B1(n_1346), .B2(n_1347), .Y(n_1345) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_605), .A2(n_631), .B1(n_633), .B2(n_634), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_605), .A2(n_632), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_605), .A2(n_632), .B1(n_1236), .B2(n_1237), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_605), .A2(n_631), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
AOI22xp5_ASAP7_75t_L g1760 ( .A1(n_605), .A2(n_632), .B1(n_1761), .B2(n_1762), .Y(n_1760) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_610), .B2(n_611), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_608), .A2(n_772), .B1(n_1304), .B2(n_1305), .Y(n_1303) );
INVx3_ASAP7_75t_L g1044 ( .A(n_609), .Y(n_1044) );
BUFx6f_ASAP7_75t_L g1285 ( .A(n_609), .Y(n_1285) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g1021 ( .A(n_614), .Y(n_1021) );
BUFx2_ASAP7_75t_L g642 ( .A(n_616), .Y(n_642) );
BUFx2_ASAP7_75t_SL g773 ( .A(n_616), .Y(n_773) );
INVx1_ASAP7_75t_L g1031 ( .A(n_616), .Y(n_1031) );
OAI31xp33_ASAP7_75t_L g1052 ( .A1(n_616), .A2(n_1053), .A3(n_1054), .B(n_1058), .Y(n_1052) );
BUFx3_ASAP7_75t_L g1129 ( .A(n_616), .Y(n_1129) );
OAI31xp33_ASAP7_75t_L g1757 ( .A1(n_616), .A2(n_1758), .A3(n_1759), .B(n_1763), .Y(n_1757) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_L g1658 ( .A(n_618), .Y(n_1658) );
OR2x2_ASAP7_75t_L g1675 ( .A(n_618), .B(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g774 ( .A(n_619), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_710), .B2(n_711), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_643), .C(n_661), .Y(n_622) );
OAI31xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_635), .A3(n_640), .B(n_642), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_627), .A2(n_945), .B1(n_946), .B2(n_947), .Y(n_944) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g767 ( .A(n_629), .Y(n_767) );
INVx1_ASAP7_75t_L g1127 ( .A(n_629), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_631), .A2(n_929), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
BUFx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_632), .A2(n_908), .B1(n_910), .B2(n_929), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_632), .A2(n_822), .B1(n_972), .B2(n_973), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_632), .A2(n_822), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_633), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_650) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g1175 ( .A(n_637), .Y(n_1175) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI31xp33_ASAP7_75t_L g817 ( .A1(n_642), .A2(n_818), .A3(n_824), .B(n_825), .Y(n_817) );
OAI31xp33_ASAP7_75t_L g858 ( .A1(n_642), .A2(n_859), .A3(n_863), .B(n_864), .Y(n_858) );
INVx1_ASAP7_75t_L g933 ( .A(n_642), .Y(n_933) );
OAI31xp33_ASAP7_75t_L g968 ( .A1(n_642), .A2(n_969), .A3(n_974), .B(n_976), .Y(n_968) );
OAI31xp33_ASAP7_75t_L g1343 ( .A1(n_642), .A2(n_1344), .A3(n_1348), .B(n_1350), .Y(n_1343) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_648), .A2(n_667), .B1(n_681), .B2(n_707), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g1160 ( .A1(n_648), .A2(n_1146), .B1(n_1161), .B2(n_1162), .Y(n_1160) );
OAI22xp33_ASAP7_75t_L g1223 ( .A1(n_648), .A2(n_707), .B1(n_1207), .B2(n_1214), .Y(n_1223) );
NAND3xp33_ASAP7_75t_L g1315 ( .A(n_649), .B(n_1316), .C(n_1317), .Y(n_1315) );
AOI222xp33_ASAP7_75t_L g1316 ( .A1(n_651), .A2(n_655), .B1(n_911), .B2(n_1307), .C1(n_1308), .C2(n_1309), .Y(n_1316) );
BUFx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
BUFx3_ASAP7_75t_L g756 ( .A(n_652), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_654), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_654), .A2(n_756), .B1(n_1125), .B2(n_1134), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_654), .A2(n_756), .B1(n_1391), .B2(n_1401), .Y(n_1400) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_655), .A2(n_972), .B1(n_982), .B2(n_983), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g1181 ( .A1(n_655), .A2(n_982), .B1(n_1172), .B2(n_1182), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_655), .A2(n_982), .B1(n_1189), .B2(n_1200), .Y(n_1199) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g750 ( .A(n_660), .Y(n_750) );
INVx1_ASAP7_75t_L g1242 ( .A(n_660), .Y(n_1242) );
NOR2xp33_ASAP7_75t_SL g661 ( .A(n_662), .B(n_694), .Y(n_661) );
OAI33xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .A3(n_669), .B1(n_676), .B2(n_682), .B3(n_686), .Y(n_662) );
INVx2_ASAP7_75t_SL g897 ( .A(n_663), .Y(n_897) );
OAI33xp33_ASAP7_75t_L g939 ( .A1(n_663), .A2(n_940), .A3(n_944), .B1(n_948), .B2(n_951), .B3(n_955), .Y(n_939) );
INVx2_ASAP7_75t_SL g1282 ( .A(n_663), .Y(n_1282) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g696 ( .A1(n_665), .A2(n_680), .B1(n_697), .B2(n_698), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_666), .A2(n_668), .B1(n_724), .B2(n_731), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_666), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_666), .A2(n_668), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_666), .A2(n_668), .B1(n_1367), .B2(n_1368), .Y(n_1366) );
OAI22xp5_ASAP7_75t_L g1377 ( .A1(n_666), .A2(n_691), .B1(n_1378), .B2(n_1379), .Y(n_1377) );
OAI22xp5_ASAP7_75t_SL g1096 ( .A1(n_668), .A2(n_1097), .B1(n_1098), .B2(n_1099), .Y(n_1096) );
OAI22xp33_ASAP7_75t_L g1205 ( .A1(n_668), .A2(n_942), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
OAI22xp33_ASAP7_75t_L g1215 ( .A1(n_668), .A2(n_942), .B1(n_1216), .B2(n_1217), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_670), .A2(n_690), .B1(n_701), .B2(n_703), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_671), .A2(n_675), .B1(n_1101), .B2(n_1102), .Y(n_1100) );
INVx1_ASAP7_75t_L g1374 ( .A(n_671), .Y(n_1374) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_672), .A2(n_693), .B1(n_703), .B2(n_705), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_673), .A2(n_677), .B1(n_1370), .B2(n_1371), .Y(n_1369) );
INVx5_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_675), .A2(n_677), .B1(n_680), .B2(n_681), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_675), .A2(n_677), .B1(n_717), .B2(n_735), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_675), .A2(n_788), .B1(n_805), .B2(n_814), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_675), .A2(n_811), .B1(n_844), .B2(n_845), .Y(n_843) );
BUFx2_ASAP7_75t_SL g1105 ( .A(n_675), .Y(n_1105) );
BUFx3_ASAP7_75t_L g1170 ( .A(n_675), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_675), .A2(n_1253), .B1(n_1263), .B2(n_1267), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_677), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx4_ASAP7_75t_L g743 ( .A(n_678), .Y(n_743) );
INVx2_ASAP7_75t_L g946 ( .A(n_678), .Y(n_946) );
INVx4_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI33xp33_ASAP7_75t_L g736 ( .A1(n_682), .A2(n_737), .A3(n_739), .B1(n_742), .B2(n_745), .B3(n_746), .Y(n_736) );
OAI33xp33_ASAP7_75t_L g1094 ( .A1(n_682), .A2(n_1095), .A3(n_1096), .B1(n_1100), .B2(n_1103), .B3(n_1107), .Y(n_1094) );
OAI33xp33_ASAP7_75t_L g1163 ( .A1(n_682), .A2(n_737), .A3(n_1164), .B1(n_1165), .B2(n_1166), .B3(n_1167), .Y(n_1163) );
OAI33xp33_ASAP7_75t_L g1365 ( .A1(n_682), .A2(n_737), .A3(n_1366), .B1(n_1369), .B2(n_1372), .B3(n_1377), .Y(n_1365) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_683), .Y(n_955) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_690), .B1(n_691), .B2(n_693), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g740 ( .A(n_688), .Y(n_740) );
INVx3_ASAP7_75t_L g942 ( .A(n_688), .Y(n_942) );
INVx2_ASAP7_75t_L g1716 ( .A(n_688), .Y(n_1716) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx4_ASAP7_75t_L g809 ( .A(n_689), .Y(n_809) );
INVx3_ASAP7_75t_L g1098 ( .A(n_689), .Y(n_1098) );
BUFx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI33xp33_ASAP7_75t_L g956 ( .A1(n_695), .A2(n_957), .A3(n_961), .B1(n_963), .B2(n_965), .B3(n_966), .Y(n_956) );
OAI33xp33_ASAP7_75t_L g1218 ( .A1(n_695), .A2(n_965), .A3(n_1219), .B1(n_1220), .B2(n_1222), .B3(n_1223), .Y(n_1218) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_697), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_697), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g1381 ( .A1(n_697), .A2(n_1367), .B1(n_1375), .B2(n_1382), .Y(n_1381) );
OAI22xp33_ASAP7_75t_L g1387 ( .A1(n_697), .A2(n_1148), .B1(n_1368), .B2(n_1376), .Y(n_1387) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_699), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g801 ( .A1(n_699), .A2(n_802), .B1(n_804), .B2(n_805), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_699), .A2(n_802), .B1(n_842), .B2(n_848), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g1082 ( .A1(n_699), .A2(n_802), .B1(n_1070), .B2(n_1076), .Y(n_1082) );
INVx2_ASAP7_75t_L g1116 ( .A(n_699), .Y(n_1116) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g1221 ( .A(n_702), .Y(n_1221) );
INVx1_ASAP7_75t_L g1384 ( .A(n_702), .Y(n_1384) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_703), .A2(n_945), .B1(n_952), .B2(n_962), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_703), .A2(n_856), .B1(n_1102), .B2(n_1109), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g1383 ( .A1(n_703), .A2(n_1370), .B1(n_1378), .B2(n_1384), .Y(n_1383) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_703), .A2(n_1371), .B1(n_1379), .B2(n_1386), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_705), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_705), .A2(n_794), .B1(n_844), .B2(n_850), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_705), .A2(n_1074), .B1(n_1080), .B2(n_1086), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1743 ( .A1(n_705), .A2(n_794), .B1(n_1744), .B2(n_1745), .Y(n_1743) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g959 ( .A(n_709), .Y(n_959) );
INVxp67_ASAP7_75t_SL g1114 ( .A(n_709), .Y(n_1114) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_747), .C(n_764), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_736), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g739 ( .A1(n_716), .A2(n_733), .B1(n_740), .B2(n_741), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_724), .B2(n_725), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_720), .A2(n_729), .B1(n_743), .B2(n_744), .Y(n_742) );
BUFx3_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx8_ASAP7_75t_L g1154 ( .A(n_722), .Y(n_1154) );
INVx5_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_SL g856 ( .A(n_723), .Y(n_856) );
INVx3_ASAP7_75t_L g1084 ( .A(n_723), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1289 ( .A(n_723), .Y(n_1289) );
OAI22xp33_ASAP7_75t_SL g1149 ( .A1(n_725), .A2(n_1084), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_725), .A2(n_1210), .B1(n_1216), .B2(n_1221), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_725), .A2(n_964), .B1(n_1211), .B2(n_1217), .Y(n_1222) );
INVx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g800 ( .A(n_727), .Y(n_800) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI33xp33_ASAP7_75t_L g838 ( .A1(n_738), .A2(n_816), .A3(n_839), .B1(n_843), .B2(n_846), .B3(n_849), .Y(n_838) );
OAI33xp33_ASAP7_75t_L g1068 ( .A1(n_738), .A2(n_816), .A3(n_1069), .B1(n_1072), .B2(n_1075), .B3(n_1078), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g1265 ( .A1(n_741), .A2(n_809), .B1(n_1252), .B2(n_1262), .Y(n_1265) );
OAI22xp33_ASAP7_75t_L g1165 ( .A1(n_743), .A2(n_819), .B1(n_1150), .B2(n_1155), .Y(n_1165) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_744), .A2(n_811), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1754 ( .A1(n_744), .A2(n_1267), .B1(n_1744), .B2(n_1747), .Y(n_1754) );
OAI31xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_751), .A3(n_759), .B(n_763), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVxp67_ASAP7_75t_SL g1148 ( .A(n_753), .Y(n_1148) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g830 ( .A(n_754), .Y(n_830) );
INVx1_ASAP7_75t_L g1399 ( .A(n_754), .Y(n_1399) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI31xp33_ASAP7_75t_L g977 ( .A1(n_763), .A2(n_978), .A3(n_979), .B(n_984), .Y(n_977) );
OAI31xp33_ASAP7_75t_L g1177 ( .A1(n_763), .A2(n_1178), .A3(n_1180), .B(n_1183), .Y(n_1177) );
OAI31xp33_ASAP7_75t_L g1194 ( .A1(n_763), .A2(n_1195), .A3(n_1196), .B(n_1201), .Y(n_1194) );
OAI31xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .A3(n_770), .B(n_773), .Y(n_764) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g926 ( .A(n_772), .Y(n_926) );
INVxp67_ASAP7_75t_SL g975 ( .A(n_772), .Y(n_975) );
OAI31xp33_ASAP7_75t_L g1186 ( .A1(n_773), .A2(n_1187), .A3(n_1192), .B(n_1193), .Y(n_1186) );
OAI31xp33_ASAP7_75t_SL g1232 ( .A1(n_773), .A2(n_1233), .A3(n_1238), .B(n_1239), .Y(n_1232) );
OAI21xp5_ASAP7_75t_L g1301 ( .A1(n_773), .A2(n_1302), .B(n_1310), .Y(n_1301) );
XNOR2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_1089), .Y(n_775) );
XOR2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_872), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
XNOR2x1_ASAP7_75t_L g779 ( .A(n_780), .B(n_835), .Y(n_779) );
XNOR2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
AND3x1_ASAP7_75t_L g782 ( .A(n_783), .B(n_817), .C(n_826), .Y(n_782) );
NOR2xp33_ASAP7_75t_SL g783 ( .A(n_784), .B(n_807), .Y(n_783) );
OAI33xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .A3(n_791), .B1(n_795), .B2(n_801), .B3(n_806), .Y(n_784) );
OAI33xp33_ASAP7_75t_L g852 ( .A1(n_785), .A2(n_806), .A3(n_853), .B1(n_854), .B2(n_855), .B3(n_857), .Y(n_852) );
OAI33xp33_ASAP7_75t_L g1081 ( .A1(n_785), .A2(n_806), .A3(n_1082), .B1(n_1083), .B2(n_1085), .B3(n_1087), .Y(n_1081) );
OAI33xp33_ASAP7_75t_L g1250 ( .A1(n_785), .A2(n_806), .A3(n_1251), .B1(n_1254), .B2(n_1257), .B3(n_1261), .Y(n_1250) );
OAI33xp33_ASAP7_75t_L g1325 ( .A1(n_785), .A2(n_806), .A3(n_1326), .B1(n_1329), .B2(n_1332), .B3(n_1335), .Y(n_1325) );
OAI33xp33_ASAP7_75t_L g1739 ( .A1(n_785), .A2(n_806), .A3(n_1740), .B1(n_1743), .B2(n_1746), .B3(n_1749), .Y(n_1739) );
OAI22xp33_ASAP7_75t_L g879 ( .A1(n_789), .A2(n_880), .B1(n_881), .B2(n_882), .Y(n_879) );
INVx3_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g967 ( .A(n_790), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_792), .A2(n_796), .B1(n_811), .B2(n_812), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_794), .A2(n_1073), .B1(n_1079), .B2(n_1084), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B1(n_799), .B2(n_800), .Y(n_795) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g962 ( .A(n_798), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_800), .A2(n_1258), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
INVx2_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
INVx3_ASAP7_75t_L g880 ( .A(n_803), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_809), .A2(n_840), .B1(n_841), .B2(n_842), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_809), .A2(n_841), .B1(n_1079), .B2(n_1080), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_812), .A2(n_1255), .B1(n_1259), .B2(n_1267), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g1340 ( .A1(n_812), .A2(n_1267), .B1(n_1330), .B2(n_1333), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_812), .A2(n_1267), .B1(n_1328), .B2(n_1337), .Y(n_1341) );
OAI33xp33_ASAP7_75t_L g895 ( .A1(n_816), .A2(n_896), .A3(n_898), .B1(n_900), .B2(n_901), .B3(n_902), .Y(n_895) );
OAI22xp33_ASAP7_75t_L g1120 ( .A1(n_829), .A2(n_1099), .B1(n_1106), .B2(n_1113), .Y(n_1120) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NAND3xp33_ASAP7_75t_SL g1008 ( .A(n_831), .B(n_1009), .C(n_1013), .Y(n_1008) );
NAND3xp33_ASAP7_75t_SL g1061 ( .A(n_831), .B(n_1062), .C(n_1064), .Y(n_1061) );
NAND3xp33_ASAP7_75t_L g1243 ( .A(n_831), .B(n_1244), .C(n_1246), .Y(n_1243) );
AND3x1_ASAP7_75t_L g836 ( .A(n_837), .B(n_858), .C(n_866), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_852), .Y(n_837) );
OAI22xp33_ASAP7_75t_L g940 ( .A1(n_841), .A2(n_941), .B1(n_942), .B2(n_943), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g1746 ( .A1(n_856), .A2(n_1086), .B1(n_1747), .B2(n_1748), .Y(n_1746) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_874), .B1(n_987), .B2(n_1088), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_935), .B1(n_936), .B2(n_986), .Y(n_874) );
INVx1_ASAP7_75t_L g986 ( .A(n_875), .Y(n_986) );
INVxp67_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
NOR4xp25_ASAP7_75t_L g934 ( .A(n_878), .B(n_895), .C(n_904), .D(n_923), .Y(n_934) );
BUFx4f_ASAP7_75t_SL g1146 ( .A(n_880), .Y(n_1146) );
INVxp67_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVxp67_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
AOI31xp33_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_912), .A3(n_916), .B(n_921), .Y(n_904) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g1136 ( .A(n_915), .Y(n_1136) );
AOI22xp5_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_916) );
INVx1_ASAP7_75t_L g1179 ( .A(n_918), .Y(n_1179) );
CKINVDCx14_ASAP7_75t_R g921 ( .A(n_922), .Y(n_921) );
AOI31xp67_ASAP7_75t_SL g923 ( .A1(n_924), .A2(n_927), .A3(n_931), .B(n_933), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g1190 ( .A(n_930), .Y(n_1190) );
INVxp67_ASAP7_75t_SL g931 ( .A(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g937 ( .A(n_938), .B(n_968), .C(n_977), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_956), .Y(n_938) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_941), .A2(n_949), .B1(n_958), .B2(n_960), .Y(n_957) );
OAI22xp33_ASAP7_75t_L g966 ( .A1(n_943), .A2(n_950), .B1(n_958), .B2(n_967), .Y(n_966) );
OAI33xp33_ASAP7_75t_L g1204 ( .A1(n_955), .A2(n_1205), .A3(n_1208), .B1(n_1209), .B2(n_1212), .B3(n_1215), .Y(n_1204) );
OAI22xp33_ASAP7_75t_L g1219 ( .A1(n_958), .A2(n_967), .B1(n_1206), .B2(n_1213), .Y(n_1219) );
INVx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g1354 ( .A(n_982), .Y(n_1354) );
INVx2_ASAP7_75t_L g1088 ( .A(n_987), .Y(n_1088) );
XNOR2x1_ASAP7_75t_L g987 ( .A(n_988), .B(n_1050), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_989), .B(n_1032), .Y(n_988) );
INVx1_ASAP7_75t_L g1034 ( .A(n_990), .Y(n_1034) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_992), .B(n_998), .Y(n_990) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
NAND3xp33_ASAP7_75t_L g1287 ( .A(n_996), .B(n_1288), .C(n_1291), .Y(n_1287) );
BUFx3_ASAP7_75t_L g1662 ( .A(n_996), .Y(n_1662) );
OAI221xp5_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1002), .B1(n_1003), .B2(n_1004), .C(n_1005), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_1001), .Y(n_1247) );
INVx2_ASAP7_75t_L g1664 ( .A(n_1003), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_1006), .B(n_1018), .Y(n_1033) );
OAI31xp33_ASAP7_75t_SL g1006 ( .A1(n_1007), .A2(n_1008), .A3(n_1016), .B(n_1017), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .Y(n_1009) );
INVx2_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1012), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1015), .B(n_1028), .Y(n_1027) );
OAI31xp33_ASAP7_75t_SL g1059 ( .A1(n_1017), .A2(n_1060), .A3(n_1061), .B(n_1066), .Y(n_1059) );
AO21x1_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1023), .B(n_1031), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .Y(n_1023) );
NAND3xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .C(n_1030), .Y(n_1025) );
INVx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
OAI31xp33_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1034), .A3(n_1035), .B(n_1047), .Y(n_1032) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1036), .Y(n_1049) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1044), .Y(n_1281) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1049), .Y(n_1047) );
NAND3xp33_ASAP7_75t_SL g1051 ( .A(n_1052), .B(n_1059), .C(n_1067), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1057), .B(n_1063), .Y(n_1062) );
NOR2xp33_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1081), .Y(n_1067) );
XNOR2xp5_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1138), .Y(n_1089) );
INVx2_ASAP7_75t_SL g1090 ( .A(n_1091), .Y(n_1090) );
NAND3xp33_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1121), .C(n_1130), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1110), .Y(n_1093) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_1097), .A2(n_1104), .B1(n_1113), .B2(n_1115), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_1105), .A2(n_1373), .B1(n_1375), .B2(n_1376), .Y(n_1372) );
OAI33xp33_ASAP7_75t_L g1110 ( .A1(n_1111), .A2(n_1112), .A3(n_1117), .B1(n_1118), .B2(n_1119), .B3(n_1120), .Y(n_1110) );
OAI33xp33_ASAP7_75t_L g1143 ( .A1(n_1111), .A2(n_1144), .A3(n_1149), .B1(n_1152), .B2(n_1157), .B3(n_1160), .Y(n_1143) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
OAI31xp33_ASAP7_75t_L g1121 ( .A1(n_1122), .A2(n_1123), .A3(n_1128), .B(n_1129), .Y(n_1121) );
OAI31xp33_ASAP7_75t_SL g1168 ( .A1(n_1129), .A2(n_1169), .A3(n_1174), .B(n_1176), .Y(n_1168) );
OAI31xp33_ASAP7_75t_L g1388 ( .A1(n_1129), .A2(n_1389), .A3(n_1393), .B(n_1394), .Y(n_1388) );
OAI31xp33_ASAP7_75t_L g1130 ( .A1(n_1131), .A2(n_1132), .A3(n_1135), .B(n_1137), .Y(n_1130) );
OAI31xp33_ASAP7_75t_L g1395 ( .A1(n_1137), .A2(n_1396), .A3(n_1397), .B(n_1402), .Y(n_1395) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1184), .B1(n_1224), .B2(n_1225), .Y(n_1138) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1139), .Y(n_1224) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
NAND3xp33_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1168), .C(n_1177), .Y(n_1141) );
NOR2xp33_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1163), .Y(n_1142) );
OAI22xp33_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1146), .B1(n_1147), .B2(n_1148), .Y(n_1144) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
AOI33xp33_ASAP7_75t_L g1661 ( .A1(n_1158), .A2(n_1662), .A3(n_1663), .B1(n_1665), .B2(n_1666), .B3(n_1668), .Y(n_1661) );
BUFx2_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
BUFx2_ASAP7_75t_L g1299 ( .A(n_1159), .Y(n_1299) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1184), .Y(n_1225) );
NAND3xp33_ASAP7_75t_SL g1185 ( .A(n_1186), .B(n_1194), .C(n_1203), .Y(n_1185) );
INVx2_ASAP7_75t_SL g1197 ( .A(n_1198), .Y(n_1197) );
NOR2xp33_ASAP7_75t_SL g1203 ( .A(n_1204), .B(n_1218), .Y(n_1203) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_1228), .A2(n_1229), .B1(n_1318), .B2(n_1319), .Y(n_1227) );
INVx2_ASAP7_75t_SL g1228 ( .A(n_1229), .Y(n_1228) );
XNOR2x1_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1272), .Y(n_1229) );
NAND3xp33_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1240), .C(n_1249), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1237), .B(n_1247), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1264), .Y(n_1249) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
NAND3xp33_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1301), .C(n_1311), .Y(n_1273) );
AND4x1_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1283), .C(n_1287), .D(n_1296), .Y(n_1274) );
NAND3xp33_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1280), .C(n_1282), .Y(n_1275) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
NAND3xp33_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1299), .C(n_1300), .Y(n_1296) );
BUFx2_ASAP7_75t_L g1667 ( .A(n_1298), .Y(n_1667) );
INVx2_ASAP7_75t_SL g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
AOI22xp5_ASAP7_75t_L g1319 ( .A1(n_1320), .A2(n_1321), .B1(n_1362), .B2(n_1403), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
NAND3xp33_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1343), .C(n_1351), .Y(n_1323) );
NOR2xp33_ASAP7_75t_SL g1324 ( .A(n_1325), .B(n_1338), .Y(n_1324) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1357), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1358), .B(n_1645), .Y(n_1644) );
INVx3_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1362), .Y(n_1403) );
NAND3xp33_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1388), .C(n_1395), .Y(n_1363) );
NOR2xp33_ASAP7_75t_SL g1364 ( .A(n_1365), .B(n_1380), .Y(n_1364) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVxp67_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
OAI221xp5_ASAP7_75t_L g1404 ( .A1(n_1405), .A2(n_1624), .B1(n_1626), .B2(n_1725), .C(n_1728), .Y(n_1404) );
AOI211xp5_ASAP7_75t_L g1405 ( .A1(n_1406), .A2(n_1529), .B(n_1536), .C(n_1602), .Y(n_1405) );
NAND5xp2_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1480), .C(n_1507), .D(n_1510), .E(n_1515), .Y(n_1406) );
AOI211xp5_ASAP7_75t_L g1407 ( .A1(n_1408), .A2(n_1438), .B(n_1447), .C(n_1475), .Y(n_1407) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
OR2x2_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1425), .Y(n_1409) );
OAI321xp33_ASAP7_75t_L g1447 ( .A1(n_1410), .A2(n_1448), .A3(n_1455), .B1(n_1460), .B2(n_1461), .C(n_1466), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1410), .B(n_1426), .Y(n_1468) );
AND3x1_ASAP7_75t_L g1501 ( .A(n_1410), .B(n_1435), .C(n_1459), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1410), .B(n_1493), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1526 ( .A(n_1410), .B(n_1435), .Y(n_1526) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1410), .B(n_1554), .Y(n_1553) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1410), .B(n_1456), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1410), .B(n_1459), .Y(n_1595) );
INVx2_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1411), .B(n_1456), .Y(n_1465) );
BUFx2_ASAP7_75t_L g1471 ( .A(n_1411), .Y(n_1471) );
OR2x2_ASAP7_75t_L g1562 ( .A(n_1411), .B(n_1548), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1411), .B(n_1493), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1420), .Y(n_1411) );
AND2x4_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1415), .Y(n_1413) );
AND2x6_ASAP7_75t_L g1418 ( .A(n_1414), .B(n_1419), .Y(n_1418) );
AND2x6_ASAP7_75t_L g1421 ( .A(n_1414), .B(n_1422), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1414), .B(n_1424), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1414), .B(n_1424), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1414), .B(n_1424), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1417), .Y(n_1415) );
INVx2_ASAP7_75t_L g1533 ( .A(n_1421), .Y(n_1533) );
OAI21xp5_ASAP7_75t_L g1772 ( .A1(n_1422), .A2(n_1773), .B(n_1774), .Y(n_1772) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1431), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1426), .B(n_1450), .Y(n_1449) );
NOR2xp33_ASAP7_75t_L g1483 ( .A(n_1426), .B(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1426), .Y(n_1518) );
NAND2xp5_ASAP7_75t_L g1544 ( .A(n_1426), .B(n_1488), .Y(n_1544) );
NOR2xp33_ASAP7_75t_L g1578 ( .A(n_1426), .B(n_1579), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1613 ( .A(n_1426), .B(n_1456), .Y(n_1613) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1427), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1427), .B(n_1471), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1427), .B(n_1440), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1548 ( .A(n_1427), .B(n_1431), .Y(n_1548) );
NOR2xp33_ASAP7_75t_L g1550 ( .A(n_1427), .B(n_1551), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1427), .B(n_1451), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1428), .B(n_1429), .Y(n_1427) );
INVxp67_ASAP7_75t_L g1535 ( .A(n_1430), .Y(n_1535) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1431), .B(n_1470), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1435), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1432), .B(n_1457), .Y(n_1456) );
INVx2_ASAP7_75t_L g1459 ( .A(n_1432), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1432), .B(n_1471), .Y(n_1484) );
NAND3xp33_ASAP7_75t_L g1557 ( .A(n_1432), .B(n_1462), .C(n_1530), .Y(n_1557) );
OR2x2_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1434), .Y(n_1432) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1435), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1435), .B(n_1459), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1435), .B(n_1471), .Y(n_1543) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1435), .B(n_1471), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1437), .Y(n_1435) );
A2O1A1Ixp33_ASAP7_75t_L g1546 ( .A1(n_1438), .A2(n_1530), .B(n_1547), .C(n_1549), .Y(n_1546) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
OR2x2_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1444), .Y(n_1439) );
CKINVDCx6p67_ASAP7_75t_R g1473 ( .A(n_1440), .Y(n_1473) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_1440), .B(n_1478), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1520 ( .A(n_1440), .B(n_1488), .Y(n_1520) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1440), .B(n_1444), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1610 ( .A(n_1440), .B(n_1530), .Y(n_1610) );
NAND2xp5_ASAP7_75t_L g1617 ( .A(n_1440), .B(n_1618), .Y(n_1617) );
OR2x6_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1443), .Y(n_1440) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1444), .Y(n_1454) );
INVx3_ASAP7_75t_L g1460 ( .A(n_1444), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1444), .B(n_1474), .Y(n_1479) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_1444), .B(n_1451), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1444), .B(n_1473), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1444), .B(n_1451), .Y(n_1497) );
OR2x2_ASAP7_75t_L g1512 ( .A(n_1444), .B(n_1473), .Y(n_1512) );
OAI221xp5_ASAP7_75t_L g1571 ( .A1(n_1444), .A2(n_1572), .B1(n_1573), .B2(n_1575), .C(n_1576), .Y(n_1571) );
OAI32xp33_ASAP7_75t_L g1598 ( .A1(n_1444), .A2(n_1460), .A3(n_1462), .B1(n_1553), .B2(n_1599), .Y(n_1598) );
AND2x4_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1446), .Y(n_1444) );
OAI32xp33_ASAP7_75t_L g1615 ( .A1(n_1448), .A2(n_1462), .A3(n_1502), .B1(n_1616), .B2(n_1617), .Y(n_1615) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1450), .Y(n_1502) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1450), .B(n_1473), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1454), .Y(n_1450) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1451), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1453), .Y(n_1451) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1458), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1456), .B(n_1470), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1457), .B(n_1459), .Y(n_1493) );
O2A1O1Ixp33_ASAP7_75t_L g1566 ( .A1(n_1457), .A2(n_1567), .B(n_1568), .C(n_1569), .Y(n_1566) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1458), .B(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1458), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1458), .B(n_1471), .Y(n_1514) );
OAI322xp33_ASAP7_75t_L g1495 ( .A1(n_1459), .A2(n_1496), .A3(n_1498), .B1(n_1500), .B2(n_1502), .C1(n_1503), .C2(n_1505), .Y(n_1495) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1459), .B(n_1471), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1459), .B(n_1471), .Y(n_1600) );
CKINVDCx14_ASAP7_75t_R g1591 ( .A(n_1460), .Y(n_1591) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1465), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1588 ( .A(n_1462), .B(n_1556), .Y(n_1588) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1463), .B(n_1506), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1463), .B(n_1504), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1463), .B(n_1556), .Y(n_1585) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1464), .B(n_1514), .Y(n_1513) );
NAND2xp5_ASAP7_75t_L g1554 ( .A(n_1464), .B(n_1493), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1464), .B(n_1504), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1621 ( .A(n_1465), .B(n_1488), .Y(n_1621) );
OAI21xp5_ASAP7_75t_L g1466 ( .A1(n_1467), .A2(n_1469), .B(n_1472), .Y(n_1466) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1467), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1468), .B(n_1493), .Y(n_1523) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1469), .Y(n_1608) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1470), .Y(n_1491) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1472), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_1472), .B(n_1574), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1474), .Y(n_1472) );
NOR2xp33_ASAP7_75t_L g1481 ( .A(n_1473), .B(n_1482), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_1473), .B(n_1504), .Y(n_1503) );
NOR2xp33_ASAP7_75t_SL g1565 ( .A(n_1473), .B(n_1502), .Y(n_1565) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1473), .B(n_1530), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1473), .B(n_1488), .Y(n_1583) );
INVx2_ASAP7_75t_L g1488 ( .A(n_1474), .Y(n_1488) );
NOR2xp33_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1477), .Y(n_1475) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1477), .Y(n_1614) );
OAI22xp5_ASAP7_75t_L g1581 ( .A1(n_1478), .A2(n_1553), .B1(n_1582), .B2(n_1584), .Y(n_1581) );
OAI211xp5_ASAP7_75t_L g1589 ( .A1(n_1478), .A2(n_1555), .B(n_1590), .C(n_1596), .Y(n_1589) );
CKINVDCx6p67_ASAP7_75t_R g1478 ( .A(n_1479), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1479), .B(n_1518), .Y(n_1517) );
AOI221xp5_ASAP7_75t_L g1480 ( .A1(n_1481), .A2(n_1483), .B1(n_1485), .B2(n_1494), .C(n_1495), .Y(n_1480) );
INVx2_ASAP7_75t_L g1504 ( .A(n_1482), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1486), .B(n_1489), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1486), .B(n_1578), .Y(n_1577) );
A2O1A1Ixp33_ASAP7_75t_L g1605 ( .A1(n_1486), .A2(n_1554), .B(n_1555), .C(n_1606), .Y(n_1605) );
INVx2_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
NAND2xp5_ASAP7_75t_L g1507 ( .A(n_1487), .B(n_1508), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1527 ( .A(n_1487), .B(n_1528), .Y(n_1527) );
NOR2xp33_ASAP7_75t_L g1607 ( .A(n_1487), .B(n_1608), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1487), .B(n_1585), .Y(n_1623) );
INVx2_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1572 ( .A(n_1488), .B(n_1490), .Y(n_1572) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
OR2x2_ASAP7_75t_L g1490 ( .A(n_1491), .B(n_1492), .Y(n_1490) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1494), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1494), .B(n_1550), .Y(n_1549) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_1496), .A2(n_1522), .B1(n_1524), .B2(n_1527), .Y(n_1521) );
NOR2xp33_ASAP7_75t_L g1597 ( .A(n_1496), .B(n_1500), .Y(n_1597) );
INVx2_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_1497), .A2(n_1501), .B1(n_1564), .B2(n_1565), .Y(n_1563) );
CKINVDCx14_ASAP7_75t_R g1498 ( .A(n_1499), .Y(n_1498) );
INVx2_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
O2A1O1Ixp33_ASAP7_75t_L g1611 ( .A1(n_1508), .A2(n_1612), .B(n_1614), .C(n_1615), .Y(n_1611) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1513), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
O2A1O1Ixp33_ASAP7_75t_L g1515 ( .A1(n_1514), .A2(n_1516), .B(n_1519), .C(n_1521), .Y(n_1515) );
NOR2xp33_ASAP7_75t_L g1616 ( .A(n_1514), .B(n_1556), .Y(n_1616) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
NOR2xp33_ASAP7_75t_L g1525 ( .A(n_1518), .B(n_1526), .Y(n_1525) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
OAI221xp5_ASAP7_75t_L g1538 ( .A1(n_1520), .A2(n_1539), .B1(n_1540), .B2(n_1545), .C(n_1546), .Y(n_1538) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
OAI31xp33_ASAP7_75t_L g1619 ( .A1(n_1528), .A2(n_1620), .A3(n_1621), .B(n_1622), .Y(n_1619) );
INVx2_ASAP7_75t_SL g1529 ( .A(n_1530), .Y(n_1529) );
INVx2_ASAP7_75t_SL g1575 ( .A(n_1530), .Y(n_1575) );
OAI22xp5_ASAP7_75t_SL g1531 ( .A1(n_1532), .A2(n_1533), .B1(n_1534), .B2(n_1535), .Y(n_1531) );
CKINVDCx20_ASAP7_75t_R g1625 ( .A(n_1533), .Y(n_1625) );
NAND3xp33_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1570), .C(n_1586), .Y(n_1536) );
NOR4xp25_ASAP7_75t_L g1537 ( .A(n_1538), .B(n_1552), .C(n_1560), .D(n_1566), .Y(n_1537) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1541), .Y(n_1540) );
OAI21xp5_ASAP7_75t_L g1576 ( .A1(n_1541), .A2(n_1577), .B(n_1580), .Y(n_1576) );
NOR2xp33_ASAP7_75t_L g1541 ( .A(n_1542), .B(n_1544), .Y(n_1541) );
A2O1A1Ixp33_ASAP7_75t_L g1603 ( .A1(n_1542), .A2(n_1604), .B(n_1605), .C(n_1609), .Y(n_1603) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
AOI31xp33_ASAP7_75t_L g1552 ( .A1(n_1553), .A2(n_1555), .A3(n_1557), .B(n_1558), .Y(n_1552) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1553), .Y(n_1620) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
OAI21xp33_ASAP7_75t_L g1560 ( .A1(n_1561), .A2(n_1562), .B(n_1563), .Y(n_1560) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1564), .Y(n_1568) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1569), .Y(n_1580) );
NOR2xp33_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1581), .Y(n_1570) );
INVx3_ASAP7_75t_L g1601 ( .A(n_1575), .Y(n_1601) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
OAI31xp33_ASAP7_75t_L g1586 ( .A1(n_1587), .A2(n_1589), .A3(n_1598), .B(n_1601), .Y(n_1586) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1592), .Y(n_1590) );
NOR2xp33_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1595), .Y(n_1592) );
CKINVDCx14_ASAP7_75t_R g1593 ( .A(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1595), .Y(n_1618) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
CKINVDCx14_ASAP7_75t_R g1599 ( .A(n_1600), .Y(n_1599) );
NAND3xp33_ASAP7_75t_L g1602 ( .A(n_1603), .B(n_1611), .C(n_1619), .Y(n_1602) );
INVxp67_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
CKINVDCx20_ASAP7_75t_R g1624 ( .A(n_1625), .Y(n_1624) );
INVx2_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
XOR2x2_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1724), .Y(n_1627) );
NAND2xp5_ASAP7_75t_SL g1628 ( .A(n_1629), .B(n_1685), .Y(n_1628) );
AOI211x1_ASAP7_75t_L g1629 ( .A1(n_1630), .A2(n_1631), .B(n_1640), .C(n_1673), .Y(n_1629) );
INVx8_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
AND2x4_ASAP7_75t_L g1632 ( .A(n_1633), .B(n_1636), .Y(n_1632) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1634), .Y(n_1682) );
OR2x2_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1638), .Y(n_1636) );
AND2x4_ASAP7_75t_L g1645 ( .A(n_1637), .B(n_1646), .Y(n_1645) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1639), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1641), .B(n_1661), .Y(n_1640) );
NOR2xp33_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1652), .Y(n_1641) );
AO22x1_ASAP7_75t_L g1642 ( .A1(n_1643), .A2(n_1644), .B1(n_1648), .B2(n_1649), .Y(n_1642) );
AND2x4_ASAP7_75t_L g1649 ( .A(n_1645), .B(n_1650), .Y(n_1649) );
INVx2_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
NAND2xp5_ASAP7_75t_SL g1652 ( .A(n_1653), .B(n_1659), .Y(n_1652) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1654), .B(n_1655), .Y(n_1653) );
NAND2xp5_ASAP7_75t_R g1703 ( .A(n_1654), .B(n_1704), .Y(n_1703) );
INVx5_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
OR2x6_ASAP7_75t_L g1656 ( .A(n_1657), .B(n_1658), .Y(n_1656) );
INVx3_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
AND2x4_ASAP7_75t_L g1674 ( .A(n_1675), .B(n_1677), .Y(n_1674) );
AOI22xp33_ASAP7_75t_L g1678 ( .A1(n_1679), .A2(n_1680), .B1(n_1683), .B2(n_1684), .Y(n_1678) );
AOI22xp33_ASAP7_75t_L g1687 ( .A1(n_1679), .A2(n_1683), .B1(n_1688), .B2(n_1692), .Y(n_1687) );
AND2x4_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1682), .Y(n_1680) );
OAI21xp5_ASAP7_75t_L g1685 ( .A1(n_1686), .A2(n_1706), .B(n_1723), .Y(n_1685) );
NAND3xp33_ASAP7_75t_SL g1686 ( .A(n_1687), .B(n_1693), .C(n_1703), .Y(n_1686) );
INVx2_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
AND2x4_ASAP7_75t_L g1704 ( .A(n_1691), .B(n_1705), .Y(n_1704) );
AOI21xp5_ASAP7_75t_L g1693 ( .A1(n_1694), .A2(n_1699), .B(n_1702), .Y(n_1693) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
INVx1_ASAP7_75t_SL g1700 ( .A(n_1701), .Y(n_1700) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
INVx4_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
INVx2_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
BUFx2_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
INVx2_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
NOR2x1_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1722), .Y(n_1720) );
CKINVDCx5p33_ASAP7_75t_R g1725 ( .A(n_1726), .Y(n_1725) );
HB1xp67_ASAP7_75t_SL g1729 ( .A(n_1730), .Y(n_1729) );
BUFx3_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
INVxp33_ASAP7_75t_SL g1732 ( .A(n_1733), .Y(n_1732) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
HB1xp67_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
NAND3xp33_ASAP7_75t_L g1737 ( .A(n_1738), .B(n_1757), .C(n_1764), .Y(n_1737) );
NOR2xp33_ASAP7_75t_SL g1738 ( .A(n_1739), .B(n_1752), .Y(n_1738) );
HB1xp67_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
INVx1_ASAP7_75t_L g1774 ( .A(n_1775), .Y(n_1774) );
endmodule