module fake_ibex_75_n_7892 (n_151, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_343, n_310, n_714, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_1052, n_852, n_789, n_880, n_654, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_1048, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_7892);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_343;
input n_310;
input n_714;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_7892;

wire n_4557;
wire n_6873;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_7170;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_7029;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_7042;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_7262;
wire n_7551;
wire n_6616;
wire n_6848;
wire n_4371;
wire n_7766;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_7063;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_6744;
wire n_7707;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_7589;
wire n_6229;
wire n_7643;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_7792;
wire n_5615;
wire n_1480;
wire n_7147;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_7067;
wire n_7816;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_6658;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_6842;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_7485;
wire n_5922;
wire n_1981;
wire n_7636;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_7450;
wire n_7492;
wire n_6760;
wire n_7396;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_7082;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_7313;
wire n_7305;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_7332;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_7673;
wire n_1778;
wire n_7151;
wire n_2839;
wire n_7013;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_7672;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_7776;
wire n_6602;
wire n_7753;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_7885;
wire n_1960;
wire n_6562;
wire n_7397;
wire n_3979;
wire n_7324;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_7105;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_7560;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_7187;
wire n_4854;
wire n_6732;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_7229;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6674;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_7099;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_7251;
wire n_7189;
wire n_1078;
wire n_4422;
wire n_5743;
wire n_6868;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_7706;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_7507;
wire n_1305;
wire n_2088;
wire n_6724;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_7097;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_7241;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_7264;
wire n_7841;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_7372;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_7855;
wire n_7607;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_7521;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_6926;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_7628;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_7888;
wire n_6638;
wire n_7358;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_6878;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_7316;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_7207;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_7112;
wire n_7083;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_7889;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_7026;
wire n_3572;
wire n_6114;
wire n_6996;
wire n_1121;
wire n_4823;
wire n_7366;
wire n_5195;
wire n_7657;
wire n_5541;
wire n_7033;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_7103;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_6864;
wire n_1781;
wire n_4331;
wire n_7733;
wire n_2028;
wire n_3678;
wire n_7790;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_7711;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_7858;
wire n_5252;
wire n_6209;
wire n_7445;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_6941;
wire n_1271;
wire n_6011;
wire n_7667;
wire n_3416;
wire n_6824;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_7140;
wire n_4225;
wire n_7169;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_7813;
wire n_6540;
wire n_4489;
wire n_6912;
wire n_3455;
wire n_6940;
wire n_1591;
wire n_7048;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_7303;
wire n_7883;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_7192;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_7639;
wire n_3365;
wire n_4974;
wire n_6802;
wire n_4725;
wire n_6691;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_7394;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_6855;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_7003;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_7161;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_7723;
wire n_7748;
wire n_6958;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_7226;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6711;
wire n_6124;
wire n_3352;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_7356;
wire n_5199;
wire n_7377;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_7315;
wire n_7360;
wire n_7804;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_7081;
wire n_6136;
wire n_7559;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_7446;
wire n_1201;
wire n_5859;
wire n_7822;
wire n_7224;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_7541;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_7583;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_7131;
wire n_2440;
wire n_4113;
wire n_7777;
wire n_1440;
wire n_4646;
wire n_7155;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6971;
wire n_7553;
wire n_6128;
wire n_2361;
wire n_6804;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_7700;
wire n_3932;
wire n_2339;
wire n_7338;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_7221;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_6714;
wire n_4114;
wire n_6983;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_6857;
wire n_4209;
wire n_3692;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_7793;
wire n_3535;
wire n_6859;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_7101;
wire n_2954;
wire n_6379;
wire n_6911;
wire n_6766;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_7692;
wire n_7173;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6893;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_7530;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_7729;
wire n_7349;
wire n_7830;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6850;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_5385;
wire n_3441;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_7749;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_7690;
wire n_1864;
wire n_7884;
wire n_6827;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_7068;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_6699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_6901;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_6773;
wire n_4416;
wire n_7430;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6765;
wire n_7703;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_7391;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_7695;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_7283;
wire n_2884;
wire n_3383;
wire n_7148;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_6704;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_7592;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_7254;
wire n_2654;
wire n_7199;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_7509;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_6939;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_6727;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_6883;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_7457;
wire n_3257;
wire n_2459;
wire n_6652;
wire n_2439;
wire n_7619;
wire n_7875;
wire n_7760;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_6950;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_7327;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6915;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_7025;
wire n_1845;
wire n_3835;
wire n_7645;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_6922;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6731;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_7090;
wire n_1857;
wire n_7587;
wire n_7574;
wire n_1997;
wire n_7174;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_7250;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_6902;
wire n_1834;
wire n_3372;
wire n_7641;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_6837;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_6767;
wire n_7102;
wire n_4858;
wire n_6733;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_6723;
wire n_3339;
wire n_7177;
wire n_6900;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_7539;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_7797;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_7233;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_7742;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_7031;
wire n_1517;
wire n_5973;
wire n_7012;
wire n_7238;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_7030;
wire n_7110;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_6856;
wire n_5770;
wire n_1763;
wire n_6976;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_6682;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_7517;
wire n_2516;
wire n_2031;
wire n_7121;
wire n_1348;
wire n_7317;
wire n_1191;
wire n_4099;
wire n_7190;
wire n_3899;
wire n_6153;
wire n_7879;
wire n_4729;
wire n_5957;
wire n_7429;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_6777;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_7390;
wire n_2410;
wire n_7145;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_7787;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_7561;
wire n_7529;
wire n_6185;
wire n_6706;
wire n_5342;
wire n_6884;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_7868;
wire n_3277;
wire n_7533;
wire n_2758;
wire n_5787;
wire n_6745;
wire n_7210;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_7563;
wire n_4022;
wire n_5843;
wire n_1072;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_7191;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_7807;
wire n_1278;
wire n_2059;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_6881;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_7136;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_7213;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_4583;
wire n_7034;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_6990;
wire n_3650;
wire n_6948;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_6816;
wire n_7512;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_6712;
wire n_5824;
wire n_6280;
wire n_7682;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_7098;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_6656;
wire n_7323;
wire n_7806;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_7149;
wire n_7219;
wire n_4919;
wire n_7320;
wire n_7175;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1878;
wire n_1374;
wire n_7357;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_7593;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_7449;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_7663;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_7218;
wire n_6863;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_7292;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_6152;
wire n_7582;
wire n_2574;
wire n_7659;
wire n_7142;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_7428;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_6805;
wire n_5260;
wire n_6416;
wire n_7602;
wire n_5069;
wire n_2364;
wire n_7133;
wire n_2641;
wire n_7306;
wire n_1077;
wire n_7202;
wire n_6771;
wire n_4751;
wire n_7730;
wire n_5930;
wire n_5309;
wire n_6695;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_7691;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_2266;
wire n_4473;
wire n_6673;
wire n_7138;
wire n_7370;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_6978;
wire n_7626;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_6910;
wire n_2394;
wire n_1572;
wire n_7236;
wire n_1245;
wire n_7877;
wire n_4867;
wire n_7387;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_7122;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_7886;
wire n_6347;
wire n_7812;
wire n_6482;
wire n_7698;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_6925;
wire n_7024;
wire n_6483;
wire n_4686;
wire n_7466;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_6800;
wire n_7410;
wire n_5186;
wire n_7257;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6944;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_6980;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_7282;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_7495;
wire n_7334;
wire n_3068;
wire n_3071;
wire n_3919;
wire n_3683;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_7346;
wire n_5267;
wire n_7649;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_7532;
wire n_7740;
wire n_6432;
wire n_6426;
wire n_7847;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_7401;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_7245;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_6946;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_6897;
wire n_2982;
wire n_2634;
wire n_3124;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_7843;
wire n_7075;
wire n_7710;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6847;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5265;
wire n_5087;
wire n_4401;
wire n_4727;
wire n_7367;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_6737;
wire n_3005;
wire n_4627;
wire n_6936;
wire n_5107;
wire n_6780;
wire n_4309;
wire n_4027;
wire n_7132;
wire n_7486;
wire n_6758;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_7419;
wire n_2279;
wire n_1536;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_7201;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_7555;
wire n_1736;
wire n_6176;
wire n_7265;
wire n_7232;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_7023;
wire n_3675;
wire n_7227;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_7789;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_7642;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_7273;
wire n_7853;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_7623;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_7774;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_6909;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_7852;
wire n_6418;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_7070;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_6989;
wire n_2510;
wire n_7634;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6662;
wire n_6461;
wire n_7046;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_7801;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_7194;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_7527;
wire n_7290;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_7146;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_6960;
wire n_1226;
wire n_7834;
wire n_7253;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_7615;
wire n_3931;
wire n_5745;
wire n_7434;
wire n_4421;
wire n_2322;
wire n_7477;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_7452;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_6823;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_7414;
wire n_2485;
wire n_5614;
wire n_7802;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_6725;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_7475;
wire n_7775;
wire n_7835;
wire n_7184;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_6914;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_7152;
wire n_4771;
wire n_4970;
wire n_4652;
wire n_6927;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_6916;
wire n_6973;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_7554;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_7114;
wire n_6566;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_7354;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_6808;
wire n_7609;
wire n_7037;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_7709;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_6747;
wire n_7335;
wire n_3856;
wire n_6496;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_7849;
wire n_2273;
wire n_5428;
wire n_7823;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_6787;
wire n_1970;
wire n_3946;
wire n_7183;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_6784;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_7433;
wire n_2269;
wire n_6741;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_7669;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_2663;
wire n_3882;
wire n_6807;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_6795;
wire n_7437;
wire n_6898;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_6785;
wire n_7384;
wire n_7588;
wire n_6738;
wire n_3030;
wire n_5631;
wire n_6818;
wire n_5983;
wire n_7516;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_7393;
wire n_4517;
wire n_6021;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_6966;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_7796;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_6899;
wire n_4850;
wire n_1869;
wire n_7614;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_7503;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_6754;
wire n_4067;
wire n_6822;
wire n_6849;
wire n_6796;
wire n_6836;
wire n_4997;
wire n_5906;
wire n_7355;
wire n_6755;
wire n_7608;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_7084;
wire n_5916;
wire n_7685;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_7515;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_7483;
wire n_6476;
wire n_5828;
wire n_7648;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_6669;
wire n_5357;
wire n_6717;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_6988;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_7256;
wire n_3573;
wire n_7652;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_7172;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_7851;
wire n_7117;
wire n_1709;
wire n_6655;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_7821;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_6790;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_7828;
wire n_4206;
wire n_5273;
wire n_7722;
wire n_7874;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_5877;
wire n_2033;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_6840;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_7287;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_6748;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6676;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_7301;
wire n_6448;
wire n_3684;
wire n_6667;
wire n_1318;
wire n_4006;
wire n_7826;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_7819;
wire n_7786;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_7156;
wire n_1772;
wire n_2858;
wire n_7780;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_7857;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_6993;
wire n_2390;
wire n_7544;
wire n_7203;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_6653;
wire n_3098;
wire n_7732;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_7658;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_7408;
wire n_7605;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_7476;
wire n_7624;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_7566;
wire n_4462;
wire n_1153;
wire n_6560;
wire n_7307;
wire n_2787;
wire n_4540;
wire n_6987;
wire n_4187;
wire n_7684;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_7409;
wire n_7087;
wire n_3503;
wire n_2441;
wire n_7280;
wire n_7680;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_7107;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_6984;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6701;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_7288;
wire n_7248;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_6907;
wire n_4554;
wire n_1260;
wire n_7038;
wire n_4097;
wire n_4861;
wire n_7833;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_6661;
wire n_6730;
wire n_7860;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_7153;
wire n_5194;
wire n_7230;
wire n_4579;
wire n_7838;
wire n_5628;
wire n_6994;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_7572;
wire n_1593;
wire n_7308;
wire n_1775;
wire n_6889;
wire n_6361;
wire n_6803;
wire n_7481;
wire n_2570;
wire n_4025;
wire n_6751;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_7403;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_7369;
wire n_5630;
wire n_7800;
wire n_3136;
wire n_3108;
wire n_6696;
wire n_2395;
wire n_7089;
wire n_6062;
wire n_4059;
wire n_7258;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_6943;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_6252;
wire n_7080;
wire n_7718;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_7002;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_7745;
wire n_6726;
wire n_7689;
wire n_3238;
wire n_6740;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_6799;
wire n_2463;
wire n_6932;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_7008;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_7049;
wire n_1251;
wire n_6657;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_7062;
wire n_7493;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_6716;
wire n_6797;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_7215;
wire n_7340;
wire n_4822;
wire n_6694;
wire n_2936;
wire n_7154;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_6965;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_6647;
wire n_7279;
wire n_7499;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_7771;
wire n_2442;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_6846;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_7052;
wire n_5018;
wire n_2386;
wire n_7662;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_7728;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_6931;
wire n_4924;
wire n_2238;
wire n_6398;
wire n_6700;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_6853;
wire n_1294;
wire n_1351;
wire n_6679;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_7158;
wire n_7820;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_7299;
wire n_1830;
wire n_6770;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_7095;
wire n_7464;
wire n_1662;
wire n_7426;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_7076;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_6660;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_7666;
wire n_1962;
wire n_5296;
wire n_7246;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_7881;
wire n_7459;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_7570;
wire n_2075;
wire n_4816;
wire n_6951;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_6949;
wire n_5096;
wire n_6480;
wire n_7380;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_7809;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_7167;
wire n_7537;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_6693;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_7455;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_7755;
wire n_1726;
wire n_5751;
wire n_6819;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5862;
wire n_5869;
wire n_1238;
wire n_3959;
wire n_6937;
wire n_4288;
wire n_7629;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_7725;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_7842;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_7474;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_6860;
wire n_7739;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_6833;
wire n_2159;
wire n_6865;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_7135;
wire n_6794;
wire n_3637;
wire n_7216;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_7487;
wire n_5277;
wire n_5900;
wire n_7421;
wire n_7694;
wire n_3647;
wire n_6240;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_7399;
wire n_1956;
wire n_7186;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_7580;
wire n_7632;
wire n_6498;
wire n_6720;
wire n_1669;
wire n_7562;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_6854;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_7197;
wire n_7015;
wire n_7747;
wire n_4408;
wire n_1175;
wire n_6832;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_7066;
wire n_4341;
wire n_4759;
wire n_7688;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_6779;
wire n_2567;
wire n_5645;
wire n_7044;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_7329;
wire n_6139;
wire n_5167;
wire n_7756;
wire n_4565;
wire n_5562;
wire n_7713;
wire n_1451;
wire n_7438;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_7871;
wire n_3121;
wire n_2121;
wire n_6887;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_7735;
wire n_2278;
wire n_6769;
wire n_6903;
wire n_2433;
wire n_7255;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_6861;
wire n_2130;
wire n_4862;
wire n_7270;
wire n_5114;
wire n_7071;
wire n_7773;
wire n_6697;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_6826;
wire n_5005;
wire n_5004;
wire n_7768;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_7235;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_7129;
wire n_4242;
wire n_7243;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_7342;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_7547;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_7581;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_7310;
wire n_2911;
wire n_1828;
wire n_6972;
wire n_1389;
wire n_6380;
wire n_7200;
wire n_7751;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_6703;
wire n_7116;
wire n_4562;
wire n_1584;
wire n_7540;
wire n_7720;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6719;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_7208;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_7337;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_7055;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_7073;
wire n_2637;
wire n_7417;
wire n_7159;
wire n_5047;
wire n_5504;
wire n_7494;
wire n_7784;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_7314;
wire n_3791;
wire n_6904;
wire n_6778;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_7294;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_7016;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_6444;
wire n_7422;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_6749;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_6985;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_7891;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_7783;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_7178;
wire n_7330;
wire n_3223;
wire n_2005;
wire n_7764;
wire n_1116;
wire n_7704;
wire n_2811;
wire n_1758;
wire n_7388;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_7697;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_5308;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5982;
wire n_6692;
wire n_7079;
wire n_6590;
wire n_7536;
wire n_3036;
wire n_7209;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_7467;
wire n_4038;
wire n_5503;
wire n_7206;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_6702;
wire n_3046;
wire n_7505;
wire n_6551;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_5644;
wire n_7501;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_7490;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_7051;
wire n_7278;
wire n_2791;
wire n_1450;
wire n_7416;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_7611;
wire n_7854;
wire n_2797;
wire n_7600;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_7447;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_7520;
wire n_4442;
wire n_7702;
wire n_5700;
wire n_7274;
wire n_2168;
wire n_1442;
wire n_7668;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_6820;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_7591;
wire n_1953;
wire n_3715;
wire n_6952;
wire n_7617;
wire n_3261;
wire n_5324;
wire n_7534;
wire n_6547;
wire n_7065;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_7837;
wire n_2559;
wire n_6589;
wire n_6995;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_7461;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_7326;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_7761;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_7423;
wire n_3270;
wire n_5168;
wire n_7443;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_7746;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_7556;
wire n_1780;
wire n_1091;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_6879;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4934;
wire n_4508;
wire n_7104;
wire n_7631;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_7845;
wire n_7106;
wire n_3615;
wire n_7693;
wire n_7198;
wire n_7656;
wire n_7381;
wire n_5970;
wire n_3363;
wire n_7731;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_7182;
wire n_6310;
wire n_6852;
wire n_5061;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_6961;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_7670;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_7126;
wire n_5132;
wire n_4883;
wire n_1079;
wire n_6249;
wire n_3559;
wire n_6956;
wire n_5184;
wire n_6440;
wire n_7564;
wire n_5747;
wire n_6575;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_7524;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_6689;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_6643;
wire n_6569;
wire n_6814;
wire n_7863;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_7176;
wire n_4159;
wire n_7056;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_7594;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_7535;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_7368;
wire n_5464;
wire n_6895;
wire n_7890;
wire n_6548;
wire n_7627;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_6890;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_6789;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_6867;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_6764;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_6935;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4975;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_7382;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_7579;
wire n_3996;
wire n_7130;
wire n_6942;
wire n_6056;
wire n_7647;
wire n_2873;
wire n_1576;
wire n_6772;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_7469;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_6955;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_7654;
wire n_6375;
wire n_7762;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_7427;
wire n_6908;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_7506;
wire n_3822;
wire n_1276;
wire n_6874;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_6736;
wire n_4259;
wire n_1620;
wire n_7376;
wire n_5196;
wire n_5086;
wire n_7018;
wire n_6025;
wire n_6168;
wire n_7498;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_7134;
wire n_3967;
wire n_2373;
wire n_7456;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_7480;
wire n_7824;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_7348;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_7383;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_7053;
wire n_7660;
wire n_5483;
wire n_6713;
wire n_6919;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_7557;
wire n_3779;
wire n_3203;
wire n_7240;
wire n_7468;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_6750;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_6981;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_6675;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_7604;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_7585;
wire n_6828;
wire n_5123;
wire n_6160;
wire n_7043;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_7074;
wire n_7119;
wire n_7596;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_6875;
wire n_1701;
wire n_5236;
wire n_7567;
wire n_6678;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_7788;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_6870;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_6715;
wire n_2529;
wire n_4126;
wire n_4103;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_7386;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_7805;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_7791;
wire n_1924;
wire n_3024;
wire n_7701;
wire n_4767;
wire n_7007;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_7027;
wire n_5999;
wire n_5147;
wire n_7616;
wire n_5407;
wire n_7432;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_7661;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_7009;
wire n_6140;
wire n_5903;
wire n_7263;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_7772;
wire n_6663;
wire n_1795;
wire n_7610;
wire n_3634;
wire n_4096;
wire n_6844;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_6999;
wire n_4571;
wire n_7214;
wire n_6982;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_7613;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_6843;
wire n_3232;
wire n_7832;
wire n_5228;
wire n_7859;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_6877;
wire n_2821;
wire n_6892;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_7162;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_7510;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_7268;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_7465;
wire n_4337;
wire n_4826;
wire n_7398;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_7815;
wire n_6473;
wire n_1748;
wire n_7304;
wire n_7036;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_7462;
wire n_2490;
wire n_3127;
wire n_7171;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_7794;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_7678;
wire n_7597;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_7850;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_7293;
wire n_1264;
wire n_6752;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_7568;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_7363;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_6698;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6977;
wire n_7798;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_7511;
wire n_7028;
wire n_1628;
wire n_6810;
wire n_1773;
wire n_7237;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1115;
wire n_1395;
wire n_7039;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_6671;
wire n_6791;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_6967;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_7442;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_7618;
wire n_6768;
wire n_2458;
wire n_7489;
wire n_7144;
wire n_3032;
wire n_3401;
wire n_7362;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_6947;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6938;
wire n_7765;
wire n_6260;
wire n_5244;
wire n_7453;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_6906;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_7758;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_7124;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_6918;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_7143;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_7606;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_6834;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_6812;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_7123;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_7072;
wire n_4175;
wire n_4458;
wire n_7488;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_7827;
wire n_5776;
wire n_5826;
wire n_6687;
wire n_2684;
wire n_2205;
wire n_1104;
wire n_3284;
wire n_2875;
wire n_1437;
wire n_2747;
wire n_7848;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_7734;
wire n_6088;
wire n_6762;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_6992;
wire n_7109;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_7644;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_7325;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_7878;
wire n_1286;
wire n_6759;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_7137;
wire n_4621;
wire n_7526;
wire n_3016;
wire n_7699;
wire n_1629;
wire n_5706;
wire n_7350;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_7311;
wire n_7458;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_7244;
wire n_1524;
wire n_7681;
wire n_7882;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_7339;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_7247;
wire n_2346;
wire n_4695;
wire n_7331;
wire n_7128;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_7284;
wire n_4163;
wire n_7321;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_7309;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_7163;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_6886;
wire n_4832;
wire n_5229;
wire n_7054;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_2555;
wire n_1587;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_6959;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_7413;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_7185;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_6710;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_6945;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_6776;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_7336;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_7814;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_7630;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_6905;
wire n_7737;
wire n_7120;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_7374;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_7491;
wire n_6964;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_7001;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_7111;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_7519;
wire n_1642;
wire n_5744;
wire n_6798;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_6665;
wire n_7538;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_7165;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_6888;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_7599;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_6677;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_7389;
wire n_1501;
wire n_7418;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_7375;
wire n_7671;
wire n_7096;
wire n_5257;
wire n_7719;
wire n_7281;
wire n_7300;
wire n_4397;
wire n_6920;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_6781;
wire n_4229;
wire n_4294;
wire n_7085;
wire n_1919;
wire n_4351;
wire n_6811;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_7683;
wire n_1515;
wire n_6921;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_7212;
wire n_7285;
wire n_7676;
wire n_3871;
wire n_2388;
wire n_6685;
wire n_7590;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_7032;
wire n_7839;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_7125;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_7160;
wire n_7100;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_7319;
wire n_6162;
wire n_7638;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_7635;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_7504;
wire n_1586;
wire n_3497;
wire n_6722;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_2128;
wire n_1697;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_7767;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_7371;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_7361;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_7440;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_7010;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_7289;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_7004;
wire n_7021;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_7234;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_6975;
wire n_7266;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_7754;
wire n_6573;
wire n_6786;
wire n_6774;
wire n_6419;
wire n_7864;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_6851;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_7211;
wire n_4335;
wire n_7141;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_4471;
wire n_1141;
wire n_3297;
wire n_6729;
wire n_7150;
wire n_6882;
wire n_1168;
wire n_5500;
wire n_7378;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_7470;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_7633;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_7420;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_7558;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6189;
wire n_6167;
wire n_1074;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_6998;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_6721;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_7640;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_7484;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_7708;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_7598;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_7271;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_7322;
wire n_7549;
wire n_7022;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_6885;
wire n_7217;
wire n_7166;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_6806;
wire n_4865;
wire n_2066;
wire n_7584;
wire n_1974;
wire n_1158;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_6933;
wire n_7844;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_7811;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_7803;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_7297;
wire n_7664;
wire n_3613;
wire n_1383;
wire n_7546;
wire n_2057;
wire n_7179;
wire n_5984;
wire n_6385;
wire n_7415;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_7057;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_6793;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_6746;
wire n_4702;
wire n_1341;
wire n_7411;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_7108;
wire n_7736;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_7220;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_7223;
wire n_2544;
wire n_7261;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_7092;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_6728;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_7275;
wire n_3768;
wire n_4224;
wire n_7272;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_7436;
wire n_3181;
wire n_7249;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_7168;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_7712;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_7743;
wire n_2569;
wire n_7705;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_7091;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_6858;
wire n_7679;
wire n_1080;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_7228;
wire n_3272;
wire n_7353;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_6841;
wire n_4668;
wire n_7696;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_7687;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_6896;
wire n_1796;
wire n_3569;
wire n_2374;
wire n_1614;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_6954;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_7000;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_7876;
wire n_7040;
wire n_6132;
wire n_7196;
wire n_2799;
wire n_7655;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6872;
wire n_6089;
wire n_5211;
wire n_7205;
wire n_1668;
wire n_7260;
wire n_7500;
wire n_5861;
wire n_7086;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_7569;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_7763;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_7810;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_7577;
wire n_4874;
wire n_7836;
wire n_1228;
wire n_7047;
wire n_7412;
wire n_4840;
wire n_7717;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_7077;
wire n_2164;
wire n_7565;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6831;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_6690;
wire n_4650;
wire n_6968;
wire n_6415;
wire n_2280;
wire n_7576;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_7523;
wire n_3809;
wire n_7887;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_7750;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_7578;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_6688;
wire n_7402;
wire n_2876;
wire n_6670;
wire n_7473;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_7840;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_6680;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_7405;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_7343;
wire n_3224;
wire n_7721;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_6046;
wire n_4981;
wire n_1799;
wire n_7252;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_7817;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_6991;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_7866;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_7831;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_6705;
wire n_3567;
wire n_7601;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_7451;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_7603;
wire n_7575;
wire n_7188;
wire n_6913;
wire n_5467;
wire n_2646;
wire n_7525;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_7528;
wire n_7113;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_7637;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_6734;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_7471;
wire n_7862;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_7296;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_7781;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_7846;
wire n_4419;
wire n_2795;
wire n_7741;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_7727;
wire n_6825;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_6743;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_7345;
wire n_7472;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4542;
wire n_4122;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1985;
wire n_1140;
wire n_4740;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_7157;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_7674;
wire n_5231;
wire n_6809;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_7622;
wire n_7115;
wire n_1884;
wire n_6632;
wire n_1589;
wire n_2717;
wire n_5720;
wire n_7286;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_7865;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_6654;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_6871;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_6672;
wire n_5214;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_7344;
wire n_2006;
wire n_7714;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_7612;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_7744;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_6953;
wire n_7779;
wire n_3145;
wire n_5682;
wire n_6891;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1464;
wire n_1566;
wire n_7127;
wire n_6565;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6601;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_7873;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_6979;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_7650;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_7050;
wire n_3554;
wire n_7431;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_6930;
wire n_7829;
wire n_1935;
wire n_7770;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_7118;
wire n_7259;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_6821;
wire n_4137;
wire n_1485;
wire n_7448;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_6775;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_7518;
wire n_3797;
wire n_6683;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6815;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_7726;
wire n_4925;
wire n_2197;
wire n_7069;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_7478;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_5000;
wire n_3390;
wire n_4425;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_7011;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_7880;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5819;
wire n_5855;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_7686;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_7716;
wire n_7856;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_7759;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_7675;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_7482;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_6763;
wire n_6782;
wire n_7621;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_7552;
wire n_6839;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_7164;
wire n_6515;
wire n_6619;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_7017;
wire n_7454;
wire n_6664;
wire n_5992;
wire n_5105;
wire n_6761;
wire n_5807;
wire n_3772;
wire n_7769;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_6974;
wire n_1898;
wire n_1254;
wire n_7312;
wire n_6894;
wire n_2524;
wire n_3927;
wire n_7045;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_7277;
wire n_6099;
wire n_5939;
wire n_7502;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_6997;
wire n_3747;
wire n_1323;
wire n_6753;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_7778;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_7359;
wire n_3632;
wire n_5200;
wire n_7225;
wire n_1874;
wire n_7651;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_7020;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_7392;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2187;
wire n_2105;
wire n_5780;
wire n_2642;
wire n_6924;
wire n_5485;
wire n_5737;
wire n_6876;
wire n_7424;
wire n_1643;
wire n_1789;
wire n_7625;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_7795;
wire n_1112;
wire n_2384;
wire n_6962;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_7059;
wire n_4084;
wire n_5149;
wire n_3174;
wire n_1527;
wire n_4848;
wire n_6970;
wire n_5185;
wire n_6829;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_7522;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_6830;
wire n_3290;
wire n_7365;
wire n_3585;
wire n_7094;
wire n_2878;
wire n_1810;
wire n_7439;
wire n_7872;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_7035;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_6838;
wire n_2698;
wire n_6869;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_6735;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_6866;
wire n_4383;
wire n_7395;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_7005;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_6742;
wire n_3063;
wire n_4543;
wire n_6969;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_7180;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_6929;
wire n_2255;
wire n_1820;
wire n_6986;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_7752;
wire n_6709;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_7724;
wire n_4068;
wire n_7385;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_7444;
wire n_6756;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_7620;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_7441;
wire n_6250;
wire n_6718;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_7078;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_7093;
wire n_1167;
wire n_7333;
wire n_3231;
wire n_6423;
wire n_6659;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_7508;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6668;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_6757;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_7496;
wire n_3649;
wire n_1838;
wire n_6880;
wire n_3824;
wire n_7425;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_7550;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_7715;
wire n_5768;
wire n_6353;
wire n_7302;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_7548;
wire n_5142;
wire n_1433;
wire n_6934;
wire n_5082;
wire n_1907;
wire n_6686;
wire n_7019;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_7595;
wire n_1088;
wire n_7088;
wire n_6666;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_7542;
wire n_4487;
wire n_7204;
wire n_7014;
wire n_1165;
wire n_6708;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_7665;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_7341;
wire n_7407;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_7757;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_7514;
wire n_6317;
wire n_7646;
wire n_7653;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_6801;
wire n_1542;
wire n_1547;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_7193;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_7373;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_7291;
wire n_2593;
wire n_7818;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_1131;
wire n_6707;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_7239;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_6835;
wire n_7406;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_6792;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_7677;
wire n_7799;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_7513;
wire n_2207;
wire n_4210;
wire n_7782;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_6928;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_7861;
wire n_4461;
wire n_2323;
wire n_7242;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_7573;
wire n_5112;
wire n_3042;
wire n_5627;
wire n_5542;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_7181;
wire n_1161;
wire n_1103;
wire n_6739;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_7139;
wire n_6194;
wire n_1911;
wire n_7586;
wire n_6381;
wire n_7404;
wire n_2870;
wire n_6862;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_7328;
wire n_6783;
wire n_4738;
wire n_7231;
wire n_6604;
wire n_1193;
wire n_2928;
wire n_3557;
wire n_3380;
wire n_7435;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_7058;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_7041;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_6788;
wire n_2668;
wire n_6684;
wire n_1386;
wire n_2931;
wire n_7364;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_7738;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_7869;
wire n_7825;
wire n_3938;
wire n_6103;
wire n_7006;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_6817;
wire n_1661;
wire n_6261;
wire n_7276;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_7571;
wire n_7269;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_6845;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_6572;
wire n_4544;
wire n_7531;
wire n_7222;
wire n_4418;
wire n_4595;
wire n_7867;
wire n_2770;
wire n_7463;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_7347;
wire n_4944;
wire n_7060;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_7064;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_6917;
wire n_7545;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_7479;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_7400;
wire n_4194;
wire n_7808;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_6813;
wire n_2670;
wire n_7379;
wire n_1745;
wire n_7318;
wire n_7352;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_7295;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_7785;
wire n_7267;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_7497;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_1113;
wire n_6963;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_7543;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_6923;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_7870;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_6681;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_7460;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_7061;
wire n_7351;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_7298;
wire n_2497;
wire n_7195;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_6957;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_822),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_894),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_826),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_165),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_407),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_762),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_958),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_697),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_789),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1039),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_114),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_1036),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_360),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_1008),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_947),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_153),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_967),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_345),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_749),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_873),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_824),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_993),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_413),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_366),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_954),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_888),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_17),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_144),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_15),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_62),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_992),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_321),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_477),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_758),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_120),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_749),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_25),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_376),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_905),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_973),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_272),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_408),
.Y(n_1113)
);

BUFx10_ASAP7_75t_L g1114 ( 
.A(n_476),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_366),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_629),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_552),
.Y(n_1117)
);

BUFx10_ASAP7_75t_L g1118 ( 
.A(n_471),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_620),
.Y(n_1119)
);

CKINVDCx16_ASAP7_75t_R g1120 ( 
.A(n_52),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_839),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_760),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_27),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_169),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_1060),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_208),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_318),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_970),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_249),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_249),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_984),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_751),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_399),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_279),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_957),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_656),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_942),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_975),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_908),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_891),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_339),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1021),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_252),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_697),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_331),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_908),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1004),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_998),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_183),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1005),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_128),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_955),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_446),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_459),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_568),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_3),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_964),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_311),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_974),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_823),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_253),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_522),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_165),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_728),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_339),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_614),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_212),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_490),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_543),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1034),
.Y(n_1170)
);

CKINVDCx16_ASAP7_75t_R g1171 ( 
.A(n_640),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_520),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_945),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_744),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_976),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1060),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_706),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_988),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_75),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_57),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_748),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_791),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1013),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_718),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_265),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_417),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_979),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_900),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_233),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_965),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_694),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_977),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_776),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_855),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1016),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_753),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1038),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_176),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_700),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_702),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_125),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_110),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_757),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_686),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1038),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_242),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_590),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_624),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_847),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_135),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_951),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1014),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_419),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_455),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_144),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1057),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_85),
.Y(n_1217)
);

BUFx5_ASAP7_75t_L g1218 ( 
.A(n_630),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_869),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_874),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_265),
.Y(n_1221)
);

BUFx10_ASAP7_75t_L g1222 ( 
.A(n_667),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_682),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_943),
.Y(n_1224)
);

CKINVDCx20_ASAP7_75t_R g1225 ( 
.A(n_919),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_910),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_57),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_938),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1029),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_945),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_861),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_456),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_668),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1033),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_812),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_944),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_424),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1015),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_821),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_161),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_947),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_796),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_578),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1064),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_727),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_982),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_193),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_140),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_660),
.Y(n_1249)
);

CKINVDCx16_ASAP7_75t_R g1250 ( 
.A(n_959),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_969),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_954),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_959),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_429),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_33),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_57),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_937),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_797),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_226),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1031),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_189),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_325),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1013),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_929),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_115),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_390),
.Y(n_1266)
);

BUFx2_ASAP7_75t_SL g1267 ( 
.A(n_201),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_940),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_408),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_650),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_277),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_882),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_407),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_911),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1026),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_322),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_977),
.Y(n_1277)
);

BUFx2_ASAP7_75t_SL g1278 ( 
.A(n_598),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_473),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_150),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1020),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1032),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_948),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_910),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_149),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_914),
.Y(n_1286)
);

CKINVDCx20_ASAP7_75t_R g1287 ( 
.A(n_1030),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_873),
.Y(n_1288)
);

BUFx5_ASAP7_75t_L g1289 ( 
.A(n_460),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_48),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_728),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_853),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_402),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1012),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1001),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_900),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_154),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_576),
.Y(n_1298)
);

CKINVDCx14_ASAP7_75t_R g1299 ( 
.A(n_935),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_467),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1051),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_241),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1023),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_868),
.Y(n_1304)
);

BUFx10_ASAP7_75t_L g1305 ( 
.A(n_856),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_614),
.Y(n_1306)
);

INVxp67_ASAP7_75t_SL g1307 ( 
.A(n_281),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1002),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_780),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_500),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1067),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_817),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_336),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_989),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_747),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_62),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_962),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1045),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_752),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_455),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1045),
.Y(n_1321)
);

BUFx2_ASAP7_75t_SL g1322 ( 
.A(n_1043),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_136),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_178),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_633),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_433),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_526),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_868),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_225),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_569),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_934),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_384),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1025),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_381),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_992),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_8),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_198),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_990),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_158),
.Y(n_1339)
);

CKINVDCx16_ASAP7_75t_R g1340 ( 
.A(n_15),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_82),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_968),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_20),
.Y(n_1343)
);

BUFx10_ASAP7_75t_L g1344 ( 
.A(n_352),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_954),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_99),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1024),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_189),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_971),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_401),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_448),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_326),
.Y(n_1352)
);

BUFx2_ASAP7_75t_SL g1353 ( 
.A(n_361),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1057),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_402),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_840),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_125),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_961),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_66),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_704),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_350),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_193),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_331),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_866),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1000),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1063),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_978),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_635),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_564),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_381),
.Y(n_1370)
);

CKINVDCx14_ASAP7_75t_R g1371 ( 
.A(n_138),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_561),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_519),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1006),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_757),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1022),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_991),
.Y(n_1377)
);

INVxp33_ASAP7_75t_SL g1378 ( 
.A(n_634),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_7),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_85),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_369),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_15),
.Y(n_1382)
);

CKINVDCx16_ASAP7_75t_R g1383 ( 
.A(n_54),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_676),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_41),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_635),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_600),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_580),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_0),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_475),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_127),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_559),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_425),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_981),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_946),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_410),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_425),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_972),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_404),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_690),
.Y(n_1400)
);

BUFx10_ASAP7_75t_L g1401 ( 
.A(n_1003),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_546),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1031),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_438),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_141),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_213),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_748),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_436),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1062),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_576),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1065),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_641),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_4),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_492),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_795),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_199),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_72),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_232),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_794),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_408),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_673),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_587),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_876),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_714),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_64),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_779),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_227),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_535),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_180),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1051),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_531),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_993),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1024),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_326),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1035),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_941),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_780),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_777),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_406),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_154),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_739),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_597),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_144),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1009),
.Y(n_1444)
);

BUFx10_ASAP7_75t_L g1445 ( 
.A(n_554),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_136),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1055),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1066),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_730),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_43),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_124),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_999),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_473),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_234),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_995),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_207),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1032),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_339),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_222),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_997),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_889),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_637),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_306),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_443),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_682),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_983),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_360),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1051),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_53),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_673),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_695),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_260),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_840),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_447),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_951),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_113),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_612),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_773),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_395),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_572),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_684),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1027),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_41),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_582),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_186),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_995),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_428),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_6),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1044),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_197),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_653),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_501),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_212),
.Y(n_1493)
);

BUFx8_ASAP7_75t_SL g1494 ( 
.A(n_23),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1044),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_700),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_607),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_245),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_960),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_45),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_870),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_709),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_224),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_840),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1052),
.Y(n_1505)
);

BUFx10_ASAP7_75t_L g1506 ( 
.A(n_33),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_894),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_291),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_981),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_558),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_902),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_457),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_750),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1044),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_952),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_896),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_713),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_605),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_536),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_131),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_435),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_404),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_996),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_189),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_134),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_163),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_583),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_704),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_804),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_949),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_98),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_68),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_264),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_589),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_26),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_620),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_829),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_482),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_641),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_644),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_79),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_583),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1037),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_793),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1041),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_426),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_472),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_232),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_950),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_30),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_790),
.Y(n_1551)
);

BUFx8_ASAP7_75t_SL g1552 ( 
.A(n_21),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_771),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_344),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_333),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_646),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1028),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_523),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_984),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1007),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_788),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_37),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_191),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1005),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_222),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_494),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_851),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_764),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1029),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_680),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_581),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1019),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1016),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_661),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_623),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1018),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_377),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_582),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_963),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1004),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_576),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_748),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1010),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_983),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_885),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_935),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1030),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_292),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_793),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_669),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_418),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1028),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_126),
.Y(n_1593)
);

BUFx2_ASAP7_75t_SL g1594 ( 
.A(n_77),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_274),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_648),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_985),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1006),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_709),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_62),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1042),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1016),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_319),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_483),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_776),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_158),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_565),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_326),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_809),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_816),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_278),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_275),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_896),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_343),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_665),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_314),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_476),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_613),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_698),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_734),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_703),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_74),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_987),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_572),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_86),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_447),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_785),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_260),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_92),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_684),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1029),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1024),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_742),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_277),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_676),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_980),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_424),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_504),
.Y(n_1638)
);

BUFx10_ASAP7_75t_L g1639 ( 
.A(n_184),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_222),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_892),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_397),
.Y(n_1642)
);

CKINVDCx16_ASAP7_75t_R g1643 ( 
.A(n_837),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1045),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_441),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_904),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_492),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_325),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_607),
.Y(n_1649)
);

INVxp67_ASAP7_75t_SL g1650 ( 
.A(n_854),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1062),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_953),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_504),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_452),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_448),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_206),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_259),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_119),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_26),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_236),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_717),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_994),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_588),
.Y(n_1663)
);

BUFx10_ASAP7_75t_L g1664 ( 
.A(n_415),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_86),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_548),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_224),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_890),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1010),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_774),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_966),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_433),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_460),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_29),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_23),
.Y(n_1675)
);

BUFx10_ASAP7_75t_L g1676 ( 
.A(n_113),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_918),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_25),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_985),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1018),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_971),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_939),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_320),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_43),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_352),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_354),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_75),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_405),
.Y(n_1688)
);

CKINVDCx16_ASAP7_75t_R g1689 ( 
.A(n_1007),
.Y(n_1689)
);

CKINVDCx14_ASAP7_75t_R g1690 ( 
.A(n_302),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_151),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_934),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_502),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_222),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_97),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_899),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_956),
.Y(n_1697)
);

BUFx10_ASAP7_75t_L g1698 ( 
.A(n_1041),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_189),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_728),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1011),
.Y(n_1701)
);

CKINVDCx20_ASAP7_75t_R g1702 ( 
.A(n_1040),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_24),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_986),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_679),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1017),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_936),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_922),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_232),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1037),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_410),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_486),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_688),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1102),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1218),
.Y(n_1715)
);

INVxp33_ASAP7_75t_L g1716 ( 
.A(n_1494),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1506),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1218),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1102),
.Y(n_1719)
);

CKINVDCx14_ASAP7_75t_R g1720 ( 
.A(n_1371),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1494),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1552),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1552),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1506),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1218),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1506),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1676),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1676),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1130),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1676),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1639),
.Y(n_1731)
);

CKINVDCx16_ASAP7_75t_R g1732 ( 
.A(n_1120),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1206),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1218),
.Y(n_1734)
);

CKINVDCx20_ASAP7_75t_R g1735 ( 
.A(n_1341),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1297),
.Y(n_1736)
);

CKINVDCx20_ASAP7_75t_R g1737 ( 
.A(n_1341),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1340),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1639),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1218),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1639),
.Y(n_1741)
);

CKINVDCx20_ASAP7_75t_R g1742 ( 
.A(n_1380),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1490),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1218),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1206),
.Y(n_1745)
);

BUFx6f_ASAP7_75t_L g1746 ( 
.A(n_1102),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1186),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1383),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1218),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1206),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1075),
.Y(n_1751)
);

INVxp33_ASAP7_75t_SL g1752 ( 
.A(n_1292),
.Y(n_1752)
);

CKINVDCx16_ASAP7_75t_R g1753 ( 
.A(n_1133),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1130),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1143),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1289),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1143),
.Y(n_1757)
);

NOR2xp67_ASAP7_75t_L g1758 ( 
.A(n_1216),
.B(n_0),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1100),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1106),
.Y(n_1760)
);

CKINVDCx14_ASAP7_75t_R g1761 ( 
.A(n_1299),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1126),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1129),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1198),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1709),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1215),
.Y(n_1766)
);

INVxp67_ASAP7_75t_SL g1767 ( 
.A(n_1189),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1709),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1217),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1227),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1261),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1265),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1690),
.Y(n_1773)
);

INVxp67_ASAP7_75t_SL g1774 ( 
.A(n_1189),
.Y(n_1774)
);

INVxp67_ASAP7_75t_SL g1775 ( 
.A(n_1357),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1389),
.Y(n_1776)
);

CKINVDCx16_ASAP7_75t_R g1777 ( 
.A(n_1171),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1289),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1391),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1082),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1413),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1289),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1087),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1454),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1380),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1476),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1483),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1498),
.Y(n_1788)
);

CKINVDCx16_ASAP7_75t_R g1789 ( 
.A(n_1200),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1524),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1525),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1316),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1099),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1101),
.Y(n_1794)
);

CKINVDCx20_ASAP7_75t_R g1795 ( 
.A(n_1687),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1699),
.Y(n_1796)
);

CKINVDCx20_ASAP7_75t_R g1797 ( 
.A(n_1687),
.Y(n_1797)
);

CKINVDCx20_ASAP7_75t_R g1798 ( 
.A(n_1076),
.Y(n_1798)
);

CKINVDCx16_ASAP7_75t_R g1799 ( 
.A(n_1250),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1108),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1123),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1703),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1533),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1124),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1535),
.Y(n_1805)
);

CKINVDCx20_ASAP7_75t_R g1806 ( 
.A(n_1076),
.Y(n_1806)
);

CKINVDCx20_ASAP7_75t_R g1807 ( 
.A(n_1090),
.Y(n_1807)
);

INVx1_ASAP7_75t_SL g1808 ( 
.A(n_1606),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1541),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1102),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1548),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1149),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1565),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1656),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1660),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1448),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1151),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1675),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1678),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1691),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1695),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1216),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1216),
.Y(n_1823)
);

INVxp33_ASAP7_75t_SL g1824 ( 
.A(n_1309),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1156),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1470),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1161),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1167),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1420),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1179),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1420),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1180),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1328),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1420),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1473),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1473),
.Y(n_1836)
);

CKINVDCx20_ASAP7_75t_R g1837 ( 
.A(n_1090),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_1107),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1201),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1202),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1107),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1473),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1662),
.Y(n_1843)
);

BUFx5_ASAP7_75t_L g1844 ( 
.A(n_1357),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1590),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1666),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1103),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1289),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1103),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1257),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1257),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1754),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1745),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1755),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1733),
.Y(n_1855)
);

CKINVDCx20_ASAP7_75t_R g1856 ( 
.A(n_1735),
.Y(n_1856)
);

INVxp33_ASAP7_75t_SL g1857 ( 
.A(n_1792),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1802),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_1737),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1808),
.Y(n_1860)
);

CKINVDCx20_ASAP7_75t_R g1861 ( 
.A(n_1742),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1767),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1757),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1729),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1765),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1768),
.Y(n_1866)
);

CKINVDCx20_ASAP7_75t_R g1867 ( 
.A(n_1785),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1780),
.Y(n_1868)
);

BUFx2_ASAP7_75t_SL g1869 ( 
.A(n_1833),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1783),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1774),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1795),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1775),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1847),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1849),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1750),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_1797),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1822),
.Y(n_1878)
);

INVxp67_ASAP7_75t_SL g1879 ( 
.A(n_1736),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1793),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1794),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1796),
.Y(n_1882)
);

INVxp33_ASAP7_75t_L g1883 ( 
.A(n_1816),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1800),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1823),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1829),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1831),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1834),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1801),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1835),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1836),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1717),
.B(n_1378),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1732),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1804),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1842),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1751),
.Y(n_1896)
);

CKINVDCx20_ASAP7_75t_R g1897 ( 
.A(n_1798),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1759),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1760),
.Y(n_1899)
);

INVxp67_ASAP7_75t_SL g1900 ( 
.A(n_1747),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1844),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1762),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1763),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_1806),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1812),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1817),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1764),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1766),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1769),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1770),
.Y(n_1910)
);

INVxp67_ASAP7_75t_SL g1911 ( 
.A(n_1771),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1772),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1776),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1825),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1844),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1844),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1827),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1807),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1779),
.Y(n_1919)
);

INVxp67_ASAP7_75t_SL g1920 ( 
.A(n_1781),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1837),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1828),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1743),
.B(n_1210),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1784),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1786),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1787),
.Y(n_1926)
);

INVxp33_ASAP7_75t_SL g1927 ( 
.A(n_1830),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1788),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1790),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1826),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1791),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1803),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1832),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1805),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1809),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1839),
.Y(n_1936)
);

CKINVDCx20_ASAP7_75t_R g1937 ( 
.A(n_1838),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1811),
.Y(n_1938)
);

CKINVDCx20_ASAP7_75t_R g1939 ( 
.A(n_1841),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1813),
.Y(n_1940)
);

CKINVDCx16_ASAP7_75t_R g1941 ( 
.A(n_1753),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1840),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1720),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1722),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1814),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1815),
.Y(n_1946)
);

CKINVDCx20_ASAP7_75t_R g1947 ( 
.A(n_1777),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1818),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1819),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1723),
.Y(n_1950)
);

CKINVDCx20_ASAP7_75t_R g1951 ( 
.A(n_1789),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1820),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1721),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1738),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1821),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1748),
.Y(n_1956)
);

INVxp67_ASAP7_75t_SL g1957 ( 
.A(n_1752),
.Y(n_1957)
);

CKINVDCx20_ASAP7_75t_R g1958 ( 
.A(n_1799),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1758),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1761),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1724),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1726),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1824),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1773),
.Y(n_1964)
);

BUFx2_ASAP7_75t_L g1965 ( 
.A(n_1845),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1727),
.B(n_1240),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1728),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1730),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1846),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1843),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1731),
.Y(n_1971)
);

CKINVDCx20_ASAP7_75t_R g1972 ( 
.A(n_1739),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1741),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1716),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1844),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1844),
.Y(n_1976)
);

CKINVDCx16_ASAP7_75t_R g1977 ( 
.A(n_1715),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1718),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1725),
.B(n_1378),
.Y(n_1979)
);

INVxp67_ASAP7_75t_L g1980 ( 
.A(n_1734),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1740),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1744),
.B(n_1247),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1749),
.B(n_1643),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1756),
.Y(n_1984)
);

CKINVDCx16_ASAP7_75t_R g1985 ( 
.A(n_1778),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1782),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1848),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1714),
.Y(n_1988)
);

INVxp67_ASAP7_75t_L g1989 ( 
.A(n_1714),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1714),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1719),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1719),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1851),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1719),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1746),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1746),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1746),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1851),
.B(n_1689),
.Y(n_1998)
);

CKINVDCx20_ASAP7_75t_R g1999 ( 
.A(n_1851),
.Y(n_1999)
);

BUFx2_ASAP7_75t_L g2000 ( 
.A(n_1810),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1810),
.Y(n_2001)
);

CKINVDCx20_ASAP7_75t_R g2002 ( 
.A(n_1810),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1850),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1850),
.Y(n_2004)
);

CKINVDCx20_ASAP7_75t_R g2005 ( 
.A(n_1850),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1735),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1745),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_1754),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1745),
.Y(n_2009)
);

CKINVDCx20_ASAP7_75t_R g2010 ( 
.A(n_1735),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1745),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1745),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1816),
.B(n_1267),
.Y(n_2013)
);

CKINVDCx20_ASAP7_75t_R g2014 ( 
.A(n_1735),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1754),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1717),
.B(n_1429),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1745),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1754),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1745),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1745),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1754),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1792),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1717),
.B(n_1144),
.Y(n_2023)
);

CKINVDCx20_ASAP7_75t_R g2024 ( 
.A(n_1735),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1754),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1745),
.Y(n_2026)
);

CKINVDCx20_ASAP7_75t_R g2027 ( 
.A(n_1735),
.Y(n_2027)
);

CKINVDCx20_ASAP7_75t_R g2028 ( 
.A(n_1735),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1745),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1745),
.Y(n_2030)
);

INVxp67_ASAP7_75t_SL g2031 ( 
.A(n_1792),
.Y(n_2031)
);

CKINVDCx20_ASAP7_75t_R g2032 ( 
.A(n_1735),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1754),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1754),
.Y(n_2034)
);

CKINVDCx20_ASAP7_75t_R g2035 ( 
.A(n_1735),
.Y(n_2035)
);

INVxp33_ASAP7_75t_SL g2036 ( 
.A(n_1792),
.Y(n_2036)
);

HB1xp67_ASAP7_75t_L g2037 ( 
.A(n_1792),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1754),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1802),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1745),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1754),
.Y(n_2041)
);

INVxp67_ASAP7_75t_SL g2042 ( 
.A(n_1792),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1745),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_1754),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1745),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1745),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1745),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1754),
.Y(n_2048)
);

CKINVDCx20_ASAP7_75t_R g2049 ( 
.A(n_1735),
.Y(n_2049)
);

CKINVDCx20_ASAP7_75t_R g2050 ( 
.A(n_1735),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1745),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1745),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1754),
.Y(n_2053)
);

CKINVDCx20_ASAP7_75t_R g2054 ( 
.A(n_1735),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1754),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1745),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1717),
.B(n_1207),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1754),
.Y(n_2058)
);

CKINVDCx20_ASAP7_75t_R g2059 ( 
.A(n_1735),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_R g2060 ( 
.A(n_1720),
.B(n_1248),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_1792),
.Y(n_2061)
);

CKINVDCx20_ASAP7_75t_R g2062 ( 
.A(n_1735),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1754),
.Y(n_2063)
);

CKINVDCx16_ASAP7_75t_R g2064 ( 
.A(n_1732),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1745),
.Y(n_2065)
);

CKINVDCx20_ASAP7_75t_R g2066 ( 
.A(n_1735),
.Y(n_2066)
);

CKINVDCx20_ASAP7_75t_R g2067 ( 
.A(n_1735),
.Y(n_2067)
);

CKINVDCx20_ASAP7_75t_R g2068 ( 
.A(n_1735),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1802),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1754),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1745),
.Y(n_2071)
);

BUFx2_ASAP7_75t_SL g2072 ( 
.A(n_1792),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1792),
.Y(n_2073)
);

HB1xp67_ASAP7_75t_L g2074 ( 
.A(n_1792),
.Y(n_2074)
);

CKINVDCx20_ASAP7_75t_R g2075 ( 
.A(n_1735),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1745),
.Y(n_2076)
);

INVxp67_ASAP7_75t_SL g2077 ( 
.A(n_1792),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1745),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1802),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1745),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_1735),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1745),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_1977),
.Y(n_2083)
);

INVx1_ASAP7_75t_SL g2084 ( 
.A(n_2072),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1874),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2039),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1911),
.B(n_1255),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1875),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2069),
.Y(n_2089)
);

BUFx8_ASAP7_75t_L g2090 ( 
.A(n_1880),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1920),
.Y(n_2091)
);

AND2x6_ASAP7_75t_L g2092 ( 
.A(n_1855),
.B(n_1417),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2079),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1983),
.B(n_1256),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2037),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2037),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2061),
.Y(n_2097)
);

OAI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_1860),
.A2(n_1280),
.B1(n_1285),
.B2(n_1259),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2000),
.Y(n_2099)
);

OAI21x1_ASAP7_75t_L g2100 ( 
.A1(n_1982),
.A2(n_1324),
.B(n_1098),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2061),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1878),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_2022),
.B(n_1072),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_2013),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1885),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1995),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1868),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1886),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1995),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1887),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1876),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_2073),
.B(n_1072),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_1973),
.B(n_1519),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_2073),
.B(n_1128),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2074),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_1985),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2074),
.B(n_1128),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1857),
.B(n_1302),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1858),
.Y(n_2119)
);

HB1xp67_ASAP7_75t_L g2120 ( 
.A(n_2036),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1966),
.B(n_1323),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1961),
.Y(n_2122)
);

AOI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_1969),
.A2(n_1892),
.B1(n_1879),
.B2(n_2031),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1962),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1870),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1869),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1888),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1967),
.B(n_1968),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_L g2129 ( 
.A(n_1881),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_2042),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1890),
.Y(n_2131)
);

INVxp33_ASAP7_75t_L g2132 ( 
.A(n_1963),
.Y(n_2132)
);

BUFx2_ASAP7_75t_L g2133 ( 
.A(n_2077),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1971),
.B(n_1329),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1891),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1895),
.Y(n_2136)
);

AND2x4_ASAP7_75t_L g2137 ( 
.A(n_1864),
.B(n_1131),
.Y(n_2137)
);

OR2x6_ASAP7_75t_L g2138 ( 
.A(n_1963),
.B(n_1278),
.Y(n_2138)
);

OAI22xp5_ASAP7_75t_SL g2139 ( 
.A1(n_1856),
.A2(n_1125),
.B1(n_1134),
.B2(n_1109),
.Y(n_2139)
);

INVx4_ASAP7_75t_L g2140 ( 
.A(n_1882),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1884),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1853),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2007),
.Y(n_2143)
);

BUFx6f_ASAP7_75t_L g2144 ( 
.A(n_1889),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1973),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_1894),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1862),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1871),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2009),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1873),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_1864),
.B(n_1131),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1970),
.A2(n_1337),
.B1(n_1343),
.B2(n_1336),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1883),
.B(n_1135),
.Y(n_2153)
);

BUFx6f_ASAP7_75t_L g2154 ( 
.A(n_1905),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2011),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_1906),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1959),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2012),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_1900),
.A2(n_1348),
.B1(n_1359),
.B2(n_1346),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_2064),
.Y(n_2160)
);

NOR2x1_ASAP7_75t_L g2161 ( 
.A(n_1923),
.B(n_1160),
.Y(n_2161)
);

OA21x2_ASAP7_75t_L g2162 ( 
.A1(n_1975),
.A2(n_1324),
.B(n_1098),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1896),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_1965),
.A2(n_1382),
.B1(n_1385),
.B2(n_1362),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_1914),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1898),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1899),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2017),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1917),
.Y(n_2169)
);

INVx4_ASAP7_75t_L g2170 ( 
.A(n_1922),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2016),
.B(n_1405),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_1927),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2019),
.Y(n_2173)
);

OAI22xp33_ASAP7_75t_R g2174 ( 
.A1(n_1957),
.A2(n_1650),
.B1(n_1307),
.B2(n_1086),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_L g2175 ( 
.A(n_1936),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1902),
.Y(n_2176)
);

AND2x4_ASAP7_75t_L g2177 ( 
.A(n_1943),
.B(n_1933),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1930),
.B(n_1135),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2016),
.B(n_1406),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2020),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1903),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2026),
.Y(n_2182)
);

OAI22xp5_ASAP7_75t_SL g2183 ( 
.A1(n_1859),
.A2(n_1867),
.B1(n_1872),
.B2(n_1861),
.Y(n_2183)
);

BUFx8_ASAP7_75t_L g2184 ( 
.A(n_1941),
.Y(n_2184)
);

BUFx6f_ASAP7_75t_L g2185 ( 
.A(n_1990),
.Y(n_2185)
);

BUFx6f_ASAP7_75t_L g2186 ( 
.A(n_1992),
.Y(n_2186)
);

OA21x2_ASAP7_75t_L g2187 ( 
.A1(n_1901),
.A2(n_1443),
.B(n_1379),
.Y(n_2187)
);

NOR2x1_ASAP7_75t_L g2188 ( 
.A(n_2023),
.B(n_2057),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2029),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1907),
.Y(n_2190)
);

INVx3_ASAP7_75t_L g2191 ( 
.A(n_2030),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1877),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2040),
.Y(n_2193)
);

NOR2x1_ASAP7_75t_L g2194 ( 
.A(n_2023),
.B(n_1972),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1908),
.B(n_1416),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1996),
.Y(n_2196)
);

BUFx6f_ASAP7_75t_L g2197 ( 
.A(n_2001),
.Y(n_2197)
);

AND2x6_ASAP7_75t_L g2198 ( 
.A(n_1979),
.B(n_1417),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1909),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1910),
.Y(n_2200)
);

INVx3_ASAP7_75t_L g2201 ( 
.A(n_2043),
.Y(n_2201)
);

INVx3_ASAP7_75t_L g2202 ( 
.A(n_2045),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1912),
.Y(n_2203)
);

OAI22x1_ASAP7_75t_R g2204 ( 
.A1(n_2006),
.A2(n_1125),
.B1(n_1134),
.B2(n_1109),
.Y(n_2204)
);

BUFx12f_ASAP7_75t_L g2205 ( 
.A(n_1960),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1933),
.B(n_1139),
.Y(n_2206)
);

OAI22xp5_ASAP7_75t_SL g2207 ( 
.A1(n_2010),
.A2(n_1175),
.B1(n_1195),
.B2(n_1172),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1913),
.Y(n_2208)
);

OAI22xp5_ASAP7_75t_SL g2209 ( 
.A1(n_2014),
.A2(n_1175),
.B1(n_1195),
.B2(n_1172),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1919),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2046),
.Y(n_2211)
);

INVxp33_ASAP7_75t_SL g2212 ( 
.A(n_2060),
.Y(n_2212)
);

INVx6_ASAP7_75t_L g2213 ( 
.A(n_1999),
.Y(n_2213)
);

CKINVDCx6p67_ASAP7_75t_R g2214 ( 
.A(n_1893),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_1943),
.B(n_1139),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1924),
.Y(n_2216)
);

BUFx6f_ASAP7_75t_L g2217 ( 
.A(n_2004),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2047),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1925),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2051),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1926),
.B(n_1418),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2052),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2056),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2065),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_1942),
.B(n_1140),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1928),
.Y(n_2226)
);

XNOR2x2_ASAP7_75t_L g2227 ( 
.A(n_1998),
.B(n_1094),
.Y(n_2227)
);

INVx5_ASAP7_75t_L g2228 ( 
.A(n_1915),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_1929),
.B(n_1620),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2071),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1931),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_1852),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_1942),
.B(n_1140),
.Y(n_2233)
);

OAI22xp33_ASAP7_75t_R g2234 ( 
.A1(n_2024),
.A2(n_2028),
.B1(n_2032),
.B2(n_2027),
.Y(n_2234)
);

AND2x6_ASAP7_75t_L g2235 ( 
.A(n_1932),
.B(n_1450),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2076),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_1934),
.B(n_1425),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1935),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_1974),
.B(n_1141),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1938),
.Y(n_2240)
);

HB1xp67_ASAP7_75t_L g2241 ( 
.A(n_1854),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1940),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_2078),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1945),
.B(n_1427),
.Y(n_2244)
);

BUFx2_ASAP7_75t_L g2245 ( 
.A(n_1863),
.Y(n_2245)
);

AND2x6_ASAP7_75t_L g2246 ( 
.A(n_1946),
.B(n_1450),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1865),
.Y(n_2247)
);

OA21x2_ASAP7_75t_L g2248 ( 
.A1(n_1916),
.A2(n_1443),
.B(n_1379),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_2035),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_1866),
.B(n_1141),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1948),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1949),
.Y(n_2252)
);

INVx3_ASAP7_75t_L g2253 ( 
.A(n_2080),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_2008),
.Y(n_2254)
);

BUFx6f_ASAP7_75t_L g2255 ( 
.A(n_2015),
.Y(n_2255)
);

INVx3_ASAP7_75t_L g2256 ( 
.A(n_2082),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1952),
.Y(n_2257)
);

HB1xp67_ASAP7_75t_L g2258 ( 
.A(n_2018),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1955),
.B(n_1446),
.Y(n_2259)
);

BUFx2_ASAP7_75t_L g2260 ( 
.A(n_2021),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1987),
.B(n_1980),
.Y(n_2261)
);

OA21x2_ASAP7_75t_L g2262 ( 
.A1(n_1978),
.A2(n_1562),
.B(n_1493),
.Y(n_2262)
);

AND2x6_ASAP7_75t_L g2263 ( 
.A(n_1981),
.B(n_1674),
.Y(n_2263)
);

NOR2x1_ASAP7_75t_L g2264 ( 
.A(n_2002),
.B(n_1160),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1984),
.Y(n_2265)
);

INVxp67_ASAP7_75t_L g2266 ( 
.A(n_2025),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1986),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_2033),
.B(n_1142),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2034),
.B(n_1451),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_2038),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1976),
.B(n_1456),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1989),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2005),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1993),
.Y(n_2274)
);

BUFx3_ASAP7_75t_L g2275 ( 
.A(n_1954),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_2041),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2044),
.Y(n_2277)
);

NAND2xp33_ASAP7_75t_L g2278 ( 
.A(n_2048),
.B(n_1289),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2053),
.Y(n_2279)
);

AND2x2_ASAP7_75t_SL g2280 ( 
.A(n_1947),
.B(n_1081),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2055),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_2049),
.Y(n_2282)
);

BUFx12f_ASAP7_75t_L g2283 ( 
.A(n_1956),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2058),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_L g2285 ( 
.A(n_2063),
.B(n_1459),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2070),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1964),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1944),
.B(n_1469),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1988),
.Y(n_2289)
);

BUFx12f_ASAP7_75t_L g2290 ( 
.A(n_1950),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1991),
.Y(n_2291)
);

BUFx6f_ASAP7_75t_L g2292 ( 
.A(n_1994),
.Y(n_2292)
);

AND2x6_ASAP7_75t_L g2293 ( 
.A(n_1997),
.B(n_1674),
.Y(n_2293)
);

BUFx12f_ASAP7_75t_L g2294 ( 
.A(n_1953),
.Y(n_2294)
);

BUFx12f_ASAP7_75t_L g2295 ( 
.A(n_1951),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2003),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1958),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2050),
.B(n_1472),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_SL g2299 ( 
.A(n_2054),
.B(n_1142),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2059),
.Y(n_2300)
);

INVx6_ASAP7_75t_L g2301 ( 
.A(n_2062),
.Y(n_2301)
);

AND2x2_ASAP7_75t_SL g2302 ( 
.A(n_2066),
.B(n_1081),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2067),
.B(n_1485),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_2081),
.B(n_1488),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2068),
.B(n_1393),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2075),
.B(n_1393),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_1897),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1904),
.Y(n_2308)
);

OAI22xp5_ASAP7_75t_SL g2309 ( 
.A1(n_1918),
.A2(n_1220),
.B1(n_1225),
.B2(n_1209),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1939),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_1921),
.B(n_1704),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_1937),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1874),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1880),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2039),
.Y(n_2315)
);

BUFx3_ASAP7_75t_L g2316 ( 
.A(n_1857),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2039),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1874),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1874),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1874),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1911),
.B(n_1500),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_1880),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2039),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_1911),
.B(n_1503),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1911),
.B(n_1520),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_1860),
.B(n_1704),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1874),
.Y(n_2327)
);

INVx3_ASAP7_75t_L g2328 ( 
.A(n_1977),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2039),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2039),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2039),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_1860),
.B(n_1707),
.Y(n_2332)
);

INVx5_ASAP7_75t_L g2333 ( 
.A(n_2000),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_1860),
.B(n_1707),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1874),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_1860),
.B(n_1710),
.Y(n_2336)
);

HB1xp67_ASAP7_75t_L g2337 ( 
.A(n_1860),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1860),
.B(n_1710),
.Y(n_2338)
);

BUFx8_ASAP7_75t_L g2339 ( 
.A(n_1880),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2039),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2039),
.Y(n_2341)
);

BUFx3_ASAP7_75t_L g2342 ( 
.A(n_1857),
.Y(n_2342)
);

AND2x4_ASAP7_75t_L g2343 ( 
.A(n_1860),
.B(n_1712),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1874),
.Y(n_2344)
);

INVx5_ASAP7_75t_L g2345 ( 
.A(n_2000),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2039),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_1860),
.B(n_1712),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1911),
.B(n_1526),
.Y(n_2348)
);

AND2x2_ASAP7_75t_SL g2349 ( 
.A(n_2064),
.B(n_1093),
.Y(n_2349)
);

OAI22xp5_ASAP7_75t_SL g2350 ( 
.A1(n_1856),
.A2(n_1220),
.B1(n_1225),
.B2(n_1209),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1911),
.B(n_1531),
.Y(n_2351)
);

OAI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_1860),
.A2(n_1550),
.B1(n_1563),
.B2(n_1532),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1874),
.Y(n_2353)
);

BUFx2_ASAP7_75t_L g2354 ( 
.A(n_1860),
.Y(n_2354)
);

AND2x2_ASAP7_75t_SL g2355 ( 
.A(n_2064),
.B(n_1093),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_1880),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_1860),
.B(n_1114),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1874),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_1880),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_1880),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_1860),
.B(n_1114),
.Y(n_2361)
);

BUFx8_ASAP7_75t_L g2362 ( 
.A(n_1880),
.Y(n_2362)
);

AOI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_1860),
.A2(n_1600),
.B1(n_1622),
.B2(n_1593),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2039),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1874),
.Y(n_2365)
);

OA21x2_ASAP7_75t_L g2366 ( 
.A1(n_1975),
.A2(n_1562),
.B(n_1493),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2039),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1874),
.Y(n_2368)
);

AND2x4_ASAP7_75t_L g2369 ( 
.A(n_1860),
.B(n_1233),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2039),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_1860),
.B(n_1114),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_1860),
.B(n_1118),
.Y(n_2372)
);

OAI22x1_ASAP7_75t_SL g2373 ( 
.A1(n_1856),
.A2(n_1236),
.B1(n_1241),
.B2(n_1233),
.Y(n_2373)
);

BUFx2_ASAP7_75t_L g2374 ( 
.A(n_1860),
.Y(n_2374)
);

HB1xp67_ASAP7_75t_L g2375 ( 
.A(n_1860),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_1977),
.Y(n_2376)
);

OR2x2_ASAP7_75t_L g2377 ( 
.A(n_1860),
.B(n_1174),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1878),
.Y(n_2378)
);

OAI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_1860),
.A2(n_1628),
.B1(n_1629),
.B2(n_1625),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_1911),
.B(n_1640),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_1977),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_1973),
.B(n_1657),
.Y(n_2382)
);

BUFx6f_ASAP7_75t_L g2383 ( 
.A(n_1880),
.Y(n_2383)
);

CKINVDCx8_ASAP7_75t_R g2384 ( 
.A(n_2072),
.Y(n_2384)
);

AND2x2_ASAP7_75t_L g2385 ( 
.A(n_1860),
.B(n_1118),
.Y(n_2385)
);

BUFx6f_ASAP7_75t_L g2386 ( 
.A(n_1880),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1911),
.B(n_1658),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2039),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_1857),
.Y(n_2389)
);

AND2x4_ASAP7_75t_L g2390 ( 
.A(n_1860),
.B(n_1236),
.Y(n_2390)
);

BUFx2_ASAP7_75t_L g2391 ( 
.A(n_1860),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1874),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_2184),
.Y(n_2393)
);

CKINVDCx20_ASAP7_75t_R g2394 ( 
.A(n_2090),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2354),
.B(n_1241),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2203),
.Y(n_2396)
);

CKINVDCx5p33_ASAP7_75t_R g2397 ( 
.A(n_2389),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_2126),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2203),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2208),
.Y(n_2400)
);

HB1xp67_ASAP7_75t_L g2401 ( 
.A(n_2354),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_2295),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_2339),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_2362),
.Y(n_2404)
);

NAND2xp33_ASAP7_75t_R g2405 ( 
.A(n_2212),
.B(n_1659),
.Y(n_2405)
);

BUFx10_ASAP7_75t_L g2406 ( 
.A(n_2177),
.Y(n_2406)
);

BUFx3_ASAP7_75t_L g2407 ( 
.A(n_2374),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_2374),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2100),
.Y(n_2409)
);

HB1xp67_ASAP7_75t_L g2410 ( 
.A(n_2391),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2172),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2120),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_R g2413 ( 
.A(n_2384),
.B(n_1284),
.Y(n_2413)
);

BUFx6f_ASAP7_75t_L g2414 ( 
.A(n_2187),
.Y(n_2414)
);

INVx3_ASAP7_75t_L g2415 ( 
.A(n_2106),
.Y(n_2415)
);

CKINVDCx5p33_ASAP7_75t_R g2416 ( 
.A(n_2316),
.Y(n_2416)
);

CKINVDCx5p33_ASAP7_75t_R g2417 ( 
.A(n_2342),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2187),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_R g2419 ( 
.A(n_2192),
.B(n_1284),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_R g2420 ( 
.A(n_2249),
.B(n_2282),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_2214),
.Y(n_2421)
);

CKINVDCx20_ASAP7_75t_R g2422 ( 
.A(n_2391),
.Y(n_2422)
);

BUFx3_ASAP7_75t_L g2423 ( 
.A(n_2213),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_R g2424 ( 
.A(n_2283),
.B(n_1287),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_2294),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_2290),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2248),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_2205),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_R g2429 ( 
.A(n_2299),
.B(n_1287),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2208),
.Y(n_2430)
);

CKINVDCx20_ASAP7_75t_R g2431 ( 
.A(n_2337),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2238),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2183),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2248),
.Y(n_2434)
);

AO22x2_ASAP7_75t_L g2435 ( 
.A1(n_2151),
.A2(n_1353),
.B1(n_1322),
.B2(n_1594),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_2375),
.Y(n_2436)
);

CKINVDCx5p33_ASAP7_75t_R g2437 ( 
.A(n_2245),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2111),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2238),
.Y(n_2439)
);

CKINVDCx20_ASAP7_75t_R g2440 ( 
.A(n_2204),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2102),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2102),
.Y(n_2442)
);

CKINVDCx5p33_ASAP7_75t_R g2443 ( 
.A(n_2245),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2105),
.Y(n_2444)
);

BUFx6f_ASAP7_75t_L g2445 ( 
.A(n_2235),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_2260),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_2260),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2270),
.Y(n_2448)
);

CKINVDCx5p33_ASAP7_75t_R g2449 ( 
.A(n_2270),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2105),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2127),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_2084),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2131),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2382),
.B(n_1667),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_2275),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_R g2456 ( 
.A(n_2160),
.B(n_1293),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2135),
.Y(n_2457)
);

BUFx2_ASAP7_75t_L g2458 ( 
.A(n_2377),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_2314),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2136),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_2314),
.Y(n_2461)
);

CKINVDCx20_ASAP7_75t_R g2462 ( 
.A(n_2139),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_2322),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2117),
.B(n_1293),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_2322),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_2356),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_2356),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2359),
.Y(n_2468)
);

CKINVDCx20_ASAP7_75t_R g2469 ( 
.A(n_2207),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2359),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2108),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2360),
.Y(n_2472)
);

CKINVDCx20_ASAP7_75t_R g2473 ( 
.A(n_2209),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2108),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_2360),
.Y(n_2475)
);

CKINVDCx20_ASAP7_75t_R g2476 ( 
.A(n_2309),
.Y(n_2476)
);

AND3x2_ASAP7_75t_L g2477 ( 
.A(n_2266),
.B(n_1311),
.C(n_1295),
.Y(n_2477)
);

CKINVDCx20_ASAP7_75t_R g2478 ( 
.A(n_2350),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_2383),
.Y(n_2479)
);

AND2x4_ASAP7_75t_L g2480 ( 
.A(n_2145),
.B(n_1158),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_2383),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2132),
.B(n_1295),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2087),
.B(n_1694),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_R g2484 ( 
.A(n_2377),
.B(n_1311),
.Y(n_2484)
);

NOR2xp33_ASAP7_75t_R g2485 ( 
.A(n_2287),
.B(n_1319),
.Y(n_2485)
);

OAI22xp33_ASAP7_75t_L g2486 ( 
.A1(n_2151),
.A2(n_2152),
.B1(n_2138),
.B2(n_2164),
.Y(n_2486)
);

HB1xp67_ASAP7_75t_L g2487 ( 
.A(n_2133),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2386),
.Y(n_2488)
);

NOR2xp33_ASAP7_75t_R g2489 ( 
.A(n_2312),
.B(n_1319),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2110),
.Y(n_2490)
);

NAND2xp33_ASAP7_75t_SL g2491 ( 
.A(n_2133),
.B(n_2140),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_R g2492 ( 
.A(n_2083),
.B(n_1403),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2265),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_2386),
.Y(n_2494)
);

CKINVDCx20_ASAP7_75t_R g2495 ( 
.A(n_2241),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_2373),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_R g2497 ( 
.A(n_2116),
.B(n_1403),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_2170),
.Y(n_2498)
);

CKINVDCx20_ASAP7_75t_R g2499 ( 
.A(n_2258),
.Y(n_2499)
);

BUFx3_ASAP7_75t_L g2500 ( 
.A(n_2213),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2110),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2378),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_R g2503 ( 
.A(n_2328),
.B(n_1509),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2138),
.Y(n_2504)
);

BUFx2_ASAP7_75t_L g2505 ( 
.A(n_2376),
.Y(n_2505)
);

INVx1_ASAP7_75t_SL g2506 ( 
.A(n_2153),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2301),
.Y(n_2507)
);

NAND2xp33_ASAP7_75t_R g2508 ( 
.A(n_2305),
.B(n_1073),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_R g2509 ( 
.A(n_2381),
.B(n_1509),
.Y(n_2509)
);

HB1xp67_ASAP7_75t_L g2510 ( 
.A(n_2137),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2378),
.Y(n_2511)
);

CKINVDCx16_ASAP7_75t_R g2512 ( 
.A(n_2276),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2301),
.Y(n_2513)
);

CKINVDCx5p33_ASAP7_75t_R g2514 ( 
.A(n_2107),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_2107),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_2125),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2125),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_2129),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2147),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_2129),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2148),
.Y(n_2521)
);

CKINVDCx5p33_ASAP7_75t_R g2522 ( 
.A(n_2141),
.Y(n_2522)
);

BUFx2_ASAP7_75t_L g2523 ( 
.A(n_2112),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2150),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_2141),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2144),
.Y(n_2526)
);

INVx3_ASAP7_75t_L g2527 ( 
.A(n_2109),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2085),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2144),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2088),
.Y(n_2530)
);

BUFx2_ASAP7_75t_L g2531 ( 
.A(n_2114),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2313),
.Y(n_2532)
);

NAND2xp33_ASAP7_75t_R g2533 ( 
.A(n_2239),
.B(n_1074),
.Y(n_2533)
);

CKINVDCx20_ASAP7_75t_R g2534 ( 
.A(n_2146),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_2146),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_2154),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_R g2537 ( 
.A(n_2280),
.B(n_1569),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2154),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_2156),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_2156),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2318),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_2165),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_2165),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2319),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_2169),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_2169),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2320),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2175),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_R g2549 ( 
.A(n_2302),
.B(n_1569),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2327),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2335),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2267),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_2175),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2344),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2142),
.Y(n_2555)
);

CKINVDCx20_ASAP7_75t_R g2556 ( 
.A(n_2232),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_2232),
.Y(n_2557)
);

BUFx2_ASAP7_75t_L g2558 ( 
.A(n_2092),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_2247),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2353),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2247),
.Y(n_2561)
);

CKINVDCx5p33_ASAP7_75t_R g2562 ( 
.A(n_2254),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2254),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2255),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2255),
.Y(n_2565)
);

CKINVDCx5p33_ASAP7_75t_R g2566 ( 
.A(n_2098),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2352),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_2379),
.Y(n_2568)
);

CKINVDCx16_ASAP7_75t_R g2569 ( 
.A(n_2369),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2143),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_2349),
.Y(n_2571)
);

BUFx4f_ASAP7_75t_L g2572 ( 
.A(n_2235),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2355),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_2390),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2358),
.Y(n_2575)
);

BUFx3_ASAP7_75t_L g2576 ( 
.A(n_2185),
.Y(n_2576)
);

CKINVDCx5p33_ASAP7_75t_R g2577 ( 
.A(n_2250),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2365),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2268),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_R g2580 ( 
.A(n_2297),
.B(n_2235),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2368),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_2363),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2392),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2326),
.B(n_1665),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2103),
.Y(n_2585)
);

BUFx2_ASAP7_75t_L g2586 ( 
.A(n_2092),
.Y(n_2586)
);

CKINVDCx20_ASAP7_75t_R g2587 ( 
.A(n_2206),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_2332),
.Y(n_2588)
);

CKINVDCx5p33_ASAP7_75t_R g2589 ( 
.A(n_2336),
.Y(n_2589)
);

AOI21x1_ASAP7_75t_L g2590 ( 
.A1(n_2262),
.A2(n_2366),
.B(n_2162),
.Y(n_2590)
);

BUFx3_ASAP7_75t_L g2591 ( 
.A(n_2185),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2246),
.Y(n_2592)
);

NOR2xp67_ASAP7_75t_L g2593 ( 
.A(n_2277),
.B(n_265),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2343),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_2347),
.Y(n_2595)
);

NAND2x1p5_ASAP7_75t_L g2596 ( 
.A(n_2186),
.B(n_1178),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2225),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_2092),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2233),
.Y(n_2599)
);

OAI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_2159),
.A2(n_1583),
.B1(n_1589),
.B2(n_1571),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2246),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2163),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2166),
.Y(n_2603)
);

NOR2xp67_ASAP7_75t_L g2604 ( 
.A(n_2279),
.B(n_266),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2334),
.B(n_1571),
.Y(n_2605)
);

CKINVDCx16_ASAP7_75t_R g2606 ( 
.A(n_2306),
.Y(n_2606)
);

INVx2_ASAP7_75t_SL g2607 ( 
.A(n_2338),
.Y(n_2607)
);

BUFx10_ASAP7_75t_L g2608 ( 
.A(n_2215),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2311),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_2297),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2304),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_2227),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_2285),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_2307),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2271),
.B(n_1703),
.Y(n_2615)
);

CKINVDCx5p33_ASAP7_75t_R g2616 ( 
.A(n_2310),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2167),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_2300),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2308),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_2178),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2186),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2176),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2181),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2196),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2246),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2149),
.Y(n_2626)
);

HB1xp67_ASAP7_75t_L g2627 ( 
.A(n_2130),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_2196),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_R g2629 ( 
.A(n_2263),
.B(n_1583),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_2197),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2190),
.Y(n_2631)
);

AND2x2_ASAP7_75t_SL g2632 ( 
.A(n_2357),
.B(n_1589),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_2197),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_2217),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2199),
.Y(n_2635)
);

INVx3_ASAP7_75t_L g2636 ( 
.A(n_2263),
.Y(n_2636)
);

CKINVDCx5p33_ASAP7_75t_R g2637 ( 
.A(n_2217),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2200),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2281),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_R g2640 ( 
.A(n_2263),
.B(n_1597),
.Y(n_2640)
);

INVx3_ASAP7_75t_L g2641 ( 
.A(n_2228),
.Y(n_2641)
);

INVxp67_ASAP7_75t_L g2642 ( 
.A(n_2261),
.Y(n_2642)
);

CKINVDCx20_ASAP7_75t_R g2643 ( 
.A(n_2118),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2155),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2210),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2158),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2095),
.B(n_1597),
.Y(n_2647)
);

BUFx10_ASAP7_75t_L g2648 ( 
.A(n_2096),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_2284),
.Y(n_2649)
);

INVxp67_ASAP7_75t_L g2650 ( 
.A(n_2361),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2168),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2216),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2173),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2097),
.B(n_1598),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_2286),
.Y(n_2655)
);

BUFx6f_ASAP7_75t_L g2656 ( 
.A(n_2262),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2101),
.B(n_1598),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2219),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_2104),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2226),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_2104),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2180),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2231),
.Y(n_2663)
);

CKINVDCx20_ASAP7_75t_R g2664 ( 
.A(n_2298),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2240),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2182),
.Y(n_2666)
);

CKINVDCx16_ASAP7_75t_R g2667 ( 
.A(n_2371),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2242),
.Y(n_2668)
);

CKINVDCx20_ASAP7_75t_R g2669 ( 
.A(n_2303),
.Y(n_2669)
);

XNOR2xp5_ASAP7_75t_L g2670 ( 
.A(n_2194),
.B(n_1614),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2251),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2252),
.Y(n_2672)
);

AND2x4_ASAP7_75t_L g2673 ( 
.A(n_2091),
.B(n_1158),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_2115),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_2273),
.Y(n_2675)
);

NAND2xp33_ASAP7_75t_R g2676 ( 
.A(n_2372),
.B(n_1077),
.Y(n_2676)
);

CKINVDCx5p33_ASAP7_75t_R g2677 ( 
.A(n_2123),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2189),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2385),
.Y(n_2679)
);

CKINVDCx20_ASAP7_75t_R g2680 ( 
.A(n_2288),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2257),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2122),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2124),
.Y(n_2683)
);

CKINVDCx20_ASAP7_75t_R g2684 ( 
.A(n_2269),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2128),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2113),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2157),
.Y(n_2687)
);

CKINVDCx20_ASAP7_75t_R g2688 ( 
.A(n_2333),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2193),
.Y(n_2689)
);

CKINVDCx20_ASAP7_75t_R g2690 ( 
.A(n_2333),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_2234),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2211),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2234),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2218),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2220),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2222),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2333),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2345),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2223),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2224),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_2345),
.Y(n_2701)
);

NAND2xp33_ASAP7_75t_R g2702 ( 
.A(n_2162),
.B(n_1078),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2230),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_2345),
.Y(n_2704)
);

CKINVDCx5p33_ASAP7_75t_R g2705 ( 
.A(n_2099),
.Y(n_2705)
);

BUFx10_ASAP7_75t_L g2706 ( 
.A(n_2237),
.Y(n_2706)
);

INVxp67_ASAP7_75t_L g2707 ( 
.A(n_2321),
.Y(n_2707)
);

CKINVDCx5p33_ASAP7_75t_R g2708 ( 
.A(n_2229),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_2198),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_R g2710 ( 
.A(n_2198),
.B(n_1614),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_2198),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2236),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2324),
.B(n_1079),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2325),
.Y(n_2714)
);

NAND3xp33_ASAP7_75t_L g2715 ( 
.A(n_2171),
.B(n_1084),
.C(n_1083),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2366),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2119),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_2348),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2264),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2086),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2351),
.Y(n_2721)
);

CKINVDCx20_ASAP7_75t_R g2722 ( 
.A(n_2380),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2387),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_2179),
.Y(n_2724)
);

CKINVDCx20_ASAP7_75t_R g2725 ( 
.A(n_2195),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_2191),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2221),
.Y(n_2727)
);

CKINVDCx5p33_ASAP7_75t_R g2728 ( 
.A(n_2201),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_2228),
.Y(n_2729)
);

HB1xp67_ASAP7_75t_L g2730 ( 
.A(n_2244),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2089),
.Y(n_2731)
);

CKINVDCx20_ASAP7_75t_R g2732 ( 
.A(n_2259),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2174),
.A2(n_1663),
.B1(n_1683),
.B2(n_1634),
.Y(n_2733)
);

BUFx6f_ASAP7_75t_L g2734 ( 
.A(n_2293),
.Y(n_2734)
);

HB1xp67_ASAP7_75t_L g2735 ( 
.A(n_2134),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2093),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_2202),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_R g2738 ( 
.A(n_2278),
.B(n_1634),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2243),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2253),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2315),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_2256),
.Y(n_2742)
);

CKINVDCx5p33_ASAP7_75t_R g2743 ( 
.A(n_2121),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2317),
.Y(n_2744)
);

CKINVDCx20_ASAP7_75t_R g2745 ( 
.A(n_2174),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2323),
.Y(n_2746)
);

HB1xp67_ASAP7_75t_L g2747 ( 
.A(n_2094),
.Y(n_2747)
);

BUFx2_ASAP7_75t_L g2748 ( 
.A(n_2293),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2329),
.Y(n_2749)
);

CKINVDCx6p67_ASAP7_75t_R g2750 ( 
.A(n_2228),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2330),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_2331),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2188),
.B(n_1197),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2340),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_2341),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_2346),
.Y(n_2756)
);

NOR2x1p5_ASAP7_75t_L g2757 ( 
.A(n_2364),
.B(n_1085),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2367),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_2370),
.Y(n_2759)
);

CKINVDCx20_ASAP7_75t_R g2760 ( 
.A(n_2388),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2293),
.Y(n_2761)
);

CKINVDCx20_ASAP7_75t_R g2762 ( 
.A(n_2272),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_2274),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_R g2764 ( 
.A(n_2291),
.B(n_1663),
.Y(n_2764)
);

CKINVDCx11_ASAP7_75t_R g2765 ( 
.A(n_2289),
.Y(n_2765)
);

CKINVDCx5p33_ASAP7_75t_R g2766 ( 
.A(n_2296),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2292),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2292),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2161),
.Y(n_2769)
);

INVx2_ASAP7_75t_SL g2770 ( 
.A(n_2354),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2184),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2132),
.B(n_1683),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_2184),
.Y(n_2773)
);

CKINVDCx5p33_ASAP7_75t_R g2774 ( 
.A(n_2184),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2203),
.Y(n_2775)
);

NOR2xp33_ASAP7_75t_SL g2776 ( 
.A(n_2126),
.B(n_1702),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_2184),
.Y(n_2777)
);

OA21x2_ASAP7_75t_L g2778 ( 
.A1(n_2100),
.A2(n_1089),
.B(n_1080),
.Y(n_2778)
);

BUFx10_ASAP7_75t_L g2779 ( 
.A(n_2126),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_R g2780 ( 
.A(n_2126),
.B(n_1702),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2203),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2354),
.B(n_1708),
.Y(n_2782)
);

AND2x6_ASAP7_75t_L g2783 ( 
.A(n_2203),
.B(n_1178),
.Y(n_2783)
);

CKINVDCx5p33_ASAP7_75t_R g2784 ( 
.A(n_2184),
.Y(n_2784)
);

INVxp67_ASAP7_75t_L g2785 ( 
.A(n_2354),
.Y(n_2785)
);

BUFx3_ASAP7_75t_L g2786 ( 
.A(n_2534),
.Y(n_2786)
);

CKINVDCx11_ASAP7_75t_R g2787 ( 
.A(n_2394),
.Y(n_2787)
);

INVx1_ASAP7_75t_SL g2788 ( 
.A(n_2407),
.Y(n_2788)
);

AND2x4_ASAP7_75t_L g2789 ( 
.A(n_2685),
.B(n_1708),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2396),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2486),
.B(n_1088),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2519),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2521),
.Y(n_2793)
);

AOI22xp33_ASAP7_75t_L g2794 ( 
.A1(n_2632),
.A2(n_1222),
.B1(n_1269),
.B2(n_1118),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2399),
.B(n_1091),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2400),
.Y(n_2796)
);

AND2x6_ASAP7_75t_L g2797 ( 
.A(n_2445),
.B(n_1263),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2430),
.B(n_1092),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2432),
.Y(n_2799)
);

BUFx3_ASAP7_75t_L g2800 ( 
.A(n_2556),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_L g2801 ( 
.A(n_2414),
.Y(n_2801)
);

BUFx2_ASAP7_75t_L g2802 ( 
.A(n_2422),
.Y(n_2802)
);

OR2x6_ASAP7_75t_L g2803 ( 
.A(n_2770),
.B(n_2785),
.Y(n_2803)
);

CKINVDCx16_ASAP7_75t_R g2804 ( 
.A(n_2429),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_SL g2805 ( 
.A(n_2785),
.B(n_1095),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2524),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2458),
.B(n_1222),
.Y(n_2807)
);

OAI22xp5_ASAP7_75t_L g2808 ( 
.A1(n_2439),
.A2(n_1338),
.B1(n_1369),
.B2(n_1263),
.Y(n_2808)
);

CKINVDCx6p67_ASAP7_75t_R g2809 ( 
.A(n_2765),
.Y(n_2809)
);

NAND3xp33_ASAP7_75t_SL g2810 ( 
.A(n_2484),
.B(n_1097),
.C(n_1096),
.Y(n_2810)
);

AO21x2_ASAP7_75t_L g2811 ( 
.A1(n_2409),
.A2(n_2590),
.B(n_2427),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2528),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2414),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2642),
.B(n_1222),
.Y(n_2814)
);

AND2x6_ASAP7_75t_L g2815 ( 
.A(n_2445),
.B(n_1338),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2441),
.Y(n_2816)
);

BUFx3_ASAP7_75t_L g2817 ( 
.A(n_2459),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2442),
.B(n_1104),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2444),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2642),
.B(n_1269),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_L g2821 ( 
.A(n_2667),
.B(n_1110),
.Y(n_2821)
);

AND2x6_ASAP7_75t_L g2822 ( 
.A(n_2445),
.B(n_1369),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2530),
.Y(n_2823)
);

INVx4_ASAP7_75t_L g2824 ( 
.A(n_2461),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2532),
.Y(n_2825)
);

AND2x4_ASAP7_75t_L g2826 ( 
.A(n_2727),
.B(n_1435),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2629),
.B(n_1113),
.Y(n_2827)
);

BUFx3_ASAP7_75t_L g2828 ( 
.A(n_2463),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2450),
.B(n_2471),
.Y(n_2829)
);

BUFx3_ASAP7_75t_L g2830 ( 
.A(n_2465),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_L g2831 ( 
.A(n_2677),
.B(n_1115),
.Y(n_2831)
);

CKINVDCx16_ASAP7_75t_R g2832 ( 
.A(n_2413),
.Y(n_2832)
);

AND3x2_ASAP7_75t_L g2833 ( 
.A(n_2776),
.B(n_1112),
.C(n_1105),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2750),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2541),
.Y(n_2835)
);

OAI22xp33_ASAP7_75t_SL g2836 ( 
.A1(n_2612),
.A2(n_1116),
.B1(n_1122),
.B2(n_1117),
.Y(n_2836)
);

AO22x2_ASAP7_75t_L g2837 ( 
.A1(n_2395),
.A2(n_1204),
.B1(n_1212),
.B2(n_1184),
.Y(n_2837)
);

AND2x6_ASAP7_75t_L g2838 ( 
.A(n_2734),
.B(n_1435),
.Y(n_2838)
);

AOI22xp33_ASAP7_75t_L g2839 ( 
.A1(n_2605),
.A2(n_1283),
.B1(n_1305),
.B2(n_1269),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2544),
.Y(n_2840)
);

INVx3_ASAP7_75t_L g2841 ( 
.A(n_2783),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_SL g2842 ( 
.A(n_2640),
.B(n_1127),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2474),
.B(n_1145),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_SL g2844 ( 
.A(n_2436),
.B(n_1146),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2547),
.Y(n_2845)
);

BUFx3_ASAP7_75t_L g2846 ( 
.A(n_2466),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2490),
.Y(n_2847)
);

BUFx10_ASAP7_75t_L g2848 ( 
.A(n_2393),
.Y(n_2848)
);

INVx1_ASAP7_75t_SL g2849 ( 
.A(n_2401),
.Y(n_2849)
);

AND2x4_ASAP7_75t_L g2850 ( 
.A(n_2707),
.B(n_1464),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2501),
.B(n_1147),
.Y(n_2851)
);

AOI22xp33_ASAP7_75t_L g2852 ( 
.A1(n_2464),
.A2(n_1305),
.B1(n_1344),
.B2(n_1283),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2550),
.Y(n_2853)
);

INVx5_ASAP7_75t_L g2854 ( 
.A(n_2783),
.Y(n_2854)
);

INVx4_ASAP7_75t_L g2855 ( 
.A(n_2467),
.Y(n_2855)
);

OAI22xp33_ASAP7_75t_L g2856 ( 
.A1(n_2733),
.A2(n_1152),
.B1(n_1153),
.B2(n_1148),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2582),
.B(n_1154),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2502),
.B(n_1157),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2551),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2511),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2775),
.B(n_1159),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2781),
.B(n_1162),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2783),
.Y(n_2863)
);

BUFx3_ASAP7_75t_L g2864 ( 
.A(n_2468),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2554),
.Y(n_2865)
);

BUFx2_ASAP7_75t_L g2866 ( 
.A(n_2431),
.Y(n_2866)
);

BUFx3_ASAP7_75t_L g2867 ( 
.A(n_2470),
.Y(n_2867)
);

BUFx6f_ASAP7_75t_L g2868 ( 
.A(n_2414),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_SL g2869 ( 
.A(n_2714),
.B(n_1165),
.Y(n_2869)
);

INVxp67_ASAP7_75t_L g2870 ( 
.A(n_2408),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2560),
.B(n_1166),
.Y(n_2871)
);

INVxp33_ASAP7_75t_L g2872 ( 
.A(n_2492),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2575),
.Y(n_2873)
);

OR2x2_ASAP7_75t_L g2874 ( 
.A(n_2782),
.B(n_1354),
.Y(n_2874)
);

INVx3_ASAP7_75t_L g2875 ( 
.A(n_2783),
.Y(n_2875)
);

INVx4_ASAP7_75t_SL g2876 ( 
.A(n_2783),
.Y(n_2876)
);

INVx2_ASAP7_75t_SL g2877 ( 
.A(n_2406),
.Y(n_2877)
);

NOR2x1p5_ASAP7_75t_L g2878 ( 
.A(n_2771),
.B(n_2773),
.Y(n_2878)
);

HB1xp67_ASAP7_75t_L g2879 ( 
.A(n_2410),
.Y(n_2879)
);

OR2x2_ASAP7_75t_L g2880 ( 
.A(n_2512),
.B(n_1474),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2415),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2578),
.B(n_1169),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2581),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_SL g2884 ( 
.A(n_2718),
.B(n_1170),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_SL g2885 ( 
.A(n_2721),
.B(n_1173),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_SL g2886 ( 
.A(n_2723),
.B(n_1177),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2583),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2724),
.B(n_1181),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2602),
.B(n_1183),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2603),
.B(n_2617),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2622),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2707),
.B(n_2487),
.Y(n_2892)
);

OR2x2_ASAP7_75t_L g2893 ( 
.A(n_2600),
.B(n_1530),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2623),
.B(n_1188),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2415),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_2472),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2780),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2631),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2635),
.B(n_1192),
.Y(n_2899)
);

AOI22xp33_ASAP7_75t_L g2900 ( 
.A1(n_2647),
.A2(n_1305),
.B1(n_1344),
.B2(n_1283),
.Y(n_2900)
);

BUFx6f_ASAP7_75t_L g2901 ( 
.A(n_2734),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2638),
.B(n_1194),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_SL g2903 ( 
.A(n_2743),
.B(n_1196),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2452),
.B(n_1199),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2645),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2527),
.Y(n_2906)
);

INVx3_ASAP7_75t_L g2907 ( 
.A(n_2527),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2652),
.Y(n_2908)
);

INVx4_ASAP7_75t_L g2909 ( 
.A(n_2475),
.Y(n_2909)
);

INVxp67_ASAP7_75t_SL g2910 ( 
.A(n_2734),
.Y(n_2910)
);

BUFx8_ASAP7_75t_SL g2911 ( 
.A(n_2774),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_L g2912 ( 
.A(n_2569),
.B(n_1203),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2658),
.B(n_1205),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2641),
.Y(n_2914)
);

AO22x2_ASAP7_75t_L g2915 ( 
.A1(n_2418),
.A2(n_1705),
.B1(n_1592),
.B2(n_1237),
.Y(n_2915)
);

INVx2_ASAP7_75t_SL g2916 ( 
.A(n_2406),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2660),
.Y(n_2917)
);

INVx4_ASAP7_75t_L g2918 ( 
.A(n_2479),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2663),
.Y(n_2919)
);

BUFx3_ASAP7_75t_L g2920 ( 
.A(n_2481),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2665),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2668),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2671),
.B(n_1211),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2672),
.B(n_1213),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2681),
.Y(n_2925)
);

CKINVDCx6p67_ASAP7_75t_R g2926 ( 
.A(n_2779),
.Y(n_2926)
);

BUFx3_ASAP7_75t_L g2927 ( 
.A(n_2488),
.Y(n_2927)
);

INVx2_ASAP7_75t_L g2928 ( 
.A(n_2682),
.Y(n_2928)
);

OR2x6_ASAP7_75t_L g2929 ( 
.A(n_2423),
.B(n_1197),
.Y(n_2929)
);

NAND2xp33_ASAP7_75t_L g2930 ( 
.A(n_2710),
.B(n_1214),
.Y(n_2930)
);

INVx5_ASAP7_75t_L g2931 ( 
.A(n_2779),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2683),
.Y(n_2932)
);

BUFx4f_ASAP7_75t_L g2933 ( 
.A(n_2596),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2438),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2451),
.Y(n_2935)
);

INVx3_ASAP7_75t_L g2936 ( 
.A(n_2641),
.Y(n_2936)
);

AND2x4_ASAP7_75t_L g2937 ( 
.A(n_2607),
.B(n_1464),
.Y(n_2937)
);

OAI22xp33_ASAP7_75t_L g2938 ( 
.A1(n_2745),
.A2(n_1219),
.B1(n_1223),
.B2(n_1221),
.Y(n_2938)
);

BUFx2_ASAP7_75t_L g2939 ( 
.A(n_2497),
.Y(n_2939)
);

INVx1_ASAP7_75t_SL g2940 ( 
.A(n_2764),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2687),
.B(n_1226),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2747),
.B(n_1228),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_2437),
.B(n_1229),
.Y(n_2943)
);

HB1xp67_ASAP7_75t_L g2944 ( 
.A(n_2494),
.Y(n_2944)
);

OR2x2_ASAP7_75t_L g2945 ( 
.A(n_2606),
.B(n_1230),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2453),
.Y(n_2946)
);

INVx1_ASAP7_75t_SL g2947 ( 
.A(n_2503),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2654),
.B(n_1344),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2778),
.Y(n_2949)
);

BUFx3_ASAP7_75t_L g2950 ( 
.A(n_2576),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_SL g2951 ( 
.A(n_2443),
.B(n_1234),
.Y(n_2951)
);

AND2x2_ASAP7_75t_L g2952 ( 
.A(n_2657),
.B(n_1401),
.Y(n_2952)
);

CKINVDCx6p67_ASAP7_75t_R g2953 ( 
.A(n_2440),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2446),
.B(n_1238),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2730),
.B(n_1239),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2457),
.Y(n_2956)
);

NOR2xp33_ASAP7_75t_L g2957 ( 
.A(n_2686),
.B(n_1243),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2778),
.Y(n_2958)
);

INVxp33_ASAP7_75t_L g2959 ( 
.A(n_2509),
.Y(n_2959)
);

AND3x2_ASAP7_75t_L g2960 ( 
.A(n_2482),
.B(n_1121),
.C(n_1119),
.Y(n_2960)
);

INVxp67_ASAP7_75t_SL g2961 ( 
.A(n_2760),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2460),
.Y(n_2962)
);

AND2x2_ASAP7_75t_L g2963 ( 
.A(n_2506),
.B(n_1401),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2708),
.B(n_1244),
.Y(n_2964)
);

INVx3_ASAP7_75t_L g2965 ( 
.A(n_2729),
.Y(n_2965)
);

NOR2xp33_ASAP7_75t_L g2966 ( 
.A(n_2679),
.B(n_1246),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2555),
.Y(n_2967)
);

CKINVDCx20_ASAP7_75t_R g2968 ( 
.A(n_2495),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2570),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2673),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2626),
.Y(n_2971)
);

INVx2_ASAP7_75t_SL g2972 ( 
.A(n_2514),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2644),
.Y(n_2973)
);

AND2x4_ASAP7_75t_L g2974 ( 
.A(n_2735),
.B(n_1465),
.Y(n_2974)
);

INVx3_ASAP7_75t_L g2975 ( 
.A(n_2729),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2673),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2753),
.B(n_1249),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2772),
.B(n_1252),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2620),
.B(n_1253),
.Y(n_2979)
);

BUFx2_ASAP7_75t_L g2980 ( 
.A(n_2419),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2692),
.Y(n_2981)
);

INVx4_ASAP7_75t_L g2982 ( 
.A(n_2498),
.Y(n_2982)
);

INVx4_ASAP7_75t_L g2983 ( 
.A(n_2621),
.Y(n_2983)
);

INVx3_ASAP7_75t_L g2984 ( 
.A(n_2636),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2694),
.Y(n_2985)
);

AOI21x1_ASAP7_75t_L g2986 ( 
.A1(n_2434),
.A2(n_1138),
.B(n_1111),
.Y(n_2986)
);

BUFx4f_ASAP7_75t_L g2987 ( 
.A(n_2596),
.Y(n_2987)
);

NOR2x1p5_ASAP7_75t_L g2988 ( 
.A(n_2777),
.B(n_1260),
.Y(n_2988)
);

INVx2_ASAP7_75t_SL g2989 ( 
.A(n_2515),
.Y(n_2989)
);

NAND3x1_ASAP7_75t_L g2990 ( 
.A(n_2477),
.B(n_1136),
.C(n_1132),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2627),
.B(n_1401),
.Y(n_2991)
);

AND2x6_ASAP7_75t_L g2992 ( 
.A(n_2592),
.B(n_1465),
.Y(n_2992)
);

AOI22xp5_ASAP7_75t_L g2993 ( 
.A1(n_2435),
.A2(n_1271),
.B1(n_1272),
.B2(n_1268),
.Y(n_2993)
);

AND2x2_ASAP7_75t_L g2994 ( 
.A(n_2597),
.B(n_2599),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2646),
.Y(n_2995)
);

AND2x4_ASAP7_75t_L g2996 ( 
.A(n_2757),
.B(n_1478),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2651),
.Y(n_2997)
);

NAND2xp33_ASAP7_75t_L g2998 ( 
.A(n_2761),
.B(n_1274),
.Y(n_2998)
);

BUFx8_ASAP7_75t_SL g2999 ( 
.A(n_2784),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2753),
.B(n_1275),
.Y(n_3000)
);

INVx4_ASAP7_75t_L g3001 ( 
.A(n_2624),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2447),
.B(n_1277),
.Y(n_3002)
);

BUFx3_ASAP7_75t_L g3003 ( 
.A(n_2591),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2653),
.Y(n_3004)
);

OAI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2448),
.A2(n_1282),
.B1(n_1286),
.B2(n_1281),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2435),
.A2(n_1664),
.B1(n_1698),
.B2(n_1445),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2695),
.Y(n_3007)
);

BUFx6f_ASAP7_75t_L g3008 ( 
.A(n_2656),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2700),
.Y(n_3009)
);

AND2x4_ASAP7_75t_L g3010 ( 
.A(n_2650),
.B(n_1478),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2650),
.B(n_1288),
.Y(n_3011)
);

INVx2_ASAP7_75t_SL g3012 ( 
.A(n_2516),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2712),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_2566),
.B(n_1296),
.Y(n_3014)
);

NAND2xp33_ASAP7_75t_SL g3015 ( 
.A(n_2580),
.B(n_1298),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_SL g3016 ( 
.A(n_2449),
.B(n_1304),
.Y(n_3016)
);

CKINVDCx5p33_ASAP7_75t_R g3017 ( 
.A(n_2403),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2717),
.Y(n_3018)
);

OAI22xp33_ASAP7_75t_L g3019 ( 
.A1(n_2533),
.A2(n_1313),
.B1(n_1314),
.B2(n_1310),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2493),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2552),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2662),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2666),
.Y(n_3023)
);

AOI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2435),
.A2(n_1317),
.B1(n_1318),
.B2(n_1315),
.Y(n_3024)
);

NOR2xp33_ASAP7_75t_L g3025 ( 
.A(n_2567),
.B(n_1320),
.Y(n_3025)
);

INVx4_ASAP7_75t_L g3026 ( 
.A(n_2628),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2483),
.B(n_1330),
.Y(n_3027)
);

BUFx6f_ASAP7_75t_L g3028 ( 
.A(n_2656),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_2568),
.B(n_1445),
.Y(n_3029)
);

INVxp67_ASAP7_75t_SL g3030 ( 
.A(n_2499),
.Y(n_3030)
);

NAND2xp33_ASAP7_75t_L g3031 ( 
.A(n_2738),
.B(n_1331),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2678),
.Y(n_3032)
);

INVx4_ASAP7_75t_L g3033 ( 
.A(n_2630),
.Y(n_3033)
);

BUFx3_ASAP7_75t_L g3034 ( 
.A(n_2500),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_2412),
.B(n_1332),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2689),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2454),
.B(n_1333),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2696),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2699),
.Y(n_3039)
);

NOR2xp33_ASAP7_75t_L g3040 ( 
.A(n_2574),
.B(n_1342),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2703),
.Y(n_3041)
);

BUFx2_ASAP7_75t_L g3042 ( 
.A(n_2485),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2720),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2480),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2725),
.B(n_1350),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2656),
.Y(n_3046)
);

BUFx2_ASAP7_75t_L g3047 ( 
.A(n_2456),
.Y(n_3047)
);

INVx6_ASAP7_75t_L g3048 ( 
.A(n_2608),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2731),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2480),
.B(n_1352),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2648),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2751),
.Y(n_3052)
);

AND2x4_ASAP7_75t_L g3053 ( 
.A(n_2592),
.B(n_1595),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2713),
.B(n_1358),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2726),
.B(n_1360),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2674),
.B(n_1366),
.Y(n_3056)
);

INVx5_ASAP7_75t_L g3057 ( 
.A(n_2608),
.Y(n_3057)
);

INVx4_ASAP7_75t_L g3058 ( 
.A(n_2633),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2648),
.Y(n_3059)
);

INVx2_ASAP7_75t_SL g3060 ( 
.A(n_2517),
.Y(n_3060)
);

INVxp33_ASAP7_75t_L g3061 ( 
.A(n_2489),
.Y(n_3061)
);

AO22x2_ASAP7_75t_L g3062 ( 
.A1(n_2549),
.A2(n_1254),
.B1(n_1351),
.B2(n_1237),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2584),
.B(n_1367),
.Y(n_3063)
);

INVx1_ASAP7_75t_SL g3064 ( 
.A(n_2659),
.Y(n_3064)
);

INVx2_ASAP7_75t_SL g3065 ( 
.A(n_2518),
.Y(n_3065)
);

CKINVDCx5p33_ASAP7_75t_R g3066 ( 
.A(n_2404),
.Y(n_3066)
);

OR2x2_ASAP7_75t_L g3067 ( 
.A(n_2609),
.B(n_1368),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_2636),
.Y(n_3068)
);

BUFx6f_ASAP7_75t_L g3069 ( 
.A(n_2716),
.Y(n_3069)
);

INVx1_ASAP7_75t_SL g3070 ( 
.A(n_2661),
.Y(n_3070)
);

AND3x2_ASAP7_75t_L g3071 ( 
.A(n_2424),
.B(n_1150),
.C(n_1137),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2728),
.B(n_1373),
.Y(n_3072)
);

AOI22xp33_ASAP7_75t_L g3073 ( 
.A1(n_2732),
.A2(n_1664),
.B1(n_1698),
.B2(n_1445),
.Y(n_3073)
);

INVx1_ASAP7_75t_SL g3074 ( 
.A(n_2705),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2736),
.Y(n_3075)
);

AOI22xp33_ASAP7_75t_L g3076 ( 
.A1(n_2722),
.A2(n_1698),
.B1(n_1664),
.B2(n_1647),
.Y(n_3076)
);

BUFx8_ASAP7_75t_SL g3077 ( 
.A(n_2402),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2741),
.Y(n_3078)
);

BUFx6f_ASAP7_75t_L g3079 ( 
.A(n_2716),
.Y(n_3079)
);

INVx2_ASAP7_75t_SL g3080 ( 
.A(n_2520),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2510),
.B(n_1375),
.Y(n_3081)
);

BUFx3_ASAP7_75t_L g3082 ( 
.A(n_2688),
.Y(n_3082)
);

AND2x6_ASAP7_75t_L g3083 ( 
.A(n_2601),
.B(n_1595),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2758),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2766),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2510),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_2716),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2593),
.B(n_1376),
.Y(n_3088)
);

BUFx6f_ASAP7_75t_L g3089 ( 
.A(n_2572),
.Y(n_3089)
);

OR2x6_ASAP7_75t_L g3090 ( 
.A(n_2505),
.B(n_1254),
.Y(n_3090)
);

INVx2_ASAP7_75t_SL g3091 ( 
.A(n_2522),
.Y(n_3091)
);

AO22x2_ASAP7_75t_L g3092 ( 
.A1(n_2537),
.A2(n_1356),
.B1(n_1461),
.B2(n_1351),
.Y(n_3092)
);

OR2x2_ASAP7_75t_L g3093 ( 
.A(n_2670),
.B(n_1377),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2615),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_SL g3095 ( 
.A(n_2737),
.B(n_1381),
.Y(n_3095)
);

BUFx4f_ASAP7_75t_L g3096 ( 
.A(n_2523),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2744),
.Y(n_3097)
);

AND2x4_ASAP7_75t_L g3098 ( 
.A(n_2601),
.B(n_1647),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2604),
.B(n_1384),
.Y(n_3099)
);

NOR2xp33_ASAP7_75t_L g3100 ( 
.A(n_2531),
.B(n_1390),
.Y(n_3100)
);

NOR2x1p5_ASAP7_75t_L g3101 ( 
.A(n_2421),
.B(n_1395),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2577),
.B(n_1400),
.Y(n_3102)
);

NAND3xp33_ASAP7_75t_L g3103 ( 
.A(n_2702),
.B(n_1258),
.C(n_1257),
.Y(n_3103)
);

BUFx3_ASAP7_75t_L g3104 ( 
.A(n_2690),
.Y(n_3104)
);

OAI22xp33_ASAP7_75t_L g3105 ( 
.A1(n_2508),
.A2(n_1402),
.B1(n_1407),
.B2(n_1404),
.Y(n_3105)
);

AND2x2_ASAP7_75t_SL g3106 ( 
.A(n_2572),
.B(n_1111),
.Y(n_3106)
);

BUFx3_ASAP7_75t_L g3107 ( 
.A(n_2634),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2625),
.Y(n_3108)
);

CKINVDCx5p33_ASAP7_75t_R g3109 ( 
.A(n_2428),
.Y(n_3109)
);

AND2x4_ASAP7_75t_L g3110 ( 
.A(n_2625),
.B(n_1711),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2746),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_2739),
.B(n_1410),
.Y(n_3112)
);

AND2x6_ASAP7_75t_L g3113 ( 
.A(n_2748),
.B(n_1711),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2579),
.B(n_1412),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2749),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2752),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2715),
.B(n_1419),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2754),
.Y(n_3118)
);

AND2x2_ASAP7_75t_L g3119 ( 
.A(n_2613),
.B(n_1421),
.Y(n_3119)
);

INVxp33_ASAP7_75t_L g3120 ( 
.A(n_2420),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2740),
.B(n_2742),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2767),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2755),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2756),
.Y(n_3124)
);

NOR2xp33_ASAP7_75t_L g3125 ( 
.A(n_2587),
.B(n_1422),
.Y(n_3125)
);

AOI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_2491),
.A2(n_1423),
.B1(n_1426),
.B2(n_1424),
.Y(n_3126)
);

INVx6_ASAP7_75t_L g3127 ( 
.A(n_2706),
.Y(n_3127)
);

INVx3_ASAP7_75t_L g3128 ( 
.A(n_2768),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2759),
.Y(n_3129)
);

INVx4_ASAP7_75t_L g3130 ( 
.A(n_2637),
.Y(n_3130)
);

AND2x2_ASAP7_75t_SL g3131 ( 
.A(n_2558),
.B(n_2586),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2706),
.B(n_1428),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2598),
.B(n_2639),
.Y(n_3133)
);

AOI22xp5_ASAP7_75t_L g3134 ( 
.A1(n_2676),
.A2(n_1430),
.B1(n_1432),
.B2(n_1431),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2719),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2763),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2697),
.Y(n_3137)
);

INVx4_ASAP7_75t_SL g3138 ( 
.A(n_2477),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2585),
.B(n_1433),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2698),
.Y(n_3140)
);

BUFx3_ASAP7_75t_L g3141 ( 
.A(n_2525),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2649),
.B(n_1437),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2701),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_L g3144 ( 
.A(n_2588),
.B(n_1438),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_SL g3145 ( 
.A(n_2398),
.B(n_1441),
.Y(n_3145)
);

NOR2xp33_ASAP7_75t_L g3146 ( 
.A(n_2589),
.B(n_1442),
.Y(n_3146)
);

AND2x4_ASAP7_75t_L g3147 ( 
.A(n_2762),
.B(n_1356),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_SL g3148 ( 
.A(n_2455),
.B(n_1447),
.Y(n_3148)
);

OR2x2_ASAP7_75t_L g3149 ( 
.A(n_2397),
.B(n_1449),
.Y(n_3149)
);

BUFx3_ASAP7_75t_L g3150 ( 
.A(n_2526),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2611),
.B(n_1453),
.Y(n_3151)
);

BUFx6f_ASAP7_75t_SL g3152 ( 
.A(n_2426),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2655),
.B(n_1457),
.Y(n_3153)
);

OR2x6_ASAP7_75t_L g3154 ( 
.A(n_2529),
.B(n_1461),
.Y(n_3154)
);

OAI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_2691),
.A2(n_1462),
.B1(n_1466),
.B2(n_1455),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2769),
.B(n_1468),
.Y(n_3156)
);

NOR2xp33_ASAP7_75t_L g3157 ( 
.A(n_2594),
.B(n_1475),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2709),
.B(n_1477),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_L g3159 ( 
.A1(n_2680),
.A2(n_2664),
.B1(n_2669),
.B2(n_2693),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_2595),
.B(n_1479),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_2704),
.B(n_1511),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2711),
.B(n_1480),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2614),
.B(n_1482),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_2416),
.B(n_1486),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2616),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2610),
.B(n_2675),
.Y(n_3166)
);

OR2x2_ASAP7_75t_L g3167 ( 
.A(n_2411),
.B(n_2417),
.Y(n_3167)
);

BUFx3_ASAP7_75t_L g3168 ( 
.A(n_2535),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2618),
.Y(n_3169)
);

NAND2x1p5_ASAP7_75t_L g3170 ( 
.A(n_2536),
.B(n_1511),
.Y(n_3170)
);

HB1xp67_ASAP7_75t_L g3171 ( 
.A(n_2538),
.Y(n_3171)
);

INVx5_ASAP7_75t_L g3172 ( 
.A(n_2539),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2571),
.B(n_1491),
.Y(n_3173)
);

BUFx6f_ASAP7_75t_L g3174 ( 
.A(n_2540),
.Y(n_3174)
);

INVx2_ASAP7_75t_SL g3175 ( 
.A(n_2542),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2619),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2543),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2573),
.B(n_1495),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_2504),
.B(n_1501),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2545),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_L g3181 ( 
.A(n_2643),
.B(n_1505),
.Y(n_3181)
);

NAND3xp33_ASAP7_75t_L g3182 ( 
.A(n_2405),
.B(n_1258),
.C(n_1257),
.Y(n_3182)
);

BUFx6f_ASAP7_75t_L g3183 ( 
.A(n_2546),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2684),
.B(n_1508),
.Y(n_3184)
);

INVx5_ASAP7_75t_L g3185 ( 
.A(n_2565),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2548),
.Y(n_3186)
);

OR2x2_ASAP7_75t_L g3187 ( 
.A(n_2553),
.B(n_1512),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2557),
.Y(n_3188)
);

INVxp67_ASAP7_75t_L g3189 ( 
.A(n_2559),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2561),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2562),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2563),
.Y(n_3192)
);

BUFx6f_ASAP7_75t_L g3193 ( 
.A(n_2564),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2507),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_2513),
.B(n_1513),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2433),
.B(n_1515),
.Y(n_3196)
);

INVx1_ASAP7_75t_SL g3197 ( 
.A(n_2462),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2469),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_2425),
.B(n_1516),
.Y(n_3199)
);

AND2x2_ASAP7_75t_L g3200 ( 
.A(n_2473),
.B(n_1517),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2476),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2478),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2496),
.Y(n_3203)
);

NAND2x1p5_ASAP7_75t_L g3204 ( 
.A(n_2572),
.B(n_1516),
.Y(n_3204)
);

INVx2_ASAP7_75t_SL g3205 ( 
.A(n_2406),
.Y(n_3205)
);

INVx3_ASAP7_75t_L g3206 ( 
.A(n_2750),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_2396),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2685),
.Y(n_3208)
);

NAND2xp33_ASAP7_75t_L g3209 ( 
.A(n_2783),
.B(n_1534),
.Y(n_3209)
);

AOI22xp5_ASAP7_75t_L g3210 ( 
.A1(n_2727),
.A2(n_1523),
.B1(n_1528),
.B2(n_1522),
.Y(n_3210)
);

OR2x6_ASAP7_75t_L g3211 ( 
.A(n_2770),
.B(n_1568),
.Y(n_3211)
);

INVx5_ASAP7_75t_L g3212 ( 
.A(n_2783),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2685),
.Y(n_3213)
);

OAI22xp33_ASAP7_75t_L g3214 ( 
.A1(n_2733),
.A2(n_1537),
.B1(n_1538),
.B2(n_1536),
.Y(n_3214)
);

OAI22xp5_ASAP7_75t_L g3215 ( 
.A1(n_2685),
.A2(n_1568),
.B1(n_1187),
.B2(n_1231),
.Y(n_3215)
);

BUFx3_ASAP7_75t_L g3216 ( 
.A(n_2534),
.Y(n_3216)
);

NOR2x1p5_ASAP7_75t_L g3217 ( 
.A(n_2393),
.B(n_1539),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2685),
.Y(n_3218)
);

AOI22xp5_ASAP7_75t_L g3219 ( 
.A1(n_2727),
.A2(n_1543),
.B1(n_1546),
.B2(n_1542),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2685),
.B(n_1553),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2486),
.B(n_1547),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_2486),
.B(n_1554),
.Y(n_3222)
);

NOR2xp33_ASAP7_75t_L g3223 ( 
.A(n_2486),
.B(n_1555),
.Y(n_3223)
);

INVx2_ASAP7_75t_SL g3224 ( 
.A(n_2406),
.Y(n_3224)
);

INVxp67_ASAP7_75t_SL g3225 ( 
.A(n_2407),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2685),
.Y(n_3226)
);

BUFx10_ASAP7_75t_L g3227 ( 
.A(n_2393),
.Y(n_3227)
);

OR2x2_ASAP7_75t_L g3228 ( 
.A(n_2458),
.B(n_1558),
.Y(n_3228)
);

INVx4_ASAP7_75t_L g3229 ( 
.A(n_2459),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2685),
.Y(n_3230)
);

INVx4_ASAP7_75t_SL g3231 ( 
.A(n_2783),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2396),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_2685),
.Y(n_3233)
);

INVxp33_ASAP7_75t_L g3234 ( 
.A(n_2484),
.Y(n_3234)
);

INVxp67_ASAP7_75t_SL g3235 ( 
.A(n_2407),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_2632),
.A2(n_1564),
.B1(n_1566),
.B2(n_1560),
.Y(n_3236)
);

INVx4_ASAP7_75t_L g3237 ( 
.A(n_2459),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2685),
.B(n_1570),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2685),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2486),
.B(n_1574),
.Y(n_3240)
);

INVx2_ASAP7_75t_SL g3241 ( 
.A(n_2406),
.Y(n_3241)
);

AND2x4_ASAP7_75t_L g3242 ( 
.A(n_2685),
.B(n_1155),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_2486),
.B(n_1575),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2685),
.B(n_1588),
.Y(n_3244)
);

AND2x2_ASAP7_75t_L g3245 ( 
.A(n_2458),
.B(n_1591),
.Y(n_3245)
);

AND2x6_ASAP7_75t_L g3246 ( 
.A(n_2445),
.B(n_1258),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2685),
.B(n_1596),
.Y(n_3247)
);

BUFx6f_ASAP7_75t_L g3248 ( 
.A(n_2414),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2685),
.Y(n_3249)
);

NAND3xp33_ASAP7_75t_SL g3250 ( 
.A(n_2429),
.B(n_1602),
.C(n_1601),
.Y(n_3250)
);

HB1xp67_ASAP7_75t_L g3251 ( 
.A(n_2407),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2685),
.B(n_1605),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2396),
.Y(n_3253)
);

OR2x2_ASAP7_75t_L g3254 ( 
.A(n_2458),
.B(n_1607),
.Y(n_3254)
);

AOI22xp33_ASAP7_75t_L g3255 ( 
.A1(n_2632),
.A2(n_1608),
.B1(n_1615),
.B2(n_1609),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_2486),
.B(n_1616),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2685),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2458),
.B(n_1618),
.Y(n_3258)
);

HB1xp67_ASAP7_75t_L g3259 ( 
.A(n_2407),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2396),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_2685),
.B(n_1619),
.Y(n_3261)
);

AOI22xp33_ASAP7_75t_L g3262 ( 
.A1(n_2632),
.A2(n_1621),
.B1(n_1627),
.B2(n_1623),
.Y(n_3262)
);

OR2x2_ASAP7_75t_L g3263 ( 
.A(n_2458),
.B(n_1631),
.Y(n_3263)
);

BUFx3_ASAP7_75t_L g3264 ( 
.A(n_2534),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2685),
.Y(n_3265)
);

NOR2xp33_ASAP7_75t_L g3266 ( 
.A(n_2486),
.B(n_1632),
.Y(n_3266)
);

INVx3_ASAP7_75t_L g3267 ( 
.A(n_2750),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_2458),
.B(n_1633),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2685),
.B(n_1635),
.Y(n_3269)
);

INVx2_ASAP7_75t_SL g3270 ( 
.A(n_2406),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2685),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_SL g3272 ( 
.A(n_2785),
.B(n_1637),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_2685),
.B(n_1642),
.Y(n_3273)
);

OAI22xp33_ASAP7_75t_L g3274 ( 
.A1(n_2733),
.A2(n_1645),
.B1(n_1651),
.B2(n_1641),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_SL g3275 ( 
.A(n_2785),
.B(n_1652),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2685),
.B(n_1654),
.Y(n_3276)
);

BUFx6f_ASAP7_75t_L g3277 ( 
.A(n_2414),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2685),
.B(n_1655),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_2396),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2685),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_2632),
.A2(n_1661),
.B1(n_1669),
.B2(n_1668),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_2785),
.B(n_1677),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2486),
.B(n_1679),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2685),
.B(n_1680),
.Y(n_3284)
);

INVx2_ASAP7_75t_SL g3285 ( 
.A(n_2406),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2685),
.Y(n_3286)
);

OR2x2_ASAP7_75t_L g3287 ( 
.A(n_2458),
.B(n_1681),
.Y(n_3287)
);

AOI22xp33_ASAP7_75t_L g3288 ( 
.A1(n_2632),
.A2(n_1682),
.B1(n_1693),
.B2(n_1686),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2685),
.Y(n_3289)
);

AND2x4_ASAP7_75t_L g3290 ( 
.A(n_2685),
.B(n_1164),
.Y(n_3290)
);

BUFx3_ASAP7_75t_L g3291 ( 
.A(n_2534),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2685),
.Y(n_3292)
);

INVx4_ASAP7_75t_L g3293 ( 
.A(n_2459),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2685),
.B(n_1696),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_SL g3295 ( 
.A(n_2785),
.B(n_1700),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_2396),
.Y(n_3296)
);

CKINVDCx20_ASAP7_75t_R g3297 ( 
.A(n_2394),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_2396),
.Y(n_3298)
);

AOI22xp33_ASAP7_75t_SL g3299 ( 
.A1(n_2429),
.A2(n_1701),
.B1(n_1289),
.B2(n_1176),
.Y(n_3299)
);

BUFx6f_ASAP7_75t_L g3300 ( 
.A(n_2414),
.Y(n_3300)
);

NAND2xp33_ASAP7_75t_L g3301 ( 
.A(n_2783),
.B(n_1289),
.Y(n_3301)
);

AND2x2_ASAP7_75t_L g3302 ( 
.A(n_2458),
.B(n_1168),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2685),
.Y(n_3303)
);

OR2x6_ASAP7_75t_L g3304 ( 
.A(n_2770),
.B(n_1138),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_2458),
.B(n_1182),
.Y(n_3305)
);

AOI22xp33_ASAP7_75t_L g3306 ( 
.A1(n_2632),
.A2(n_1290),
.B1(n_1339),
.B2(n_1163),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2685),
.Y(n_3307)
);

BUFx6f_ASAP7_75t_L g3308 ( 
.A(n_2414),
.Y(n_3308)
);

INVx4_ASAP7_75t_L g3309 ( 
.A(n_2459),
.Y(n_3309)
);

BUFx3_ASAP7_75t_L g3310 ( 
.A(n_2534),
.Y(n_3310)
);

NOR2xp33_ASAP7_75t_L g3311 ( 
.A(n_2486),
.B(n_1185),
.Y(n_3311)
);

INVx2_ASAP7_75t_SL g3312 ( 
.A(n_2406),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2685),
.Y(n_3313)
);

AOI22xp5_ASAP7_75t_L g3314 ( 
.A1(n_2727),
.A2(n_1290),
.B1(n_1339),
.B2(n_1163),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_2785),
.B(n_1440),
.Y(n_3315)
);

NOR2x1p5_ASAP7_75t_L g3316 ( 
.A(n_2393),
.B(n_1648),
.Y(n_3316)
);

INVx2_ASAP7_75t_SL g3317 ( 
.A(n_2406),
.Y(n_3317)
);

AND2x2_ASAP7_75t_L g3318 ( 
.A(n_2458),
.B(n_1190),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_2458),
.B(n_1191),
.Y(n_3319)
);

AND2x4_ASAP7_75t_L g3320 ( 
.A(n_2685),
.B(n_1193),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2685),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2685),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_SL g3323 ( 
.A(n_2785),
.B(n_1440),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_2785),
.B(n_1684),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2685),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_2458),
.B(n_1208),
.Y(n_3326)
);

INVx1_ASAP7_75t_SL g3327 ( 
.A(n_2407),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2396),
.Y(n_3328)
);

OR2x2_ASAP7_75t_L g3329 ( 
.A(n_2458),
.B(n_1224),
.Y(n_3329)
);

CKINVDCx5p33_ASAP7_75t_R g3330 ( 
.A(n_2393),
.Y(n_3330)
);

INVx2_ASAP7_75t_SL g3331 ( 
.A(n_2406),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_SL g3332 ( 
.A(n_2785),
.B(n_1684),
.Y(n_3332)
);

BUFx6f_ASAP7_75t_L g3333 ( 
.A(n_2414),
.Y(n_3333)
);

BUFx3_ASAP7_75t_L g3334 ( 
.A(n_2534),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2685),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2685),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_SL g3337 ( 
.A(n_2785),
.B(n_1187),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2685),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_SL g3339 ( 
.A(n_2785),
.B(n_1231),
.Y(n_3339)
);

AOI22xp5_ASAP7_75t_L g3340 ( 
.A1(n_2727),
.A2(n_1235),
.B1(n_1242),
.B2(n_1232),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_2685),
.Y(n_3341)
);

INVx3_ASAP7_75t_L g3342 ( 
.A(n_2750),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_2785),
.B(n_1276),
.Y(n_3343)
);

INVx2_ASAP7_75t_SL g3344 ( 
.A(n_2406),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_L g3345 ( 
.A(n_2486),
.B(n_1245),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_2396),
.Y(n_3346)
);

NAND2x1p5_ASAP7_75t_L g3347 ( 
.A(n_2572),
.B(n_1258),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_2685),
.B(n_1251),
.Y(n_3348)
);

OR2x6_ASAP7_75t_L g3349 ( 
.A(n_2770),
.B(n_1276),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2685),
.B(n_1262),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_2396),
.Y(n_3351)
);

INVx4_ASAP7_75t_L g3352 ( 
.A(n_2459),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_2458),
.B(n_1264),
.Y(n_3353)
);

NAND3xp33_ASAP7_75t_SL g3354 ( 
.A(n_2429),
.B(n_1270),
.C(n_1266),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_L g3355 ( 
.A(n_2486),
.B(n_1273),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_L g3356 ( 
.A1(n_2632),
.A2(n_1291),
.B1(n_1300),
.B2(n_1279),
.Y(n_3356)
);

NOR2xp33_ASAP7_75t_L g3357 ( 
.A(n_2486),
.B(n_1303),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_SL g3358 ( 
.A(n_2785),
.B(n_1294),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2396),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_2396),
.Y(n_3360)
);

INVx4_ASAP7_75t_L g3361 ( 
.A(n_2459),
.Y(n_3361)
);

AND2x2_ASAP7_75t_L g3362 ( 
.A(n_2458),
.B(n_1306),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_2458),
.B(n_1308),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2685),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2685),
.Y(n_3365)
);

INVx4_ASAP7_75t_L g3366 ( 
.A(n_2459),
.Y(n_3366)
);

BUFx3_ASAP7_75t_L g3367 ( 
.A(n_2534),
.Y(n_3367)
);

BUFx2_ASAP7_75t_L g3368 ( 
.A(n_2422),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_2458),
.B(n_1321),
.Y(n_3369)
);

INVx4_ASAP7_75t_L g3370 ( 
.A(n_2459),
.Y(n_3370)
);

AND2x4_ASAP7_75t_L g3371 ( 
.A(n_2685),
.B(n_1325),
.Y(n_3371)
);

INVxp33_ASAP7_75t_L g3372 ( 
.A(n_2484),
.Y(n_3372)
);

BUFx10_ASAP7_75t_L g3373 ( 
.A(n_2393),
.Y(n_3373)
);

CKINVDCx20_ASAP7_75t_R g3374 ( 
.A(n_2394),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_2632),
.A2(n_1327),
.B1(n_1334),
.B2(n_1326),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2685),
.Y(n_3376)
);

INVx5_ASAP7_75t_L g3377 ( 
.A(n_2783),
.Y(n_3377)
);

OAI21xp33_ASAP7_75t_SL g3378 ( 
.A1(n_2418),
.A2(n_1301),
.B(n_1294),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_2685),
.B(n_1335),
.Y(n_3379)
);

INVx2_ASAP7_75t_SL g3380 ( 
.A(n_2406),
.Y(n_3380)
);

INVx3_ASAP7_75t_L g3381 ( 
.A(n_2750),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_2486),
.B(n_1345),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2685),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_2396),
.Y(n_3384)
);

INVx4_ASAP7_75t_SL g3385 ( 
.A(n_2783),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_2458),
.B(n_1347),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2685),
.Y(n_3387)
);

INVx2_ASAP7_75t_SL g3388 ( 
.A(n_2406),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_2685),
.B(n_1349),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_2396),
.Y(n_3390)
);

BUFx6f_ASAP7_75t_L g3391 ( 
.A(n_2414),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_2396),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_2785),
.B(n_1672),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_L g3394 ( 
.A(n_2486),
.B(n_1361),
.Y(n_3394)
);

INVx2_ASAP7_75t_SL g3395 ( 
.A(n_2406),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2685),
.Y(n_3396)
);

NOR2xp33_ASAP7_75t_L g3397 ( 
.A(n_2486),
.B(n_1363),
.Y(n_3397)
);

NAND3xp33_ASAP7_75t_L g3398 ( 
.A(n_2702),
.B(n_1502),
.C(n_1444),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_2396),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2685),
.Y(n_3400)
);

NAND3xp33_ASAP7_75t_L g3401 ( 
.A(n_2702),
.B(n_1502),
.C(n_1444),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_2685),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2685),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2685),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_SL g3405 ( 
.A(n_2785),
.B(n_1301),
.Y(n_3405)
);

INVxp67_ASAP7_75t_L g3406 ( 
.A(n_2401),
.Y(n_3406)
);

INVxp33_ASAP7_75t_SL g3407 ( 
.A(n_2429),
.Y(n_3407)
);

BUFx3_ASAP7_75t_L g3408 ( 
.A(n_2534),
.Y(n_3408)
);

INVx1_ASAP7_75t_SL g3409 ( 
.A(n_2407),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_2396),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_2685),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_2486),
.B(n_1364),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_2458),
.B(n_1365),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_2486),
.B(n_1370),
.Y(n_3414)
);

BUFx6f_ASAP7_75t_L g3415 ( 
.A(n_2414),
.Y(n_3415)
);

OAI22xp33_ASAP7_75t_L g3416 ( 
.A1(n_2733),
.A2(n_1374),
.B1(n_1386),
.B2(n_1372),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_2396),
.Y(n_3417)
);

INVxp33_ASAP7_75t_L g3418 ( 
.A(n_2484),
.Y(n_3418)
);

INVx3_ASAP7_75t_L g3419 ( 
.A(n_2750),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2685),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2685),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2685),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_2396),
.Y(n_3423)
);

BUFx6f_ASAP7_75t_L g3424 ( 
.A(n_2414),
.Y(n_3424)
);

INVx1_ASAP7_75t_SL g3425 ( 
.A(n_2407),
.Y(n_3425)
);

AOI22xp33_ASAP7_75t_L g3426 ( 
.A1(n_2632),
.A2(n_1388),
.B1(n_1392),
.B2(n_1387),
.Y(n_3426)
);

INVx4_ASAP7_75t_L g3427 ( 
.A(n_2459),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_SL g3428 ( 
.A(n_2785),
.B(n_1672),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_2396),
.Y(n_3429)
);

INVx6_ASAP7_75t_L g3430 ( 
.A(n_2779),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_2685),
.Y(n_3431)
);

NAND2xp33_ASAP7_75t_SL g3432 ( 
.A(n_2629),
.B(n_1312),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_2396),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_2396),
.Y(n_3434)
);

BUFx6f_ASAP7_75t_L g3435 ( 
.A(n_2414),
.Y(n_3435)
);

INVxp67_ASAP7_75t_SL g3436 ( 
.A(n_2407),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_2685),
.B(n_1394),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_SL g3438 ( 
.A(n_2572),
.B(n_1312),
.Y(n_3438)
);

BUFx10_ASAP7_75t_L g3439 ( 
.A(n_2393),
.Y(n_3439)
);

INVx1_ASAP7_75t_SL g3440 ( 
.A(n_2407),
.Y(n_3440)
);

AND2x6_ASAP7_75t_L g3441 ( 
.A(n_2445),
.B(n_1444),
.Y(n_3441)
);

INVx4_ASAP7_75t_L g3442 ( 
.A(n_2459),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_SL g3443 ( 
.A(n_2785),
.B(n_1355),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_2685),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_SL g3445 ( 
.A(n_2785),
.B(n_1355),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3234),
.B(n_1396),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3444),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_2892),
.B(n_1397),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_2804),
.B(n_1444),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3208),
.B(n_1398),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3213),
.Y(n_3451)
);

OAI22xp5_ASAP7_75t_L g3452 ( 
.A1(n_2915),
.A2(n_1411),
.B1(n_1415),
.B2(n_1399),
.Y(n_3452)
);

INVx2_ASAP7_75t_SL g3453 ( 
.A(n_2931),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3218),
.B(n_1408),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3431),
.Y(n_3455)
);

NOR2xp33_ASAP7_75t_SL g3456 ( 
.A(n_2854),
.B(n_1399),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3226),
.Y(n_3457)
);

INVxp67_ASAP7_75t_SL g3458 ( 
.A(n_3031),
.Y(n_3458)
);

OR2x2_ASAP7_75t_L g3459 ( 
.A(n_2789),
.B(n_1706),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3230),
.B(n_1409),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3233),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3239),
.B(n_1414),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3249),
.B(n_3257),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3265),
.B(n_1434),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_2940),
.B(n_3407),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_SL g3466 ( 
.A(n_2940),
.B(n_1502),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3271),
.Y(n_3467)
);

NOR3xp33_ASAP7_75t_L g3468 ( 
.A(n_2810),
.B(n_1439),
.C(n_1436),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3280),
.B(n_1452),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3286),
.B(n_1458),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3289),
.Y(n_3471)
);

NOR2xp33_ASAP7_75t_L g3472 ( 
.A(n_3372),
.B(n_3418),
.Y(n_3472)
);

NAND2xp33_ASAP7_75t_L g3473 ( 
.A(n_2854),
.B(n_1502),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3292),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3303),
.Y(n_3475)
);

CKINVDCx5p33_ASAP7_75t_R g3476 ( 
.A(n_2787),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3307),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_2892),
.B(n_1460),
.Y(n_3478)
);

AOI22xp33_ASAP7_75t_SL g3479 ( 
.A1(n_2837),
.A2(n_3092),
.B1(n_3062),
.B2(n_2915),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_SL g3480 ( 
.A(n_2789),
.B(n_1587),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3313),
.Y(n_3481)
);

NOR2xp67_ASAP7_75t_L g3482 ( 
.A(n_2931),
.B(n_266),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_SL g3483 ( 
.A(n_3074),
.B(n_1587),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3321),
.B(n_1463),
.Y(n_3484)
);

NAND2x1_ASAP7_75t_L g3485 ( 
.A(n_3246),
.B(n_3441),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_SL g3486 ( 
.A(n_3074),
.B(n_1587),
.Y(n_3486)
);

INVx5_ASAP7_75t_L g3487 ( 
.A(n_3174),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3322),
.B(n_1467),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3325),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3335),
.B(n_1487),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3336),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3338),
.B(n_1489),
.Y(n_3492)
);

OAI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_2993),
.A2(n_1496),
.B1(n_1497),
.B2(n_1492),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3341),
.Y(n_3494)
);

INVx2_ASAP7_75t_SL g3495 ( 
.A(n_2931),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3126),
.B(n_2947),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3364),
.B(n_3365),
.Y(n_3497)
);

O2A1O1Ixp33_ASAP7_75t_L g3498 ( 
.A1(n_2836),
.A2(n_1504),
.B(n_1507),
.C(n_1499),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3376),
.B(n_1510),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_2837),
.B(n_1521),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_L g3501 ( 
.A(n_2831),
.B(n_1527),
.Y(n_3501)
);

OAI22xp33_ASAP7_75t_L g3502 ( 
.A1(n_2993),
.A2(n_1540),
.B1(n_1544),
.B2(n_1529),
.Y(n_3502)
);

INVx2_ASAP7_75t_SL g3503 ( 
.A(n_3172),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3383),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3387),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_2857),
.B(n_1549),
.Y(n_3506)
);

AO22x2_ASAP7_75t_L g3507 ( 
.A1(n_3138),
.A2(n_1415),
.B1(n_1471),
.B2(n_1411),
.Y(n_3507)
);

INVx2_ASAP7_75t_SL g3508 ( 
.A(n_3172),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_SL g3509 ( 
.A(n_3126),
.B(n_1587),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3396),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3400),
.B(n_1551),
.Y(n_3511)
);

AND2x6_ASAP7_75t_SL g3512 ( 
.A(n_3154),
.B(n_1556),
.Y(n_3512)
);

OAI221xp5_ASAP7_75t_L g3513 ( 
.A1(n_3306),
.A2(n_2794),
.B1(n_3375),
.B2(n_3426),
.C(n_3356),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3402),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3403),
.Y(n_3515)
);

AND2x2_ASAP7_75t_SL g3516 ( 
.A(n_3106),
.B(n_1626),
.Y(n_3516)
);

AOI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_2791),
.A2(n_1626),
.B1(n_1481),
.B2(n_1484),
.Y(n_3517)
);

AOI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_3209),
.A2(n_1481),
.B(n_1471),
.Y(n_3518)
);

AOI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_3354),
.A2(n_1561),
.B1(n_1567),
.B2(n_1559),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_L g3520 ( 
.A(n_3221),
.B(n_1572),
.Y(n_3520)
);

NAND2xp33_ASAP7_75t_SL g3521 ( 
.A(n_3006),
.B(n_1484),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3404),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_SL g3523 ( 
.A(n_2947),
.B(n_1626),
.Y(n_3523)
);

INVxp67_ASAP7_75t_L g3524 ( 
.A(n_2866),
.Y(n_3524)
);

INVxp67_ASAP7_75t_L g3525 ( 
.A(n_2879),
.Y(n_3525)
);

AOI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3045),
.A2(n_1576),
.B1(n_1577),
.B2(n_1573),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_3411),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3420),
.B(n_1578),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_SL g3529 ( 
.A(n_2788),
.B(n_3327),
.Y(n_3529)
);

AOI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_3125),
.A2(n_1580),
.B1(n_1581),
.B2(n_1579),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3421),
.Y(n_3531)
);

NOR2xp33_ASAP7_75t_L g3532 ( 
.A(n_3222),
.B(n_1582),
.Y(n_3532)
);

BUFx6f_ASAP7_75t_L g3533 ( 
.A(n_2801),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_SL g3534 ( 
.A(n_2788),
.B(n_3327),
.Y(n_3534)
);

NOR2xp33_ASAP7_75t_L g3535 ( 
.A(n_3223),
.B(n_1584),
.Y(n_3535)
);

NOR3xp33_ASAP7_75t_L g3536 ( 
.A(n_3250),
.B(n_3432),
.C(n_3345),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_2814),
.B(n_1585),
.Y(n_3537)
);

NAND3xp33_ASAP7_75t_L g3538 ( 
.A(n_3103),
.B(n_1626),
.C(n_1603),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3422),
.B(n_1599),
.Y(n_3539)
);

OAI22xp5_ASAP7_75t_L g3540 ( 
.A1(n_3024),
.A2(n_1518),
.B1(n_1545),
.B2(n_1514),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_2917),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3311),
.B(n_1604),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_2921),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3240),
.B(n_3243),
.Y(n_3544)
);

NOR2xp67_ASAP7_75t_L g3545 ( 
.A(n_3057),
.B(n_266),
.Y(n_3545)
);

BUFx3_ASAP7_75t_L g3546 ( 
.A(n_3174),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3355),
.B(n_1610),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3357),
.B(n_1611),
.Y(n_3548)
);

AND2x4_ASAP7_75t_L g3549 ( 
.A(n_2876),
.B(n_1514),
.Y(n_3549)
);

NOR2xp33_ASAP7_75t_L g3550 ( 
.A(n_3256),
.B(n_1612),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3382),
.B(n_1617),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_3409),
.B(n_1518),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_2928),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3394),
.B(n_1624),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_3409),
.B(n_1545),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_2932),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_2790),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_3425),
.B(n_1557),
.Y(n_3558)
);

INVxp67_ASAP7_75t_L g3559 ( 
.A(n_2880),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3397),
.B(n_1636),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3412),
.B(n_1638),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3266),
.B(n_1644),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3414),
.B(n_1649),
.Y(n_3563)
);

INVx2_ASAP7_75t_SL g3564 ( 
.A(n_3172),
.Y(n_3564)
);

OAI22xp33_ASAP7_75t_L g3565 ( 
.A1(n_3024),
.A2(n_1670),
.B1(n_1671),
.B2(n_1653),
.Y(n_3565)
);

OAI22xp33_ASAP7_75t_L g3566 ( 
.A1(n_2893),
.A2(n_1685),
.B1(n_1688),
.B2(n_1673),
.Y(n_3566)
);

NOR2xp33_ASAP7_75t_L g3567 ( 
.A(n_3283),
.B(n_1692),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_2796),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3340),
.B(n_1697),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_2792),
.Y(n_3570)
);

INVx8_ASAP7_75t_L g3571 ( 
.A(n_3057),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3340),
.B(n_1713),
.Y(n_3572)
);

BUFx6f_ASAP7_75t_SL g3573 ( 
.A(n_2848),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_L g3574 ( 
.A(n_3014),
.B(n_1557),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3242),
.B(n_1586),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3242),
.B(n_1586),
.Y(n_3576)
);

NAND2xp33_ASAP7_75t_L g3577 ( 
.A(n_2854),
.B(n_1613),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3290),
.B(n_1613),
.Y(n_3578)
);

CKINVDCx5p33_ASAP7_75t_R g3579 ( 
.A(n_2911),
.Y(n_3579)
);

INVx4_ASAP7_75t_L g3580 ( 
.A(n_3174),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3290),
.B(n_1630),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3320),
.B(n_1630),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3320),
.B(n_1646),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_2793),
.Y(n_3584)
);

BUFx6f_ASAP7_75t_L g3585 ( 
.A(n_2801),
.Y(n_3585)
);

INVx2_ASAP7_75t_SL g3586 ( 
.A(n_3185),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_2806),
.Y(n_3587)
);

HB1xp67_ASAP7_75t_L g3588 ( 
.A(n_3304),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_2799),
.Y(n_3589)
);

NOR2xp33_ASAP7_75t_L g3590 ( 
.A(n_3025),
.B(n_1646),
.Y(n_3590)
);

NAND2xp5_ASAP7_75t_SL g3591 ( 
.A(n_3425),
.B(n_267),
.Y(n_3591)
);

NOR2xp33_ASAP7_75t_L g3592 ( 
.A(n_2856),
.B(n_267),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3437),
.B(n_267),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_2816),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3437),
.B(n_268),
.Y(n_3595)
);

NOR2xp33_ASAP7_75t_L g3596 ( 
.A(n_3214),
.B(n_268),
.Y(n_3596)
);

NAND2x1_ASAP7_75t_L g3597 ( 
.A(n_3246),
.B(n_268),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3371),
.B(n_269),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_2820),
.B(n_269),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_2812),
.Y(n_3600)
);

INVx2_ASAP7_75t_SL g3601 ( 
.A(n_3185),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_2823),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_SL g3603 ( 
.A(n_3440),
.B(n_269),
.Y(n_3603)
);

AND2x2_ASAP7_75t_L g3604 ( 
.A(n_2948),
.B(n_270),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3371),
.B(n_270),
.Y(n_3605)
);

NOR2xp33_ASAP7_75t_L g3606 ( 
.A(n_3274),
.B(n_2872),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_2825),
.Y(n_3607)
);

AOI221xp5_ASAP7_75t_L g3608 ( 
.A1(n_3416),
.A2(n_272),
.B1(n_273),
.B2(n_271),
.C(n_270),
.Y(n_3608)
);

BUFx2_ASAP7_75t_L g3609 ( 
.A(n_2968),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_2835),
.Y(n_3610)
);

NOR2xp67_ASAP7_75t_L g3611 ( 
.A(n_3057),
.B(n_271),
.Y(n_3611)
);

CKINVDCx5p33_ASAP7_75t_R g3612 ( 
.A(n_2999),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_2850),
.B(n_271),
.Y(n_3613)
);

NOR2xp33_ASAP7_75t_L g3614 ( 
.A(n_2959),
.B(n_272),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_2850),
.B(n_273),
.Y(n_3615)
);

BUFx6f_ASAP7_75t_L g3616 ( 
.A(n_2801),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_2840),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_2845),
.Y(n_3618)
);

AOI22xp33_ASAP7_75t_L g3619 ( 
.A1(n_3062),
.A2(n_274),
.B1(n_275),
.B2(n_273),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3210),
.B(n_274),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_L g3621 ( 
.A(n_3085),
.B(n_275),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_2853),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_2952),
.B(n_276),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_2859),
.Y(n_3624)
);

AND2x4_ASAP7_75t_L g3625 ( 
.A(n_2876),
.B(n_276),
.Y(n_3625)
);

INVx3_ASAP7_75t_L g3626 ( 
.A(n_3212),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_2819),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_2865),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_2847),
.Y(n_3629)
);

NOR2xp33_ASAP7_75t_L g3630 ( 
.A(n_2945),
.B(n_276),
.Y(n_3630)
);

BUFx6f_ASAP7_75t_L g3631 ( 
.A(n_2813),
.Y(n_3631)
);

NOR2xp67_ASAP7_75t_SL g3632 ( 
.A(n_2832),
.B(n_277),
.Y(n_3632)
);

CKINVDCx5p33_ASAP7_75t_R g3633 ( 
.A(n_3077),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3210),
.B(n_278),
.Y(n_3634)
);

AOI22xp5_ASAP7_75t_L g3635 ( 
.A1(n_2888),
.A2(n_279),
.B1(n_280),
.B2(n_278),
.Y(n_3635)
);

NAND3xp33_ASAP7_75t_L g3636 ( 
.A(n_3103),
.B(n_280),
.C(n_279),
.Y(n_3636)
);

NOR2xp33_ASAP7_75t_L g3637 ( 
.A(n_3184),
.B(n_280),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_2873),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3219),
.B(n_281),
.Y(n_3639)
);

NAND3xp33_ASAP7_75t_L g3640 ( 
.A(n_3398),
.B(n_282),
.C(n_281),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_3219),
.B(n_282),
.Y(n_3641)
);

NOR2xp33_ASAP7_75t_SL g3642 ( 
.A(n_3212),
.B(n_282),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_2860),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3207),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_2890),
.B(n_3220),
.Y(n_3645)
);

INVxp67_ASAP7_75t_L g3646 ( 
.A(n_3304),
.Y(n_3646)
);

NOR2x1p5_ASAP7_75t_L g3647 ( 
.A(n_2809),
.B(n_2953),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_2890),
.B(n_283),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3245),
.B(n_283),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3220),
.B(n_283),
.Y(n_3650)
);

AOI22xp33_ASAP7_75t_L g3651 ( 
.A1(n_3092),
.A2(n_285),
.B1(n_286),
.B2(n_284),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_L g3652 ( 
.A(n_3184),
.B(n_284),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3238),
.B(n_284),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3238),
.B(n_285),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3232),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3244),
.B(n_285),
.Y(n_3656)
);

NOR2xp33_ASAP7_75t_L g3657 ( 
.A(n_3029),
.B(n_286),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3244),
.B(n_286),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3247),
.B(n_287),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_2883),
.Y(n_3660)
);

INVxp67_ASAP7_75t_SL g3661 ( 
.A(n_3030),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3440),
.B(n_287),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_2887),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3253),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_2891),
.Y(n_3665)
);

CKINVDCx5p33_ASAP7_75t_R g3666 ( 
.A(n_3297),
.Y(n_3666)
);

NAND2xp33_ASAP7_75t_L g3667 ( 
.A(n_3212),
.B(n_287),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3247),
.B(n_3252),
.Y(n_3668)
);

NOR2xp33_ASAP7_75t_L g3669 ( 
.A(n_3093),
.B(n_288),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_SL g3670 ( 
.A(n_3096),
.B(n_2933),
.Y(n_3670)
);

NOR2xp33_ASAP7_75t_L g3671 ( 
.A(n_2821),
.B(n_288),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3252),
.B(n_288),
.Y(n_3672)
);

OR2x2_ASAP7_75t_L g3673 ( 
.A(n_2874),
.B(n_289),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3261),
.B(n_289),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_SL g3675 ( 
.A(n_3096),
.B(n_2933),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3261),
.B(n_289),
.Y(n_3676)
);

O2A1O1Ixp33_ASAP7_75t_L g3677 ( 
.A1(n_2836),
.A2(n_3269),
.B(n_3276),
.C(n_3273),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3260),
.Y(n_3678)
);

INVx2_ASAP7_75t_SL g3679 ( 
.A(n_3185),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3269),
.B(n_290),
.Y(n_3680)
);

NOR2xp67_ASAP7_75t_SL g3681 ( 
.A(n_3377),
.B(n_290),
.Y(n_3681)
);

NAND2xp33_ASAP7_75t_L g3682 ( 
.A(n_3377),
.B(n_290),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3273),
.B(n_291),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3279),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3276),
.B(n_291),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3278),
.B(n_292),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_2898),
.Y(n_3687)
);

NOR2xp33_ASAP7_75t_L g3688 ( 
.A(n_3061),
.B(n_292),
.Y(n_3688)
);

O2A1O1Ixp33_ASAP7_75t_L g3689 ( 
.A1(n_3278),
.A2(n_3284),
.B(n_3294),
.C(n_3027),
.Y(n_3689)
);

HB1xp67_ASAP7_75t_L g3690 ( 
.A(n_3304),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_SL g3691 ( 
.A(n_2987),
.B(n_293),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3296),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3284),
.B(n_293),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3294),
.B(n_293),
.Y(n_3694)
);

INVx2_ASAP7_75t_SL g3695 ( 
.A(n_3183),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_2802),
.B(n_3368),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_2905),
.B(n_294),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_2908),
.B(n_294),
.Y(n_3698)
);

BUFx6f_ASAP7_75t_L g3699 ( 
.A(n_2813),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_2919),
.B(n_294),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_SL g3701 ( 
.A(n_3377),
.B(n_295),
.Y(n_3701)
);

INVxp67_ASAP7_75t_SL g3702 ( 
.A(n_2870),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3298),
.Y(n_3703)
);

NOR3xp33_ASAP7_75t_L g3704 ( 
.A(n_2964),
.B(n_296),
.C(n_295),
.Y(n_3704)
);

AOI22xp33_ASAP7_75t_L g3705 ( 
.A1(n_3147),
.A2(n_296),
.B1(n_297),
.B2(n_295),
.Y(n_3705)
);

INVx2_ASAP7_75t_SL g3706 ( 
.A(n_3183),
.Y(n_3706)
);

INVx4_ASAP7_75t_L g3707 ( 
.A(n_3183),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3328),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_2922),
.Y(n_3709)
);

NAND3xp33_ASAP7_75t_L g3710 ( 
.A(n_3398),
.B(n_297),
.C(n_296),
.Y(n_3710)
);

NOR2xp67_ASAP7_75t_L g3711 ( 
.A(n_2982),
.B(n_297),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_2925),
.B(n_298),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3302),
.B(n_298),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_2981),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3346),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3351),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3305),
.B(n_298),
.Y(n_3717)
);

INVx2_ASAP7_75t_SL g3718 ( 
.A(n_3193),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_L g3719 ( 
.A1(n_3147),
.A2(n_300),
.B1(n_301),
.B2(n_299),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_SL g3720 ( 
.A(n_2987),
.B(n_3438),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3318),
.B(n_299),
.Y(n_3721)
);

NOR2xp33_ASAP7_75t_L g3722 ( 
.A(n_2912),
.B(n_299),
.Y(n_3722)
);

BUFx6f_ASAP7_75t_L g3723 ( 
.A(n_2813),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_3319),
.B(n_300),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3326),
.B(n_300),
.Y(n_3725)
);

O2A1O1Ixp5_ASAP7_75t_L g3726 ( 
.A1(n_2808),
.A2(n_302),
.B(n_303),
.C(n_301),
.Y(n_3726)
);

NAND2xp33_ASAP7_75t_L g3727 ( 
.A(n_3113),
.B(n_301),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3353),
.B(n_302),
.Y(n_3728)
);

BUFx6f_ASAP7_75t_SL g3729 ( 
.A(n_2848),
.Y(n_3729)
);

BUFx24_ASAP7_75t_SL g3730 ( 
.A(n_3134),
.Y(n_3730)
);

INVx4_ASAP7_75t_L g3731 ( 
.A(n_3193),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_2808),
.A2(n_304),
.B1(n_305),
.B2(n_303),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_2985),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3359),
.Y(n_3734)
);

NAND2xp33_ASAP7_75t_L g3735 ( 
.A(n_3113),
.B(n_303),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3362),
.B(n_304),
.Y(n_3736)
);

NOR2xp33_ASAP7_75t_L g3737 ( 
.A(n_3035),
.B(n_304),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3007),
.Y(n_3738)
);

OAI22xp5_ASAP7_75t_L g3739 ( 
.A1(n_2829),
.A2(n_306),
.B1(n_307),
.B2(n_305),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3363),
.B(n_3369),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3258),
.B(n_305),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3386),
.B(n_306),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3413),
.B(n_307),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3314),
.B(n_307),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_SL g3745 ( 
.A(n_3438),
.B(n_308),
.Y(n_3745)
);

NOR2xp33_ASAP7_75t_L g3746 ( 
.A(n_3166),
.B(n_308),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3360),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3009),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_SL g3749 ( 
.A(n_3042),
.B(n_308),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3314),
.B(n_309),
.Y(n_3750)
);

INVx3_ASAP7_75t_L g3751 ( 
.A(n_3089),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3013),
.Y(n_3752)
);

AND2x4_ASAP7_75t_SL g3753 ( 
.A(n_2926),
.B(n_309),
.Y(n_3753)
);

AOI22xp33_ASAP7_75t_L g3754 ( 
.A1(n_3236),
.A2(n_310),
.B1(n_311),
.B2(n_309),
.Y(n_3754)
);

INVx8_ASAP7_75t_L g3755 ( 
.A(n_3349),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3384),
.Y(n_3756)
);

OR2x6_ASAP7_75t_L g3757 ( 
.A(n_3349),
.B(n_310),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_SL g3758 ( 
.A(n_2939),
.B(n_310),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3018),
.Y(n_3759)
);

INVxp67_ASAP7_75t_L g3760 ( 
.A(n_3349),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3075),
.Y(n_3761)
);

INVx3_ASAP7_75t_L g3762 ( 
.A(n_3089),
.Y(n_3762)
);

NOR2xp33_ASAP7_75t_L g3763 ( 
.A(n_3166),
.B(n_311),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_3149),
.B(n_312),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_SL g3765 ( 
.A(n_3047),
.B(n_312),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3078),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_2829),
.B(n_312),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3390),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3348),
.B(n_313),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3348),
.B(n_313),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_2934),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_2935),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3392),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3350),
.B(n_313),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3399),
.Y(n_3775)
);

BUFx2_ASAP7_75t_L g3776 ( 
.A(n_3374),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_2946),
.Y(n_3777)
);

AOI22xp5_ASAP7_75t_L g3778 ( 
.A1(n_2957),
.A2(n_315),
.B1(n_316),
.B2(n_314),
.Y(n_3778)
);

NOR2xp33_ASAP7_75t_L g3779 ( 
.A(n_3169),
.B(n_314),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3350),
.B(n_315),
.Y(n_3780)
);

AND2x4_ASAP7_75t_L g3781 ( 
.A(n_3231),
.B(n_315),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3379),
.B(n_316),
.Y(n_3782)
);

OR2x6_ASAP7_75t_L g3783 ( 
.A(n_2982),
.B(n_316),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3379),
.B(n_317),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3005),
.B(n_317),
.Y(n_3785)
);

INVxp33_ASAP7_75t_L g3786 ( 
.A(n_3164),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_SL g3787 ( 
.A(n_2849),
.B(n_317),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3410),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3389),
.B(n_318),
.Y(n_3789)
);

INVxp67_ASAP7_75t_L g3790 ( 
.A(n_2849),
.Y(n_3790)
);

NOR2xp33_ASAP7_75t_L g3791 ( 
.A(n_3067),
.B(n_318),
.Y(n_3791)
);

NOR2xp33_ASAP7_75t_L g3792 ( 
.A(n_3176),
.B(n_319),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_SL g3793 ( 
.A(n_2980),
.B(n_319),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_2956),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_2966),
.B(n_320),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3417),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3389),
.B(n_3215),
.Y(n_3797)
);

BUFx6f_ASAP7_75t_L g3798 ( 
.A(n_2868),
.Y(n_3798)
);

NOR2xp67_ASAP7_75t_L g3799 ( 
.A(n_2824),
.B(n_320),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_2979),
.B(n_321),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_3215),
.B(n_321),
.Y(n_3801)
);

AOI22xp5_ASAP7_75t_L g3802 ( 
.A1(n_2930),
.A2(n_323),
.B1(n_324),
.B2(n_322),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_2962),
.Y(n_3803)
);

INVx3_ASAP7_75t_L g3804 ( 
.A(n_3089),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_2826),
.B(n_322),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3268),
.B(n_323),
.Y(n_3806)
);

NOR2xp33_ASAP7_75t_L g3807 ( 
.A(n_3151),
.B(n_323),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_2826),
.B(n_324),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3170),
.B(n_324),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_2811),
.A2(n_327),
.B(n_325),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3020),
.Y(n_3811)
);

NOR2xp33_ASAP7_75t_L g3812 ( 
.A(n_3102),
.B(n_327),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_SL g3813 ( 
.A(n_3170),
.B(n_3019),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3021),
.Y(n_3814)
);

AOI22xp5_ASAP7_75t_L g3815 ( 
.A1(n_3134),
.A2(n_328),
.B1(n_329),
.B2(n_327),
.Y(n_3815)
);

OAI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3378),
.A2(n_0),
.B(n_1),
.Y(n_3816)
);

AOI22xp5_ASAP7_75t_L g3817 ( 
.A1(n_3119),
.A2(n_329),
.B1(n_330),
.B2(n_328),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_2811),
.A2(n_329),
.B(n_328),
.Y(n_3818)
);

AOI22xp33_ASAP7_75t_L g3819 ( 
.A1(n_3255),
.A2(n_331),
.B1(n_332),
.B2(n_330),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3105),
.B(n_3138),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_SL g3821 ( 
.A(n_2897),
.B(n_330),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_L g3822 ( 
.A(n_3114),
.B(n_332),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_2974),
.B(n_332),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3231),
.B(n_333),
.Y(n_3824)
);

AOI22xp5_ASAP7_75t_L g3825 ( 
.A1(n_3181),
.A2(n_334),
.B1(n_335),
.B2(n_333),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_2974),
.B(n_334),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3032),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3423),
.Y(n_3828)
);

NOR2xp33_ASAP7_75t_L g3829 ( 
.A(n_2827),
.B(n_334),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_SL g3830 ( 
.A(n_3385),
.B(n_335),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_2871),
.B(n_335),
.Y(n_3831)
);

O2A1O1Ixp5_ASAP7_75t_L g3832 ( 
.A1(n_3401),
.A2(n_337),
.B(n_338),
.C(n_336),
.Y(n_3832)
);

INVx3_ASAP7_75t_L g3833 ( 
.A(n_2901),
.Y(n_3833)
);

BUFx5_ASAP7_75t_L g3834 ( 
.A(n_3246),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3038),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_2871),
.B(n_336),
.Y(n_3836)
);

NOR2xp33_ASAP7_75t_L g3837 ( 
.A(n_2842),
.B(n_337),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_2882),
.B(n_337),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3039),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3429),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_2882),
.B(n_338),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_2889),
.B(n_338),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_2889),
.B(n_340),
.Y(n_3843)
);

NAND2xp5_ASAP7_75t_L g3844 ( 
.A(n_2894),
.B(n_340),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_2894),
.B(n_340),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_2899),
.B(n_341),
.Y(n_3846)
);

INVx2_ASAP7_75t_L g3847 ( 
.A(n_3433),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3434),
.Y(n_3848)
);

BUFx6f_ASAP7_75t_L g3849 ( 
.A(n_2868),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_2899),
.B(n_341),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_3385),
.B(n_341),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_SL g3852 ( 
.A(n_3131),
.B(n_342),
.Y(n_3852)
);

INVxp67_ASAP7_75t_SL g3853 ( 
.A(n_3406),
.Y(n_3853)
);

AOI22xp5_ASAP7_75t_L g3854 ( 
.A1(n_2978),
.A2(n_343),
.B1(n_344),
.B2(n_342),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_2967),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_2902),
.B(n_342),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_SL g3857 ( 
.A(n_3064),
.B(n_343),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_2902),
.B(n_344),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3086),
.Y(n_3859)
);

AO22x2_ASAP7_75t_L g3860 ( 
.A1(n_3401),
.A2(n_346),
.B1(n_347),
.B2(n_345),
.Y(n_3860)
);

AOI22xp33_ASAP7_75t_L g3861 ( 
.A1(n_3262),
.A2(n_346),
.B1(n_347),
.B2(n_345),
.Y(n_3861)
);

NOR2xp33_ASAP7_75t_L g3862 ( 
.A(n_2903),
.B(n_346),
.Y(n_3862)
);

INVxp67_ASAP7_75t_SL g3863 ( 
.A(n_2961),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_2969),
.Y(n_3864)
);

CKINVDCx5p33_ASAP7_75t_R g3865 ( 
.A(n_3017),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3084),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3064),
.B(n_347),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_2913),
.B(n_348),
.Y(n_3868)
);

NOR2x1p5_ASAP7_75t_L g3869 ( 
.A(n_3066),
.B(n_348),
.Y(n_3869)
);

AOI22xp33_ASAP7_75t_L g3870 ( 
.A1(n_3281),
.A2(n_349),
.B1(n_350),
.B2(n_348),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_2970),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_2971),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_2913),
.B(n_349),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_2976),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_2923),
.B(n_349),
.Y(n_3875)
);

INVxp67_ASAP7_75t_L g3876 ( 
.A(n_3211),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_2973),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_L g3878 ( 
.A(n_2923),
.B(n_350),
.Y(n_3878)
);

OR2x6_ASAP7_75t_L g3879 ( 
.A(n_3430),
.B(n_351),
.Y(n_3879)
);

OAI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3211),
.A2(n_352),
.B1(n_353),
.B2(n_351),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_2963),
.B(n_2807),
.Y(n_3881)
);

CKINVDCx16_ASAP7_75t_R g3882 ( 
.A(n_3152),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_2995),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_2924),
.B(n_351),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_2924),
.B(n_353),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_SL g3886 ( 
.A(n_3070),
.B(n_353),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_3070),
.B(n_354),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_L g3888 ( 
.A(n_3142),
.B(n_354),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_2997),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3004),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_3182),
.B(n_2996),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_2941),
.B(n_355),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3022),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3023),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_2941),
.B(n_355),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_2795),
.B(n_355),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_SL g3897 ( 
.A(n_3182),
.B(n_356),
.Y(n_3897)
);

OR2x2_ASAP7_75t_L g3898 ( 
.A(n_3228),
.B(n_356),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3036),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_2795),
.B(n_356),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_2798),
.B(n_357),
.Y(n_3901)
);

NOR2xp33_ASAP7_75t_L g3902 ( 
.A(n_3142),
.B(n_3153),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_2798),
.B(n_357),
.Y(n_3903)
);

INVxp67_ASAP7_75t_L g3904 ( 
.A(n_3211),
.Y(n_3904)
);

INVx3_ASAP7_75t_L g3905 ( 
.A(n_2901),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_2818),
.B(n_357),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_2803),
.Y(n_3907)
);

INVxp67_ASAP7_75t_L g3908 ( 
.A(n_3090),
.Y(n_3908)
);

OAI221xp5_ASAP7_75t_L g3909 ( 
.A1(n_3288),
.A2(n_360),
.B1(n_361),
.B2(n_359),
.C(n_358),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_2818),
.B(n_358),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_2938),
.A2(n_359),
.B1(n_361),
.B2(n_358),
.Y(n_3911)
);

AOI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3139),
.A2(n_362),
.B1(n_363),
.B2(n_359),
.Y(n_3912)
);

OAI22xp5_ASAP7_75t_L g3913 ( 
.A1(n_2843),
.A2(n_363),
.B1(n_364),
.B2(n_362),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_2991),
.B(n_362),
.Y(n_3914)
);

OAI21xp5_ASAP7_75t_L g3915 ( 
.A1(n_3378),
.A2(n_0),
.B(n_1),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_2843),
.B(n_363),
.Y(n_3916)
);

OR2x2_ASAP7_75t_L g3917 ( 
.A(n_3254),
.B(n_3263),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_SL g3918 ( 
.A(n_2996),
.B(n_364),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_3153),
.B(n_364),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3041),
.Y(n_3920)
);

AOI22xp5_ASAP7_75t_L g3921 ( 
.A1(n_3144),
.A2(n_366),
.B1(n_367),
.B2(n_365),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3043),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_2851),
.B(n_2858),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3044),
.Y(n_3924)
);

OAI22xp5_ASAP7_75t_L g3925 ( 
.A1(n_2851),
.A2(n_367),
.B1(n_368),
.B2(n_365),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_SL g3926 ( 
.A(n_3193),
.B(n_365),
.Y(n_3926)
);

AOI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3301),
.A2(n_368),
.B(n_367),
.Y(n_3927)
);

INVx3_ASAP7_75t_L g3928 ( 
.A(n_2901),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3049),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_SL g3930 ( 
.A(n_2824),
.B(n_368),
.Y(n_3930)
);

OAI22xp5_ASAP7_75t_L g3931 ( 
.A1(n_2858),
.A2(n_370),
.B1(n_371),
.B2(n_369),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_SL g3932 ( 
.A(n_2855),
.B(n_369),
.Y(n_3932)
);

BUFx3_ASAP7_75t_L g3933 ( 
.A(n_2817),
.Y(n_3933)
);

AOI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_2949),
.A2(n_371),
.B(n_370),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3052),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_SL g3936 ( 
.A(n_2855),
.B(n_370),
.Y(n_3936)
);

AOI22xp5_ASAP7_75t_L g3937 ( 
.A1(n_3146),
.A2(n_372),
.B1(n_373),
.B2(n_371),
.Y(n_3937)
);

BUFx3_ASAP7_75t_L g3938 ( 
.A(n_2828),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_L g3939 ( 
.A(n_2861),
.B(n_2862),
.Y(n_3939)
);

CKINVDCx5p33_ASAP7_75t_R g3940 ( 
.A(n_3152),
.Y(n_3940)
);

NOR2xp33_ASAP7_75t_L g3941 ( 
.A(n_3056),
.B(n_372),
.Y(n_3941)
);

NAND2xp33_ASAP7_75t_SL g3942 ( 
.A(n_2841),
.B(n_372),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_SL g3943 ( 
.A(n_2909),
.B(n_373),
.Y(n_3943)
);

OR2x2_ASAP7_75t_L g3944 ( 
.A(n_3287),
.B(n_373),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3299),
.A2(n_375),
.B1(n_376),
.B2(n_374),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3010),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_2861),
.B(n_2862),
.Y(n_3947)
);

NOR2xp33_ASAP7_75t_L g3948 ( 
.A(n_3056),
.B(n_2869),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_2942),
.B(n_374),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_2942),
.B(n_374),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_2955),
.B(n_375),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_2986),
.Y(n_3952)
);

INVx4_ASAP7_75t_L g3953 ( 
.A(n_3430),
.Y(n_3953)
);

INVxp67_ASAP7_75t_SL g3954 ( 
.A(n_3225),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_2958),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_2955),
.B(n_375),
.Y(n_3956)
);

OAI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3347),
.A2(n_377),
.B1(n_378),
.B2(n_376),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3087),
.A2(n_378),
.B(n_377),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_2881),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_SL g3960 ( 
.A(n_2909),
.B(n_378),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_2895),
.Y(n_3961)
);

OR2x2_ASAP7_75t_L g3962 ( 
.A(n_2994),
.B(n_379),
.Y(n_3962)
);

INVx4_ASAP7_75t_L g3963 ( 
.A(n_2983),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_SL g3964 ( 
.A(n_2918),
.B(n_3229),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3010),
.B(n_379),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3027),
.B(n_379),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_2937),
.Y(n_3967)
);

INVx3_ASAP7_75t_L g3968 ( 
.A(n_3347),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_2906),
.Y(n_3969)
);

NOR2xp33_ASAP7_75t_L g3970 ( 
.A(n_2884),
.B(n_380),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_2907),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_2937),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_2977),
.B(n_3000),
.Y(n_3973)
);

OAI22xp33_ASAP7_75t_L g3974 ( 
.A1(n_3154),
.A2(n_381),
.B1(n_382),
.B2(n_380),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3037),
.B(n_1),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_2907),
.Y(n_3976)
);

OAI22xp33_ASAP7_75t_L g3977 ( 
.A1(n_3154),
.A2(n_382),
.B1(n_383),
.B2(n_380),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_2803),
.Y(n_3978)
);

NOR2xp67_ASAP7_75t_L g3979 ( 
.A(n_2918),
.B(n_382),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_2977),
.B(n_383),
.Y(n_3980)
);

OAI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_2841),
.A2(n_384),
.B1(n_385),
.B2(n_383),
.Y(n_3981)
);

INVx2_ASAP7_75t_L g3982 ( 
.A(n_3094),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3000),
.B(n_384),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_SL g3984 ( 
.A(n_3229),
.B(n_385),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_2803),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3135),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3037),
.B(n_385),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3235),
.B(n_3436),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3054),
.B(n_3329),
.Y(n_3989)
);

INVxp67_ASAP7_75t_L g3990 ( 
.A(n_3090),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3251),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3053),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_SL g3993 ( 
.A(n_3237),
.B(n_386),
.Y(n_3993)
);

NAND3xp33_ASAP7_75t_L g3994 ( 
.A(n_2960),
.B(n_387),
.C(n_386),
.Y(n_3994)
);

AND2x4_ASAP7_75t_L g3995 ( 
.A(n_3051),
.B(n_386),
.Y(n_3995)
);

OR2x2_ASAP7_75t_SL g3996 ( 
.A(n_3127),
.B(n_387),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_SL g3997 ( 
.A(n_3237),
.B(n_387),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3053),
.Y(n_3998)
);

OAI22xp5_ASAP7_75t_L g3999 ( 
.A1(n_2863),
.A2(n_389),
.B1(n_390),
.B2(n_388),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3293),
.B(n_388),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3098),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3259),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_3293),
.B(n_388),
.Y(n_4003)
);

OR2x6_ASAP7_75t_L g4004 ( 
.A(n_2929),
.B(n_389),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_3309),
.B(n_3352),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3054),
.B(n_389),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3098),
.Y(n_4007)
);

INVx3_ASAP7_75t_L g4008 ( 
.A(n_2863),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_SL g4009 ( 
.A(n_3309),
.B(n_390),
.Y(n_4009)
);

NOR2xp33_ASAP7_75t_SL g4010 ( 
.A(n_3246),
.B(n_391),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3059),
.Y(n_4011)
);

OAI22xp33_ASAP7_75t_SL g4012 ( 
.A1(n_3090),
.A2(n_392),
.B1(n_394),
.B2(n_391),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3110),
.Y(n_4013)
);

NOR2xp33_ASAP7_75t_L g4014 ( 
.A(n_2885),
.B(n_391),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_SL g4015 ( 
.A(n_3352),
.B(n_392),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3110),
.Y(n_4016)
);

NAND2xp33_ASAP7_75t_L g4017 ( 
.A(n_3113),
.B(n_392),
.Y(n_4017)
);

BUFx4_ASAP7_75t_L g4018 ( 
.A(n_3180),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3011),
.B(n_393),
.Y(n_4019)
);

AO22x1_ASAP7_75t_L g4020 ( 
.A1(n_3452),
.A2(n_3120),
.B1(n_2797),
.B2(n_2822),
.Y(n_4020)
);

AOI22xp33_ASAP7_75t_SL g4021 ( 
.A1(n_3516),
.A2(n_3113),
.B1(n_2797),
.B2(n_2822),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3740),
.B(n_3136),
.Y(n_4022)
);

NOR3xp33_ASAP7_75t_L g4023 ( 
.A(n_3479),
.B(n_2886),
.C(n_3157),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3451),
.Y(n_4024)
);

NAND2x1p5_ASAP7_75t_L g4025 ( 
.A(n_3487),
.B(n_2983),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3649),
.B(n_3050),
.Y(n_4026)
);

NOR2x1p5_ASAP7_75t_L g4027 ( 
.A(n_3476),
.B(n_2830),
.Y(n_4027)
);

INVxp67_ASAP7_75t_L g4028 ( 
.A(n_3702),
.Y(n_4028)
);

OR2x6_ASAP7_75t_L g4029 ( 
.A(n_3755),
.B(n_2878),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_3544),
.B(n_3200),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3989),
.B(n_2833),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3457),
.Y(n_4032)
);

AOI22xp33_ASAP7_75t_L g4033 ( 
.A1(n_3536),
.A2(n_3161),
.B1(n_2929),
.B2(n_3099),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3645),
.B(n_3165),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3556),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3557),
.Y(n_4036)
);

AND2x4_ASAP7_75t_L g4037 ( 
.A(n_3757),
.B(n_2875),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3471),
.Y(n_4038)
);

OR2x2_ASAP7_75t_L g4039 ( 
.A(n_3917),
.B(n_2944),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3902),
.B(n_3129),
.Y(n_4040)
);

INVx2_ASAP7_75t_SL g4041 ( 
.A(n_3571),
.Y(n_4041)
);

NOR2xp33_ASAP7_75t_L g4042 ( 
.A(n_3786),
.B(n_3196),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_SL g4043 ( 
.A(n_3452),
.B(n_2875),
.Y(n_4043)
);

AND2x4_ASAP7_75t_L g4044 ( 
.A(n_3757),
.B(n_3968),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3481),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3568),
.Y(n_4046)
);

NOR2xp33_ASAP7_75t_L g4047 ( 
.A(n_3606),
.B(n_3512),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3566),
.B(n_3097),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_SL g4049 ( 
.A(n_3642),
.B(n_3361),
.Y(n_4049)
);

NOR2xp67_ASAP7_75t_L g4050 ( 
.A(n_3968),
.B(n_2914),
.Y(n_4050)
);

NOR2xp33_ASAP7_75t_L g4051 ( 
.A(n_3512),
.B(n_3202),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3973),
.B(n_3111),
.Y(n_4052)
);

OR2x6_ASAP7_75t_L g4053 ( 
.A(n_3755),
.B(n_3001),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3520),
.B(n_3115),
.Y(n_4054)
);

O2A1O1Ixp5_ASAP7_75t_L g4055 ( 
.A1(n_3891),
.A2(n_2910),
.B(n_3339),
.C(n_3337),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3642),
.B(n_3361),
.Y(n_4056)
);

O2A1O1Ixp33_ASAP7_75t_L g4057 ( 
.A1(n_3689),
.A2(n_3155),
.B(n_3088),
.C(n_3099),
.Y(n_4057)
);

INVxp67_ASAP7_75t_L g4058 ( 
.A(n_3853),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3491),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3494),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3532),
.B(n_3116),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3535),
.B(n_3118),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_L g4063 ( 
.A(n_3550),
.B(n_3123),
.Y(n_4063)
);

AND2x6_ASAP7_75t_SL g4064 ( 
.A(n_3696),
.B(n_3198),
.Y(n_4064)
);

AOI22xp5_ASAP7_75t_L g4065 ( 
.A1(n_3757),
.A2(n_2990),
.B1(n_3100),
.B2(n_3040),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3504),
.Y(n_4066)
);

AND2x6_ASAP7_75t_SL g4067 ( 
.A(n_4004),
.B(n_3201),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3510),
.Y(n_4068)
);

AOI22xp5_ASAP7_75t_L g4069 ( 
.A1(n_4004),
.A2(n_3316),
.B1(n_3160),
.B2(n_3197),
.Y(n_4069)
);

INVx3_ASAP7_75t_L g4070 ( 
.A(n_3571),
.Y(n_4070)
);

INVxp67_ASAP7_75t_L g4071 ( 
.A(n_3988),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3589),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3562),
.B(n_3124),
.Y(n_4073)
);

INVx2_ASAP7_75t_SL g4074 ( 
.A(n_3571),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_SL g4075 ( 
.A1(n_3996),
.A2(n_4004),
.B1(n_3783),
.B2(n_3879),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3514),
.Y(n_4076)
);

AOI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_3513),
.A2(n_3161),
.B1(n_2929),
.B2(n_3088),
.Y(n_4077)
);

AND2x4_ASAP7_75t_L g4078 ( 
.A(n_3580),
.B(n_2914),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_3567),
.B(n_3050),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3531),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3447),
.Y(n_4081)
);

INVx3_ASAP7_75t_L g4082 ( 
.A(n_3485),
.Y(n_4082)
);

OAI22xp33_ASAP7_75t_L g4083 ( 
.A1(n_3783),
.A2(n_3197),
.B1(n_3204),
.B2(n_3366),
.Y(n_4083)
);

INVx2_ASAP7_75t_L g4084 ( 
.A(n_3594),
.Y(n_4084)
);

BUFx3_ASAP7_75t_L g4085 ( 
.A(n_3487),
.Y(n_4085)
);

AOI22xp33_ASAP7_75t_L g4086 ( 
.A1(n_3704),
.A2(n_3358),
.B1(n_3393),
.B2(n_3343),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3455),
.Y(n_4087)
);

BUFx3_ASAP7_75t_L g4088 ( 
.A(n_3487),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3461),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3627),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3629),
.Y(n_4091)
);

AND2x6_ASAP7_75t_SL g4092 ( 
.A(n_3783),
.B(n_3330),
.Y(n_4092)
);

NOR2xp33_ASAP7_75t_SL g4093 ( 
.A(n_3573),
.B(n_3366),
.Y(n_4093)
);

INVxp67_ASAP7_75t_L g4094 ( 
.A(n_3954),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3668),
.B(n_3081),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3537),
.B(n_3081),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3493),
.B(n_3122),
.Y(n_4097)
);

AOI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3540),
.A2(n_3405),
.B1(n_3443),
.B2(n_3428),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3502),
.B(n_3128),
.Y(n_4099)
);

BUFx6f_ASAP7_75t_L g4100 ( 
.A(n_3533),
.Y(n_4100)
);

BUFx6f_ASAP7_75t_L g4101 ( 
.A(n_3533),
.Y(n_4101)
);

INVx2_ASAP7_75t_SL g4102 ( 
.A(n_3546),
.Y(n_4102)
);

AOI22xp33_ASAP7_75t_L g4103 ( 
.A1(n_3671),
.A2(n_3445),
.B1(n_3199),
.B2(n_3071),
.Y(n_4103)
);

AOI22xp5_ASAP7_75t_L g4104 ( 
.A1(n_3540),
.A2(n_3195),
.B1(n_3199),
.B2(n_3163),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_L g4105 ( 
.A(n_3565),
.B(n_3128),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_3741),
.B(n_2900),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3643),
.Y(n_4107)
);

NOR2x2_ASAP7_75t_L g4108 ( 
.A(n_3879),
.B(n_3203),
.Y(n_4108)
);

NAND2x1p5_ASAP7_75t_L g4109 ( 
.A(n_3963),
.B(n_3001),
.Y(n_4109)
);

NOR2xp67_ASAP7_75t_L g4110 ( 
.A(n_3636),
.B(n_3640),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_3923),
.B(n_2852),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3939),
.B(n_3177),
.Y(n_4112)
);

BUFx6f_ASAP7_75t_L g4113 ( 
.A(n_3533),
.Y(n_4113)
);

NOR2xp33_ASAP7_75t_L g4114 ( 
.A(n_3559),
.B(n_3188),
.Y(n_4114)
);

NOR2xp33_ASAP7_75t_L g4115 ( 
.A(n_3908),
.B(n_3190),
.Y(n_4115)
);

INVx1_ASAP7_75t_SL g4116 ( 
.A(n_3933),
.Y(n_4116)
);

INVx3_ASAP7_75t_L g4117 ( 
.A(n_3963),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3467),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_3947),
.B(n_3186),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3501),
.B(n_3163),
.Y(n_4120)
);

BUFx6f_ASAP7_75t_L g4121 ( 
.A(n_3585),
.Y(n_4121)
);

O2A1O1Ixp5_ASAP7_75t_L g4122 ( 
.A1(n_3483),
.A2(n_3015),
.B(n_3272),
.C(n_2805),
.Y(n_4122)
);

OR2x2_ASAP7_75t_L g4123 ( 
.A(n_3790),
.B(n_2786),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_3506),
.B(n_2839),
.Y(n_4124)
);

AOI22xp33_ASAP7_75t_L g4125 ( 
.A1(n_3795),
.A2(n_3315),
.B1(n_3324),
.B2(n_3323),
.Y(n_4125)
);

NAND2xp33_ASAP7_75t_L g4126 ( 
.A(n_3834),
.B(n_2797),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_L g4127 ( 
.A(n_3448),
.B(n_3191),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_SL g4128 ( 
.A(n_3701),
.B(n_3370),
.Y(n_4128)
);

AOI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_3669),
.A2(n_3179),
.B1(n_3132),
.B2(n_3076),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_SL g4130 ( 
.A(n_3701),
.B(n_3370),
.Y(n_4130)
);

O2A1O1Ixp33_ASAP7_75t_L g4131 ( 
.A1(n_3677),
.A2(n_3132),
.B(n_3332),
.C(n_3282),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_SL g4132 ( 
.A(n_4010),
.B(n_3456),
.Y(n_4132)
);

AND2x4_ASAP7_75t_L g4133 ( 
.A(n_3580),
.B(n_2936),
.Y(n_4133)
);

CKINVDCx11_ASAP7_75t_R g4134 ( 
.A(n_3882),
.Y(n_4134)
);

NOR2xp33_ASAP7_75t_L g4135 ( 
.A(n_3990),
.B(n_3192),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3478),
.B(n_3881),
.Y(n_4136)
);

NOR2xp33_ASAP7_75t_L g4137 ( 
.A(n_3524),
.B(n_3171),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3542),
.B(n_3063),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3547),
.B(n_3063),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3644),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_L g4141 ( 
.A1(n_3800),
.A2(n_2822),
.B1(n_2815),
.B2(n_2797),
.Y(n_4141)
);

NOR2xp33_ASAP7_75t_L g4142 ( 
.A(n_3609),
.B(n_3876),
.Y(n_4142)
);

BUFx6f_ASAP7_75t_L g4143 ( 
.A(n_3585),
.Y(n_4143)
);

AOI22xp33_ASAP7_75t_L g4144 ( 
.A1(n_3592),
.A2(n_2815),
.B1(n_2838),
.B2(n_2822),
.Y(n_4144)
);

OR2x2_ASAP7_75t_L g4145 ( 
.A(n_3673),
.B(n_2800),
.Y(n_4145)
);

AOI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_3807),
.A2(n_3127),
.B1(n_3101),
.B2(n_2988),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_3548),
.B(n_3275),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3474),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3551),
.B(n_3295),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_3655),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_4010),
.B(n_3427),
.Y(n_4151)
);

NAND2x1p5_ASAP7_75t_L g4152 ( 
.A(n_3953),
.B(n_3026),
.Y(n_4152)
);

INVxp67_ASAP7_75t_L g4153 ( 
.A(n_3806),
.Y(n_4153)
);

INVx3_ASAP7_75t_L g4154 ( 
.A(n_3755),
.Y(n_4154)
);

AND2x6_ASAP7_75t_SL g4155 ( 
.A(n_3879),
.B(n_3227),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3475),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3477),
.Y(n_4157)
);

BUFx6f_ASAP7_75t_L g4158 ( 
.A(n_3585),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_3664),
.Y(n_4159)
);

NOR2xp33_ASAP7_75t_L g4160 ( 
.A(n_3904),
.B(n_3189),
.Y(n_4160)
);

NOR2x2_ASAP7_75t_L g4161 ( 
.A(n_3573),
.B(n_3194),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_3678),
.Y(n_4162)
);

AOI22xp5_ASAP7_75t_L g4163 ( 
.A1(n_3657),
.A2(n_3217),
.B1(n_3159),
.B2(n_3073),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3489),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3554),
.B(n_3133),
.Y(n_4165)
);

OAI22xp5_ASAP7_75t_SL g4166 ( 
.A1(n_3666),
.A2(n_3442),
.B1(n_3427),
.B2(n_3264),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_3560),
.B(n_3133),
.Y(n_4167)
);

OR2x2_ASAP7_75t_L g4168 ( 
.A(n_3898),
.B(n_3216),
.Y(n_4168)
);

CKINVDCx5p33_ASAP7_75t_R g4169 ( 
.A(n_3579),
.Y(n_4169)
);

BUFx3_ASAP7_75t_L g4170 ( 
.A(n_3938),
.Y(n_4170)
);

CKINVDCx20_ASAP7_75t_R g4171 ( 
.A(n_3633),
.Y(n_4171)
);

AOI22xp33_ASAP7_75t_SL g4172 ( 
.A1(n_3507),
.A2(n_2838),
.B1(n_2815),
.B2(n_3204),
.Y(n_4172)
);

NOR2xp33_ASAP7_75t_L g4173 ( 
.A(n_3813),
.B(n_3291),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3505),
.Y(n_4174)
);

INVx3_ASAP7_75t_L g4175 ( 
.A(n_3707),
.Y(n_4175)
);

NOR2xp33_ASAP7_75t_L g4176 ( 
.A(n_3646),
.B(n_3310),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_3684),
.Y(n_4177)
);

NOR2xp33_ASAP7_75t_L g4178 ( 
.A(n_3760),
.B(n_3334),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3515),
.Y(n_4179)
);

NOR2xp33_ASAP7_75t_L g4180 ( 
.A(n_3496),
.B(n_3367),
.Y(n_4180)
);

OAI22xp5_ASAP7_75t_SL g4181 ( 
.A1(n_3776),
.A2(n_3442),
.B1(n_3408),
.B2(n_3033),
.Y(n_4181)
);

AOI22xp33_ASAP7_75t_SL g4182 ( 
.A1(n_3507),
.A2(n_2838),
.B1(n_2815),
.B2(n_2992),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3522),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_3692),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3561),
.B(n_2950),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_3703),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3527),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3563),
.B(n_3003),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_3708),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3463),
.Y(n_4190)
);

NOR2xp33_ASAP7_75t_L g4191 ( 
.A(n_3948),
.B(n_2844),
.Y(n_4191)
);

NOR2x2_ASAP7_75t_L g4192 ( 
.A(n_3729),
.B(n_3227),
.Y(n_4192)
);

NAND2xp5_ASAP7_75t_L g4193 ( 
.A(n_3497),
.B(n_3459),
.Y(n_4193)
);

NAND2x1p5_ASAP7_75t_L g4194 ( 
.A(n_3953),
.B(n_3026),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3797),
.B(n_3570),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_3584),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_3587),
.Y(n_4197)
);

CKINVDCx5p33_ASAP7_75t_R g4198 ( 
.A(n_3612),
.Y(n_4198)
);

INVx2_ASAP7_75t_L g4199 ( 
.A(n_3715),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_SL g4200 ( 
.A1(n_3619),
.A2(n_3058),
.B1(n_3130),
.B2(n_3033),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_3600),
.B(n_3173),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3602),
.B(n_3607),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_3716),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3610),
.B(n_3173),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_3617),
.B(n_3178),
.Y(n_4205)
);

BUFx4f_ASAP7_75t_L g4206 ( 
.A(n_3753),
.Y(n_4206)
);

HB1xp67_ASAP7_75t_L g4207 ( 
.A(n_3525),
.Y(n_4207)
);

AND2x4_ASAP7_75t_L g4208 ( 
.A(n_3707),
.B(n_2936),
.Y(n_4208)
);

NAND2x1_ASAP7_75t_L g4209 ( 
.A(n_3626),
.B(n_3441),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_SL g4210 ( 
.A(n_3456),
.B(n_3058),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_3734),
.Y(n_4211)
);

AOI221xp5_ASAP7_75t_L g4212 ( 
.A1(n_3637),
.A2(n_3178),
.B1(n_3156),
.B2(n_2954),
.C(n_3002),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_3618),
.B(n_2877),
.Y(n_4213)
);

A2O1A1Ixp33_ASAP7_75t_L g4214 ( 
.A1(n_3727),
.A2(n_3117),
.B(n_2965),
.C(n_2975),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3622),
.Y(n_4215)
);

AOI22xp33_ASAP7_75t_L g4216 ( 
.A1(n_3596),
.A2(n_2838),
.B1(n_3117),
.B2(n_3104),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_SL g4217 ( 
.A(n_3834),
.B(n_3130),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_3624),
.B(n_2916),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_3628),
.B(n_3205),
.Y(n_4219)
);

AND2x2_ASAP7_75t_L g4220 ( 
.A(n_3500),
.B(n_2867),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3747),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_SL g4222 ( 
.A(n_3834),
.B(n_2846),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_SL g4223 ( 
.A(n_3834),
.B(n_2864),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_3638),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_3660),
.B(n_3224),
.Y(n_4225)
);

NOR2xp33_ASAP7_75t_L g4226 ( 
.A(n_3852),
.B(n_3167),
.Y(n_4226)
);

NAND2xp33_ASAP7_75t_L g4227 ( 
.A(n_3834),
.B(n_3441),
.Y(n_4227)
);

OR2x2_ASAP7_75t_L g4228 ( 
.A(n_3944),
.B(n_3187),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_3663),
.B(n_3241),
.Y(n_4229)
);

INVx1_ASAP7_75t_SL g4230 ( 
.A(n_4018),
.Y(n_4230)
);

AOI22xp5_ASAP7_75t_L g4231 ( 
.A1(n_3812),
.A2(n_2989),
.B1(n_3012),
.B2(n_2972),
.Y(n_4231)
);

BUFx6f_ASAP7_75t_L g4232 ( 
.A(n_3616),
.Y(n_4232)
);

NOR2xp33_ASAP7_75t_L g4233 ( 
.A(n_3962),
.B(n_2943),
.Y(n_4233)
);

AOI22xp33_ASAP7_75t_SL g4234 ( 
.A1(n_3588),
.A2(n_2992),
.B1(n_3083),
.B2(n_3441),
.Y(n_4234)
);

AOI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_3822),
.A2(n_3060),
.B1(n_3080),
.B2(n_3065),
.Y(n_4235)
);

HB1xp67_ASAP7_75t_L g4236 ( 
.A(n_3690),
.Y(n_4236)
);

INVxp67_ASAP7_75t_L g4237 ( 
.A(n_3746),
.Y(n_4237)
);

NAND3xp33_ASAP7_75t_SL g4238 ( 
.A(n_3651),
.B(n_3121),
.C(n_3109),
.Y(n_4238)
);

NOR2xp33_ASAP7_75t_L g4239 ( 
.A(n_3661),
.B(n_2951),
.Y(n_4239)
);

NOR2xp33_ASAP7_75t_SL g4240 ( 
.A(n_3729),
.B(n_2896),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_SL g4241 ( 
.A(n_3816),
.B(n_2920),
.Y(n_4241)
);

A2O1A1Ixp33_ASAP7_75t_L g4242 ( 
.A1(n_3735),
.A2(n_2965),
.B(n_2975),
.C(n_2984),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_3665),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_3816),
.B(n_2927),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_L g4245 ( 
.A(n_3722),
.B(n_3016),
.Y(n_4245)
);

NOR2xp33_ASAP7_75t_SL g4246 ( 
.A(n_3940),
.B(n_3107),
.Y(n_4246)
);

CKINVDCx5p33_ASAP7_75t_R g4247 ( 
.A(n_3865),
.Y(n_4247)
);

BUFx3_ASAP7_75t_L g4248 ( 
.A(n_3731),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_3687),
.B(n_3270),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_3709),
.B(n_3285),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_3569),
.B(n_3312),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_3572),
.B(n_3317),
.Y(n_4252)
);

AOI22xp33_ASAP7_75t_L g4253 ( 
.A1(n_3521),
.A2(n_3082),
.B1(n_3140),
.B2(n_3083),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_3530),
.B(n_3331),
.Y(n_4254)
);

CKINVDCx5p33_ASAP7_75t_R g4255 ( 
.A(n_3647),
.Y(n_4255)
);

INVx2_ASAP7_75t_SL g4256 ( 
.A(n_3731),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_3526),
.B(n_3344),
.Y(n_4257)
);

INVx2_ASAP7_75t_SL g4258 ( 
.A(n_3453),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_SL g4259 ( 
.A(n_3915),
.B(n_2868),
.Y(n_4259)
);

NOR2xp67_ASAP7_75t_L g4260 ( 
.A(n_3636),
.B(n_3248),
.Y(n_4260)
);

AOI22xp5_ASAP7_75t_L g4261 ( 
.A1(n_3764),
.A2(n_3737),
.B1(n_3791),
.B2(n_4017),
.Y(n_4261)
);

INVx2_ASAP7_75t_L g4262 ( 
.A(n_3756),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_3714),
.B(n_3380),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_3733),
.B(n_3388),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_SL g4265 ( 
.A(n_3915),
.B(n_3248),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_3738),
.Y(n_4266)
);

AOI22xp5_ASAP7_75t_L g4267 ( 
.A1(n_3630),
.A2(n_3091),
.B1(n_3175),
.B2(n_2998),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_3748),
.Y(n_4268)
);

NOR3x1_ASAP7_75t_L g4269 ( 
.A(n_3994),
.B(n_3121),
.C(n_3395),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_3752),
.Y(n_4270)
);

NOR2xp33_ASAP7_75t_L g4271 ( 
.A(n_3918),
.B(n_2904),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_3759),
.B(n_3137),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_3768),
.Y(n_4273)
);

BUFx3_ASAP7_75t_L g4274 ( 
.A(n_3695),
.Y(n_4274)
);

OR2x2_ASAP7_75t_L g4275 ( 
.A(n_3541),
.B(n_3141),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3761),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_SL g4277 ( 
.A(n_3458),
.B(n_3248),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3766),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3975),
.B(n_3143),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_3975),
.B(n_3156),
.Y(n_4280)
);

OR2x2_ASAP7_75t_L g4281 ( 
.A(n_3543),
.B(n_3150),
.Y(n_4281)
);

OR2x2_ASAP7_75t_L g4282 ( 
.A(n_3553),
.B(n_3168),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_L g4283 ( 
.A(n_3859),
.B(n_2834),
.Y(n_4283)
);

INVx2_ASAP7_75t_SL g4284 ( 
.A(n_3495),
.Y(n_4284)
);

INVx3_ASAP7_75t_L g4285 ( 
.A(n_3626),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_3648),
.B(n_2834),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_3773),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_3771),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_3772),
.Y(n_4289)
);

INVx6_ASAP7_75t_L g4290 ( 
.A(n_3869),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_3769),
.B(n_3206),
.Y(n_4291)
);

BUFx3_ASAP7_75t_L g4292 ( 
.A(n_3706),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_3777),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_SL g4294 ( 
.A(n_3732),
.B(n_3277),
.Y(n_4294)
);

NOR2xp33_ASAP7_75t_L g4295 ( 
.A(n_3691),
.B(n_3145),
.Y(n_4295)
);

AOI22xp5_ASAP7_75t_L g4296 ( 
.A1(n_3652),
.A2(n_3055),
.B1(n_3095),
.B2(n_3072),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_3770),
.B(n_3206),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_SL g4298 ( 
.A(n_3732),
.B(n_3277),
.Y(n_4298)
);

NAND2x1p5_ASAP7_75t_L g4299 ( 
.A(n_3670),
.B(n_3675),
.Y(n_4299)
);

OAI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_3994),
.A2(n_3801),
.B1(n_3802),
.B2(n_3880),
.Y(n_4300)
);

AND2x2_ASAP7_75t_L g4301 ( 
.A(n_3604),
.B(n_3267),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_3774),
.B(n_3267),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_3794),
.Y(n_4303)
);

AOI22xp33_ASAP7_75t_L g4304 ( 
.A1(n_3785),
.A2(n_2992),
.B1(n_3083),
.B2(n_3342),
.Y(n_4304)
);

NOR2xp33_ASAP7_75t_L g4305 ( 
.A(n_3480),
.B(n_3148),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_SL g4306 ( 
.A(n_3711),
.B(n_3277),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_3803),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_3811),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_3623),
.B(n_3342),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_L g4310 ( 
.A(n_3863),
.B(n_3112),
.Y(n_4310)
);

AOI22xp33_ASAP7_75t_L g4311 ( 
.A1(n_3574),
.A2(n_2992),
.B1(n_3083),
.B2(n_3381),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_3914),
.B(n_3381),
.Y(n_4312)
);

AND2x6_ASAP7_75t_SL g4313 ( 
.A(n_3472),
.B(n_3373),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_3780),
.B(n_3419),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3814),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_3599),
.B(n_3419),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_3775),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_3782),
.B(n_3158),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_3827),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_3784),
.B(n_3158),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3835),
.Y(n_4321)
);

INVx4_ASAP7_75t_L g4322 ( 
.A(n_3625),
.Y(n_4322)
);

OR2x2_ASAP7_75t_L g4323 ( 
.A(n_3788),
.B(n_3034),
.Y(n_4323)
);

BUFx6f_ASAP7_75t_SL g4324 ( 
.A(n_3995),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_3789),
.B(n_3162),
.Y(n_4325)
);

AOI22xp33_ASAP7_75t_L g4326 ( 
.A1(n_3590),
.A2(n_3068),
.B1(n_2984),
.B2(n_3162),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_3888),
.B(n_3048),
.Y(n_4327)
);

AND2x2_ASAP7_75t_L g4328 ( 
.A(n_3995),
.B(n_3048),
.Y(n_4328)
);

AND2x2_ASAP7_75t_L g4329 ( 
.A(n_3796),
.B(n_393),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_3828),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_SL g4331 ( 
.A(n_3640),
.B(n_3300),
.Y(n_4331)
);

INVx4_ASAP7_75t_L g4332 ( 
.A(n_3625),
.Y(n_4332)
);

AND2x4_ASAP7_75t_L g4333 ( 
.A(n_3840),
.B(n_3068),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_3839),
.Y(n_4334)
);

INVx2_ASAP7_75t_SL g4335 ( 
.A(n_3718),
.Y(n_4335)
);

NAND2x1p5_ASAP7_75t_L g4336 ( 
.A(n_3720),
.B(n_3373),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_3866),
.Y(n_4337)
);

NOR2xp67_ASAP7_75t_L g4338 ( 
.A(n_3710),
.B(n_3300),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_3847),
.Y(n_4339)
);

INVx3_ASAP7_75t_L g4340 ( 
.A(n_3781),
.Y(n_4340)
);

AOI22xp33_ASAP7_75t_L g4341 ( 
.A1(n_3919),
.A2(n_3108),
.B1(n_3308),
.B2(n_3300),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_3941),
.B(n_393),
.Y(n_4342)
);

OR2x2_ASAP7_75t_L g4343 ( 
.A(n_3848),
.B(n_394),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_3986),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_SL g4345 ( 
.A(n_3710),
.B(n_3308),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_3519),
.B(n_394),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_3877),
.Y(n_4347)
);

CKINVDCx5p33_ASAP7_75t_R g4348 ( 
.A(n_3964),
.Y(n_4348)
);

A2O1A1Ixp33_ASAP7_75t_L g4349 ( 
.A1(n_3942),
.A2(n_3333),
.B(n_3391),
.C(n_3308),
.Y(n_4349)
);

AOI21xp5_ASAP7_75t_L g4350 ( 
.A1(n_3473),
.A2(n_3391),
.B(n_3333),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_3713),
.B(n_395),
.Y(n_4351)
);

NOR2xp33_ASAP7_75t_L g4352 ( 
.A(n_3809),
.B(n_3439),
.Y(n_4352)
);

AOI22xp33_ASAP7_75t_SL g4353 ( 
.A1(n_4012),
.A2(n_3391),
.B1(n_3415),
.B2(n_3333),
.Y(n_4353)
);

OAI21xp5_ASAP7_75t_L g4354 ( 
.A1(n_3832),
.A2(n_3028),
.B(n_3008),
.Y(n_4354)
);

AOI22xp33_ASAP7_75t_L g4355 ( 
.A1(n_3763),
.A2(n_3424),
.B1(n_3435),
.B2(n_3415),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_SL g4356 ( 
.A(n_3799),
.B(n_3415),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_3883),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_3889),
.Y(n_4358)
);

NOR2xp33_ASAP7_75t_L g4359 ( 
.A(n_3717),
.B(n_3439),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_3890),
.Y(n_4360)
);

AOI22xp33_ASAP7_75t_SL g4361 ( 
.A1(n_4012),
.A2(n_3435),
.B1(n_3424),
.B2(n_3028),
.Y(n_4361)
);

AOI22xp33_ASAP7_75t_L g4362 ( 
.A1(n_3730),
.A2(n_3435),
.B1(n_3424),
.B2(n_3028),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_3894),
.Y(n_4363)
);

BUFx6f_ASAP7_75t_L g4364 ( 
.A(n_3616),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_3721),
.B(n_3724),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_3621),
.B(n_1069),
.Y(n_4366)
);

CKINVDCx5p33_ASAP7_75t_R g4367 ( 
.A(n_4005),
.Y(n_4367)
);

INVx2_ASAP7_75t_L g4368 ( 
.A(n_3855),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_3864),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_3899),
.Y(n_4370)
);

INVx3_ASAP7_75t_L g4371 ( 
.A(n_3781),
.Y(n_4371)
);

AOI22xp33_ASAP7_75t_L g4372 ( 
.A1(n_3909),
.A2(n_3046),
.B1(n_3069),
.B2(n_3008),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_SL g4373 ( 
.A(n_3979),
.B(n_3482),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_3725),
.B(n_395),
.Y(n_4374)
);

INVx3_ASAP7_75t_L g4375 ( 
.A(n_3597),
.Y(n_4375)
);

INVx2_ASAP7_75t_SL g4376 ( 
.A(n_3503),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_3728),
.B(n_396),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_3920),
.Y(n_4378)
);

BUFx4f_ASAP7_75t_L g4379 ( 
.A(n_3508),
.Y(n_4379)
);

AOI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_3880),
.A2(n_3046),
.B1(n_3069),
.B2(n_3008),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_3736),
.B(n_3742),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_3743),
.B(n_396),
.Y(n_4382)
);

BUFx3_ASAP7_75t_L g4383 ( 
.A(n_3564),
.Y(n_4383)
);

OAI22xp5_ASAP7_75t_L g4384 ( 
.A1(n_3815),
.A2(n_3069),
.B1(n_3079),
.B2(n_3046),
.Y(n_4384)
);

AOI22xp5_ASAP7_75t_L g4385 ( 
.A1(n_3862),
.A2(n_3079),
.B1(n_397),
.B2(n_398),
.Y(n_4385)
);

AND2x4_ASAP7_75t_L g4386 ( 
.A(n_3978),
.B(n_3079),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_3929),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_SL g4388 ( 
.A(n_3545),
.B(n_396),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_3792),
.B(n_1071),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_3872),
.Y(n_4390)
);

NOR2xp33_ASAP7_75t_SL g4391 ( 
.A(n_3957),
.B(n_3632),
.Y(n_4391)
);

BUFx3_ASAP7_75t_L g4392 ( 
.A(n_3586),
.Y(n_4392)
);

INVxp33_ASAP7_75t_L g4393 ( 
.A(n_3465),
.Y(n_4393)
);

OAI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_3854),
.A2(n_3913),
.B1(n_3931),
.B2(n_3925),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_3767),
.B(n_397),
.Y(n_4395)
);

NOR2xp33_ASAP7_75t_L g4396 ( 
.A(n_3823),
.B(n_398),
.Y(n_4396)
);

INVx4_ASAP7_75t_L g4397 ( 
.A(n_3601),
.Y(n_4397)
);

INVx4_ASAP7_75t_L g4398 ( 
.A(n_3679),
.Y(n_4398)
);

INVx8_ASAP7_75t_L g4399 ( 
.A(n_3549),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_3620),
.B(n_398),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_3935),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_SL g4402 ( 
.A(n_3611),
.B(n_399),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_3634),
.B(n_3639),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_3641),
.B(n_399),
.Y(n_4404)
);

BUFx2_ASAP7_75t_L g4405 ( 
.A(n_3907),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_3871),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_SL g4407 ( 
.A(n_3549),
.B(n_400),
.Y(n_4407)
);

AOI22xp33_ASAP7_75t_L g4408 ( 
.A1(n_3820),
.A2(n_401),
.B1(n_402),
.B2(n_400),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_3650),
.B(n_400),
.Y(n_4409)
);

AOI22xp5_ASAP7_75t_L g4410 ( 
.A1(n_3970),
.A2(n_403),
.B1(n_404),
.B2(n_401),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_3893),
.Y(n_4411)
);

AOI22xp5_ASAP7_75t_L g4412 ( 
.A1(n_4014),
.A2(n_405),
.B1(n_406),
.B2(n_403),
.Y(n_4412)
);

AOI22xp33_ASAP7_75t_L g4413 ( 
.A1(n_3744),
.A2(n_405),
.B1(n_406),
.B2(n_403),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_3653),
.B(n_407),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_3654),
.B(n_409),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_3656),
.B(n_409),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_3874),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_L g4418 ( 
.A(n_3658),
.B(n_409),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_SL g4419 ( 
.A(n_3957),
.B(n_410),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_L g4420 ( 
.A(n_3659),
.B(n_411),
.Y(n_4420)
);

OAI22xp5_ASAP7_75t_L g4421 ( 
.A1(n_3913),
.A2(n_412),
.B1(n_413),
.B2(n_411),
.Y(n_4421)
);

AND2x2_ASAP7_75t_L g4422 ( 
.A(n_3468),
.B(n_1068),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_3924),
.Y(n_4423)
);

AND2x4_ASAP7_75t_SL g4424 ( 
.A(n_3992),
.B(n_3998),
.Y(n_4424)
);

AOI22xp5_ASAP7_75t_L g4425 ( 
.A1(n_3829),
.A2(n_412),
.B1(n_413),
.B2(n_411),
.Y(n_4425)
);

AOI22xp33_ASAP7_75t_L g4426 ( 
.A1(n_3750),
.A2(n_414),
.B1(n_415),
.B2(n_412),
.Y(n_4426)
);

NAND2xp5_ASAP7_75t_L g4427 ( 
.A(n_3672),
.B(n_414),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_SL g4428 ( 
.A(n_3739),
.B(n_414),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_SL g4429 ( 
.A(n_3739),
.B(n_415),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_SL g4430 ( 
.A(n_3925),
.B(n_416),
.Y(n_4430)
);

CKINVDCx20_ASAP7_75t_R g4431 ( 
.A(n_3529),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_3674),
.B(n_416),
.Y(n_4432)
);

AOI22xp33_ASAP7_75t_L g4433 ( 
.A1(n_3837),
.A2(n_4019),
.B1(n_3608),
.B2(n_3931),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_3697),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_3698),
.Y(n_4435)
);

AOI22xp33_ASAP7_75t_L g4436 ( 
.A1(n_3446),
.A2(n_417),
.B1(n_418),
.B2(n_416),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_3922),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_3700),
.Y(n_4438)
);

AOI22xp5_ASAP7_75t_L g4439 ( 
.A1(n_3974),
.A2(n_3977),
.B1(n_3911),
.B2(n_3779),
.Y(n_4439)
);

BUFx6f_ASAP7_75t_SL g4440 ( 
.A(n_3991),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_3712),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_3676),
.B(n_417),
.Y(n_4442)
);

AOI22xp5_ASAP7_75t_L g4443 ( 
.A1(n_3817),
.A2(n_419),
.B1(n_420),
.B2(n_418),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_3680),
.B(n_419),
.Y(n_4444)
);

OR2x6_ASAP7_75t_L g4445 ( 
.A(n_3449),
.B(n_420),
.Y(n_4445)
);

AOI22xp33_ASAP7_75t_SL g4446 ( 
.A1(n_3667),
.A2(n_421),
.B1(n_422),
.B2(n_420),
.Y(n_4446)
);

INVx4_ASAP7_75t_L g4447 ( 
.A(n_3616),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_3955),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_3683),
.B(n_421),
.Y(n_4449)
);

AOI22xp5_ASAP7_75t_L g4450 ( 
.A1(n_3778),
.A2(n_422),
.B1(n_423),
.B2(n_421),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_3685),
.B(n_422),
.Y(n_4451)
);

AOI22xp33_ASAP7_75t_L g4452 ( 
.A1(n_3591),
.A2(n_424),
.B1(n_425),
.B2(n_423),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_3686),
.B(n_423),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_3693),
.B(n_426),
.Y(n_4454)
);

AOI22xp5_ASAP7_75t_L g4455 ( 
.A1(n_3787),
.A2(n_427),
.B1(n_428),
.B2(n_426),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_SL g4456 ( 
.A(n_3534),
.B(n_427),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4011),
.Y(n_4457)
);

NOR2xp33_ASAP7_75t_L g4458 ( 
.A(n_3826),
.B(n_427),
.Y(n_4458)
);

NOR2xp33_ASAP7_75t_L g4459 ( 
.A(n_3946),
.B(n_428),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_3470),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_3470),
.Y(n_4461)
);

INVx2_ASAP7_75t_L g4462 ( 
.A(n_3982),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_SL g4463 ( 
.A(n_3981),
.B(n_429),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_3450),
.Y(n_4464)
);

AOI22xp33_ASAP7_75t_L g4465 ( 
.A1(n_3603),
.A2(n_430),
.B1(n_431),
.B2(n_429),
.Y(n_4465)
);

AOI22xp33_ASAP7_75t_L g4466 ( 
.A1(n_3662),
.A2(n_3987),
.B1(n_3682),
.B2(n_4006),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_SL g4467 ( 
.A(n_3981),
.B(n_430),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_3694),
.B(n_430),
.Y(n_4468)
);

INVx2_ASAP7_75t_L g4469 ( 
.A(n_3959),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_3831),
.B(n_431),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4002),
.B(n_431),
.Y(n_4471)
);

O2A1O1Ixp33_ASAP7_75t_L g4472 ( 
.A1(n_3930),
.A2(n_433),
.B(n_434),
.C(n_432),
.Y(n_4472)
);

NOR2x2_ASAP7_75t_L g4473 ( 
.A(n_4001),
.B(n_4007),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_3836),
.B(n_432),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_3838),
.B(n_432),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_3454),
.Y(n_4476)
);

AOI22xp5_ASAP7_75t_L g4477 ( 
.A1(n_3932),
.A2(n_435),
.B1(n_436),
.B2(n_434),
.Y(n_4477)
);

AOI22xp33_ASAP7_75t_L g4478 ( 
.A1(n_3966),
.A2(n_435),
.B1(n_436),
.B2(n_434),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_SL g4479 ( 
.A(n_3999),
.B(n_3726),
.Y(n_4479)
);

OR2x6_ASAP7_75t_L g4480 ( 
.A(n_3999),
.B(n_437),
.Y(n_4480)
);

A2O1A1Ixp33_ASAP7_75t_L g4481 ( 
.A1(n_3927),
.A2(n_3498),
.B(n_3577),
.C(n_3518),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_SL g4482 ( 
.A(n_3486),
.B(n_437),
.Y(n_4482)
);

AOI22xp5_ASAP7_75t_L g4483 ( 
.A1(n_3936),
.A2(n_438),
.B1(n_439),
.B2(n_437),
.Y(n_4483)
);

AOI22xp33_ASAP7_75t_SL g4484 ( 
.A1(n_3860),
.A2(n_439),
.B1(n_440),
.B2(n_438),
.Y(n_4484)
);

AOI22xp5_ASAP7_75t_L g4485 ( 
.A1(n_3943),
.A2(n_440),
.B1(n_441),
.B2(n_439),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_SL g4486 ( 
.A(n_3745),
.B(n_440),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_3961),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_3841),
.B(n_441),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_L g4489 ( 
.A(n_3842),
.B(n_442),
.Y(n_4489)
);

BUFx6f_ASAP7_75t_L g4490 ( 
.A(n_3631),
.Y(n_4490)
);

INVx3_ASAP7_75t_L g4491 ( 
.A(n_3631),
.Y(n_4491)
);

INVx2_ASAP7_75t_L g4492 ( 
.A(n_3969),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_3460),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_3843),
.B(n_442),
.Y(n_4494)
);

AOI22xp33_ASAP7_75t_L g4495 ( 
.A1(n_3754),
.A2(n_443),
.B1(n_444),
.B2(n_442),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_3844),
.B(n_443),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_3705),
.B(n_1069),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_3462),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_3464),
.Y(n_4499)
);

AOI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_3952),
.A2(n_445),
.B(n_444),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_3469),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_3845),
.B(n_444),
.Y(n_4502)
);

AND3x1_ASAP7_75t_SL g4503 ( 
.A(n_3985),
.B(n_446),
.C(n_445),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_SL g4504 ( 
.A(n_3897),
.B(n_3824),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_SL g4505 ( 
.A(n_3830),
.B(n_445),
.Y(n_4505)
);

NAND2xp5_ASAP7_75t_SL g4506 ( 
.A(n_3851),
.B(n_446),
.Y(n_4506)
);

AND2x6_ASAP7_75t_SL g4507 ( 
.A(n_3614),
.B(n_1),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_3846),
.B(n_447),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_3850),
.B(n_448),
.Y(n_4509)
);

AND2x6_ASAP7_75t_L g4510 ( 
.A(n_4008),
.B(n_452),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_3833),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_3856),
.B(n_449),
.Y(n_4512)
);

NOR2xp33_ASAP7_75t_L g4513 ( 
.A(n_3593),
.B(n_449),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_SL g4514 ( 
.A(n_3631),
.B(n_449),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_3858),
.B(n_450),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_3484),
.Y(n_4516)
);

INVx2_ASAP7_75t_L g4517 ( 
.A(n_3833),
.Y(n_4517)
);

BUFx3_ASAP7_75t_L g4518 ( 
.A(n_3751),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_3868),
.B(n_450),
.Y(n_4519)
);

HB1xp67_ASAP7_75t_L g4520 ( 
.A(n_3613),
.Y(n_4520)
);

NOR3xp33_ASAP7_75t_L g4521 ( 
.A(n_3960),
.B(n_451),
.C(n_450),
.Y(n_4521)
);

AOI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_3538),
.A2(n_452),
.B(n_451),
.Y(n_4522)
);

AOI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_3538),
.A2(n_453),
.B(n_451),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_3719),
.B(n_1063),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_SL g4525 ( 
.A(n_3699),
.B(n_453),
.Y(n_4525)
);

AOI22xp33_ASAP7_75t_L g4526 ( 
.A1(n_3819),
.A2(n_454),
.B1(n_455),
.B2(n_453),
.Y(n_4526)
);

INVx5_ASAP7_75t_L g4527 ( 
.A(n_3699),
.Y(n_4527)
);

AOI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_3984),
.A2(n_456),
.B1(n_457),
.B2(n_454),
.Y(n_4528)
);

INVx2_ASAP7_75t_L g4529 ( 
.A(n_3905),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_3873),
.B(n_454),
.Y(n_4530)
);

INVx3_ASAP7_75t_L g4531 ( 
.A(n_3699),
.Y(n_4531)
);

INVx2_ASAP7_75t_SL g4532 ( 
.A(n_3751),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_3575),
.B(n_1066),
.Y(n_4533)
);

BUFx3_ASAP7_75t_L g4534 ( 
.A(n_3762),
.Y(n_4534)
);

AOI21xp5_ASAP7_75t_L g4535 ( 
.A1(n_3509),
.A2(n_457),
.B(n_456),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_3488),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_3490),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_3875),
.B(n_458),
.Y(n_4538)
);

NOR2xp33_ASAP7_75t_L g4539 ( 
.A(n_3595),
.B(n_458),
.Y(n_4539)
);

CKINVDCx20_ASAP7_75t_R g4540 ( 
.A(n_3688),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_3492),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_SL g4542 ( 
.A(n_3723),
.B(n_3798),
.Y(n_4542)
);

BUFx12f_ASAP7_75t_L g4543 ( 
.A(n_3723),
.Y(n_4543)
);

AOI21xp5_ASAP7_75t_L g4544 ( 
.A1(n_3723),
.A2(n_459),
.B(n_458),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_3905),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_SL g4546 ( 
.A(n_3798),
.B(n_459),
.Y(n_4546)
);

INVx2_ASAP7_75t_L g4547 ( 
.A(n_3928),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_3878),
.B(n_460),
.Y(n_4548)
);

BUFx5_ASAP7_75t_L g4549 ( 
.A(n_4013),
.Y(n_4549)
);

A2O1A1Ixp33_ASAP7_75t_SL g4550 ( 
.A1(n_3681),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_4550)
);

INVx1_ASAP7_75t_SL g4551 ( 
.A(n_3615),
.Y(n_4551)
);

O2A1O1Ixp5_ASAP7_75t_L g4552 ( 
.A1(n_3523),
.A2(n_462),
.B(n_463),
.C(n_461),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_3884),
.B(n_461),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_3885),
.B(n_461),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_3892),
.B(n_3895),
.Y(n_4555)
);

AOI21xp5_ASAP7_75t_L g4556 ( 
.A1(n_3798),
.A2(n_463),
.B(n_462),
.Y(n_4556)
);

NOR2xp33_ASAP7_75t_L g4557 ( 
.A(n_3598),
.B(n_462),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_3928),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_3896),
.B(n_463),
.Y(n_4559)
);

NAND2x1p5_ASAP7_75t_L g4560 ( 
.A(n_3762),
.B(n_467),
.Y(n_4560)
);

AND2x2_ASAP7_75t_SL g4561 ( 
.A(n_3605),
.B(n_464),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_3900),
.B(n_464),
.Y(n_4562)
);

AND2x6_ASAP7_75t_L g4563 ( 
.A(n_4008),
.B(n_467),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_3499),
.Y(n_4564)
);

INVx3_ASAP7_75t_L g4565 ( 
.A(n_3849),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_3901),
.B(n_464),
.Y(n_4566)
);

HB1xp67_ASAP7_75t_L g4567 ( 
.A(n_3805),
.Y(n_4567)
);

OR2x6_ASAP7_75t_L g4568 ( 
.A(n_3993),
.B(n_465),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_3903),
.B(n_465),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_SL g4570 ( 
.A(n_3849),
.B(n_465),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_3906),
.Y(n_4571)
);

AOI22xp33_ASAP7_75t_SL g4572 ( 
.A1(n_3860),
.A2(n_468),
.B1(n_469),
.B2(n_466),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_3576),
.B(n_1061),
.Y(n_4573)
);

INVxp67_ASAP7_75t_L g4574 ( 
.A(n_3965),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_L g4575 ( 
.A(n_3910),
.B(n_466),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_L g4576 ( 
.A(n_3916),
.B(n_3949),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_3950),
.B(n_466),
.Y(n_4577)
);

NOR2xp33_ASAP7_75t_L g4578 ( 
.A(n_3808),
.B(n_3967),
.Y(n_4578)
);

O2A1O1Ixp33_ASAP7_75t_L g4579 ( 
.A1(n_3997),
.A2(n_469),
.B(n_470),
.C(n_468),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_SL g4580 ( 
.A(n_3849),
.B(n_468),
.Y(n_4580)
);

NOR2xp33_ASAP7_75t_L g4581 ( 
.A(n_3972),
.B(n_469),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_3951),
.B(n_470),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_3956),
.B(n_3980),
.Y(n_4583)
);

INVx2_ASAP7_75t_L g4584 ( 
.A(n_3971),
.Y(n_4584)
);

HB1xp67_ASAP7_75t_L g4585 ( 
.A(n_3578),
.Y(n_4585)
);

INVx3_ASAP7_75t_L g4586 ( 
.A(n_4109),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4457),
.Y(n_4587)
);

AND2x4_ASAP7_75t_L g4588 ( 
.A(n_4322),
.B(n_4016),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4035),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4024),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4190),
.B(n_3581),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_4193),
.B(n_3582),
.Y(n_4592)
);

NOR2xp33_ASAP7_75t_L g4593 ( 
.A(n_4051),
.B(n_3793),
.Y(n_4593)
);

NAND2xp5_ASAP7_75t_SL g4594 ( 
.A(n_4075),
.B(n_3810),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4071),
.B(n_3583),
.Y(n_4595)
);

BUFx3_ASAP7_75t_L g4596 ( 
.A(n_4170),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4032),
.Y(n_4597)
);

INVx2_ASAP7_75t_L g4598 ( 
.A(n_4036),
.Y(n_4598)
);

AOI22xp5_ASAP7_75t_L g4599 ( 
.A1(n_4391),
.A2(n_4003),
.B1(n_4009),
.B2(n_4000),
.Y(n_4599)
);

AO22x1_ASAP7_75t_L g4600 ( 
.A1(n_4269),
.A2(n_3804),
.B1(n_3983),
.B2(n_3976),
.Y(n_4600)
);

BUFx6f_ASAP7_75t_L g4601 ( 
.A(n_4248),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4460),
.B(n_3825),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_4461),
.B(n_3635),
.Y(n_4603)
);

AND2x4_ASAP7_75t_L g4604 ( 
.A(n_4322),
.B(n_3804),
.Y(n_4604)
);

NOR2xp33_ASAP7_75t_R g4605 ( 
.A(n_4206),
.B(n_470),
.Y(n_4605)
);

INVx3_ASAP7_75t_L g4606 ( 
.A(n_4379),
.Y(n_4606)
);

HB1xp67_ASAP7_75t_L g4607 ( 
.A(n_4094),
.Y(n_4607)
);

BUFx2_ASAP7_75t_L g4608 ( 
.A(n_4473),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_L g4609 ( 
.A(n_4464),
.B(n_3912),
.Y(n_4609)
);

BUFx2_ASAP7_75t_L g4610 ( 
.A(n_4332),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4046),
.Y(n_4611)
);

AND2x4_ASAP7_75t_SL g4612 ( 
.A(n_4029),
.B(n_3921),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4476),
.B(n_3937),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4038),
.Y(n_4614)
);

NOR2xp67_ASAP7_75t_L g4615 ( 
.A(n_4397),
.B(n_4015),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4072),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4493),
.B(n_3511),
.Y(n_4617)
);

BUFx6f_ASAP7_75t_L g4618 ( 
.A(n_4543),
.Y(n_4618)
);

AND2x4_ASAP7_75t_L g4619 ( 
.A(n_4332),
.B(n_3818),
.Y(n_4619)
);

INVx2_ASAP7_75t_SL g4620 ( 
.A(n_4206),
.Y(n_4620)
);

BUFx2_ASAP7_75t_L g4621 ( 
.A(n_4100),
.Y(n_4621)
);

BUFx3_ASAP7_75t_L g4622 ( 
.A(n_4379),
.Y(n_4622)
);

NAND2xp33_ASAP7_75t_R g4623 ( 
.A(n_4255),
.B(n_474),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4045),
.Y(n_4624)
);

NOR3xp33_ASAP7_75t_SL g4625 ( 
.A(n_4083),
.B(n_3821),
.C(n_3758),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4498),
.B(n_3528),
.Y(n_4626)
);

AND2x4_ASAP7_75t_L g4627 ( 
.A(n_4340),
.B(n_3926),
.Y(n_4627)
);

OR2x6_ASAP7_75t_L g4628 ( 
.A(n_4399),
.B(n_3857),
.Y(n_4628)
);

BUFx6f_ASAP7_75t_L g4629 ( 
.A(n_4399),
.Y(n_4629)
);

AOI22xp5_ASAP7_75t_L g4630 ( 
.A1(n_4030),
.A2(n_3765),
.B1(n_3749),
.B2(n_3867),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4026),
.B(n_471),
.Y(n_4631)
);

BUFx6f_ASAP7_75t_L g4632 ( 
.A(n_4399),
.Y(n_4632)
);

INVx2_ASAP7_75t_L g4633 ( 
.A(n_4084),
.Y(n_4633)
);

INVx4_ASAP7_75t_L g4634 ( 
.A(n_4155),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4059),
.Y(n_4635)
);

BUFx3_ASAP7_75t_L g4636 ( 
.A(n_4152),
.Y(n_4636)
);

NOR3xp33_ASAP7_75t_SL g4637 ( 
.A(n_4169),
.B(n_3887),
.C(n_3886),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_L g4638 ( 
.A(n_4499),
.B(n_3539),
.Y(n_4638)
);

AND2x4_ASAP7_75t_L g4639 ( 
.A(n_4340),
.B(n_3552),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4501),
.B(n_4516),
.Y(n_4640)
);

AND2x4_ASAP7_75t_L g4641 ( 
.A(n_4371),
.B(n_3555),
.Y(n_4641)
);

AOI22xp33_ASAP7_75t_L g4642 ( 
.A1(n_4047),
.A2(n_3870),
.B1(n_3861),
.B2(n_3945),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4060),
.Y(n_4643)
);

AOI22xp5_ASAP7_75t_SL g4644 ( 
.A1(n_4230),
.A2(n_3934),
.B1(n_3958),
.B2(n_1065),
.Y(n_4644)
);

BUFx3_ASAP7_75t_L g4645 ( 
.A(n_4194),
.Y(n_4645)
);

INVx2_ASAP7_75t_L g4646 ( 
.A(n_4090),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4066),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4068),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4091),
.Y(n_4649)
);

AND2x4_ASAP7_75t_L g4650 ( 
.A(n_4371),
.B(n_3558),
.Y(n_4650)
);

BUFx6f_ASAP7_75t_L g4651 ( 
.A(n_4085),
.Y(n_4651)
);

OAI21xp5_ASAP7_75t_L g4652 ( 
.A1(n_4057),
.A2(n_3517),
.B(n_3466),
.Y(n_4652)
);

BUFx6f_ASAP7_75t_L g4653 ( 
.A(n_4088),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4076),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4080),
.Y(n_4655)
);

INVx3_ASAP7_75t_L g4656 ( 
.A(n_4070),
.Y(n_4656)
);

BUFx3_ASAP7_75t_L g4657 ( 
.A(n_4025),
.Y(n_4657)
);

INVx4_ASAP7_75t_L g4658 ( 
.A(n_4092),
.Y(n_4658)
);

INVx2_ASAP7_75t_SL g4659 ( 
.A(n_4041),
.Y(n_4659)
);

INVx3_ASAP7_75t_SL g4660 ( 
.A(n_4192),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4136),
.B(n_4153),
.Y(n_4661)
);

AOI22xp33_ASAP7_75t_L g4662 ( 
.A1(n_4480),
.A2(n_4394),
.B1(n_4023),
.B2(n_4300),
.Y(n_4662)
);

AOI22xp33_ASAP7_75t_SL g4663 ( 
.A1(n_4324),
.A2(n_472),
.B1(n_473),
.B2(n_471),
.Y(n_4663)
);

BUFx2_ASAP7_75t_L g4664 ( 
.A(n_4100),
.Y(n_4664)
);

AOI22xp5_ASAP7_75t_L g4665 ( 
.A1(n_4561),
.A2(n_1068),
.B1(n_1069),
.B2(n_1067),
.Y(n_4665)
);

AND2x4_ASAP7_75t_L g4666 ( 
.A(n_4044),
.B(n_472),
.Y(n_4666)
);

INVx2_ASAP7_75t_SL g4667 ( 
.A(n_4074),
.Y(n_4667)
);

AOI22xp33_ASAP7_75t_L g4668 ( 
.A1(n_4480),
.A2(n_475),
.B1(n_476),
.B2(n_474),
.Y(n_4668)
);

NAND2x1_ASAP7_75t_L g4669 ( 
.A(n_4082),
.B(n_474),
.Y(n_4669)
);

AO22x1_ASAP7_75t_L g4670 ( 
.A1(n_4269),
.A2(n_477),
.B1(n_478),
.B2(n_475),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4536),
.B(n_477),
.Y(n_4671)
);

AOI22xp5_ASAP7_75t_L g4672 ( 
.A1(n_4104),
.A2(n_1057),
.B1(n_1058),
.B2(n_1056),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_L g4673 ( 
.A(n_4537),
.B(n_478),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4196),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4197),
.Y(n_4675)
);

INVx6_ASAP7_75t_L g4676 ( 
.A(n_4053),
.Y(n_4676)
);

NOR3xp33_ASAP7_75t_SL g4677 ( 
.A(n_4198),
.B(n_479),
.C(n_478),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4215),
.Y(n_4678)
);

NAND3xp33_ASAP7_75t_L g4679 ( 
.A(n_4033),
.B(n_480),
.C(n_479),
.Y(n_4679)
);

BUFx2_ASAP7_75t_L g4680 ( 
.A(n_4100),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_4107),
.Y(n_4681)
);

OAI22xp33_ASAP7_75t_L g4682 ( 
.A1(n_4261),
.A2(n_4568),
.B1(n_4065),
.B2(n_4069),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4541),
.B(n_479),
.Y(n_4683)
);

OR2x6_ASAP7_75t_L g4684 ( 
.A(n_4029),
.B(n_480),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4140),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_SL g4686 ( 
.A(n_4021),
.B(n_480),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4150),
.Y(n_4687)
);

HB1xp67_ASAP7_75t_L g4688 ( 
.A(n_4028),
.Y(n_4688)
);

BUFx4f_ASAP7_75t_L g4689 ( 
.A(n_4290),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4564),
.B(n_481),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4034),
.B(n_481),
.Y(n_4691)
);

INVx4_ASAP7_75t_L g4692 ( 
.A(n_4070),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4224),
.Y(n_4693)
);

INVx3_ASAP7_75t_L g4694 ( 
.A(n_4117),
.Y(n_4694)
);

BUFx3_ASAP7_75t_L g4695 ( 
.A(n_4116),
.Y(n_4695)
);

CKINVDCx8_ASAP7_75t_R g4696 ( 
.A(n_4067),
.Y(n_4696)
);

AOI22xp33_ASAP7_75t_L g4697 ( 
.A1(n_4238),
.A2(n_482),
.B1(n_483),
.B2(n_481),
.Y(n_4697)
);

AND2x4_ASAP7_75t_L g4698 ( 
.A(n_4044),
.B(n_482),
.Y(n_4698)
);

INVx2_ASAP7_75t_L g4699 ( 
.A(n_4159),
.Y(n_4699)
);

BUFx6f_ASAP7_75t_L g4700 ( 
.A(n_4053),
.Y(n_4700)
);

INVxp67_ASAP7_75t_L g4701 ( 
.A(n_4323),
.Y(n_4701)
);

INVx4_ASAP7_75t_L g4702 ( 
.A(n_4117),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4243),
.Y(n_4703)
);

AND2x4_ASAP7_75t_L g4704 ( 
.A(n_4082),
.B(n_483),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4266),
.Y(n_4705)
);

INVx2_ASAP7_75t_L g4706 ( 
.A(n_4162),
.Y(n_4706)
);

INVx2_ASAP7_75t_L g4707 ( 
.A(n_4177),
.Y(n_4707)
);

NAND2xp33_ASAP7_75t_R g4708 ( 
.A(n_4348),
.B(n_1063),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4268),
.Y(n_4709)
);

AND2x2_ASAP7_75t_L g4710 ( 
.A(n_4220),
.B(n_484),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4270),
.B(n_484),
.Y(n_4711)
);

INVx1_ASAP7_75t_SL g4712 ( 
.A(n_4161),
.Y(n_4712)
);

INVx2_ASAP7_75t_SL g4713 ( 
.A(n_4027),
.Y(n_4713)
);

NOR3xp33_ASAP7_75t_SL g4714 ( 
.A(n_4247),
.B(n_485),
.C(n_484),
.Y(n_4714)
);

INVx3_ASAP7_75t_L g4715 ( 
.A(n_4397),
.Y(n_4715)
);

HB1xp67_ASAP7_75t_L g4716 ( 
.A(n_4058),
.Y(n_4716)
);

INVx3_ASAP7_75t_L g4717 ( 
.A(n_4398),
.Y(n_4717)
);

NOR3xp33_ASAP7_75t_SL g4718 ( 
.A(n_4367),
.B(n_486),
.C(n_485),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4316),
.B(n_485),
.Y(n_4719)
);

AND2x4_ASAP7_75t_L g4720 ( 
.A(n_4037),
.B(n_486),
.Y(n_4720)
);

BUFx4f_ASAP7_75t_L g4721 ( 
.A(n_4290),
.Y(n_4721)
);

AND2x4_ASAP7_75t_L g4722 ( 
.A(n_4037),
.B(n_487),
.Y(n_4722)
);

INVx5_ASAP7_75t_L g4723 ( 
.A(n_4510),
.Y(n_4723)
);

INVx3_ASAP7_75t_L g4724 ( 
.A(n_4398),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4276),
.B(n_487),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4207),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4278),
.B(n_487),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_SL g4728 ( 
.A(n_4182),
.B(n_488),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4288),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_L g4730 ( 
.A(n_4585),
.B(n_488),
.Y(n_4730)
);

BUFx6f_ASAP7_75t_L g4731 ( 
.A(n_4383),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_4289),
.B(n_488),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_SL g4733 ( 
.A(n_4172),
.B(n_4175),
.Y(n_4733)
);

INVx3_ASAP7_75t_L g4734 ( 
.A(n_4154),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4293),
.B(n_489),
.Y(n_4735)
);

NOR2xp33_ASAP7_75t_L g4736 ( 
.A(n_4237),
.B(n_489),
.Y(n_4736)
);

INVx4_ASAP7_75t_L g4737 ( 
.A(n_4134),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4303),
.B(n_489),
.Y(n_4738)
);

INVxp67_ASAP7_75t_L g4739 ( 
.A(n_4275),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4184),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4307),
.Y(n_4741)
);

BUFx10_ASAP7_75t_L g4742 ( 
.A(n_4324),
.Y(n_4742)
);

BUFx2_ASAP7_75t_L g4743 ( 
.A(n_4101),
.Y(n_4743)
);

INVx4_ASAP7_75t_L g4744 ( 
.A(n_4154),
.Y(n_4744)
);

BUFx2_ASAP7_75t_L g4745 ( 
.A(n_4101),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4308),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4315),
.Y(n_4747)
);

NOR2xp33_ASAP7_75t_L g4748 ( 
.A(n_4393),
.B(n_490),
.Y(n_4748)
);

HB1xp67_ASAP7_75t_L g4749 ( 
.A(n_4236),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4319),
.B(n_490),
.Y(n_4750)
);

BUFx2_ASAP7_75t_L g4751 ( 
.A(n_4101),
.Y(n_4751)
);

NAND3xp33_ASAP7_75t_SL g4752 ( 
.A(n_4093),
.B(n_2),
.C(n_3),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4301),
.B(n_491),
.Y(n_4753)
);

BUFx6f_ASAP7_75t_L g4754 ( 
.A(n_4392),
.Y(n_4754)
);

INVxp67_ASAP7_75t_L g4755 ( 
.A(n_4281),
.Y(n_4755)
);

INVx2_ASAP7_75t_L g4756 ( 
.A(n_4186),
.Y(n_4756)
);

AND2x4_ASAP7_75t_L g4757 ( 
.A(n_4175),
.B(n_491),
.Y(n_4757)
);

NAND2x1p5_ASAP7_75t_L g4758 ( 
.A(n_4210),
.B(n_491),
.Y(n_4758)
);

INVx3_ASAP7_75t_L g4759 ( 
.A(n_4336),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4321),
.Y(n_4760)
);

AND2x2_ASAP7_75t_L g4761 ( 
.A(n_4309),
.B(n_492),
.Y(n_4761)
);

INVx2_ASAP7_75t_SL g4762 ( 
.A(n_4282),
.Y(n_4762)
);

OR2x2_ASAP7_75t_L g4763 ( 
.A(n_4039),
.B(n_493),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4334),
.Y(n_4764)
);

INVx3_ASAP7_75t_SL g4765 ( 
.A(n_4108),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4337),
.Y(n_4766)
);

AOI22xp33_ASAP7_75t_L g4767 ( 
.A1(n_4419),
.A2(n_494),
.B1(n_495),
.B2(n_493),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_4344),
.B(n_493),
.Y(n_4768)
);

INVx3_ASAP7_75t_L g4769 ( 
.A(n_4256),
.Y(n_4769)
);

OAI221xp5_ASAP7_75t_L g4770 ( 
.A1(n_4077),
.A2(n_496),
.B1(n_497),
.B2(n_495),
.C(n_494),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4312),
.B(n_495),
.Y(n_4771)
);

INVx2_ASAP7_75t_L g4772 ( 
.A(n_4189),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4199),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4471),
.B(n_496),
.Y(n_4774)
);

INVx3_ASAP7_75t_L g4775 ( 
.A(n_4274),
.Y(n_4775)
);

CKINVDCx20_ASAP7_75t_R g4776 ( 
.A(n_4171),
.Y(n_4776)
);

INVx2_ASAP7_75t_L g4777 ( 
.A(n_4203),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4081),
.B(n_4087),
.Y(n_4778)
);

AND2x4_ASAP7_75t_L g4779 ( 
.A(n_4527),
.B(n_496),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4211),
.Y(n_4780)
);

INVx2_ASAP7_75t_L g4781 ( 
.A(n_4221),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4202),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4089),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_SL g4784 ( 
.A(n_4234),
.B(n_497),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4118),
.B(n_497),
.Y(n_4785)
);

BUFx6f_ASAP7_75t_L g4786 ( 
.A(n_4527),
.Y(n_4786)
);

AND2x4_ASAP7_75t_L g4787 ( 
.A(n_4527),
.B(n_498),
.Y(n_4787)
);

INVx5_ASAP7_75t_L g4788 ( 
.A(n_4510),
.Y(n_4788)
);

AOI22xp5_ASAP7_75t_L g4789 ( 
.A1(n_4245),
.A2(n_1062),
.B1(n_1064),
.B2(n_1061),
.Y(n_4789)
);

BUFx12f_ASAP7_75t_L g4790 ( 
.A(n_4313),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4148),
.Y(n_4791)
);

NOR2xp33_ASAP7_75t_SL g4792 ( 
.A(n_4240),
.B(n_1064),
.Y(n_4792)
);

INVx3_ASAP7_75t_L g4793 ( 
.A(n_4292),
.Y(n_4793)
);

INVx6_ASAP7_75t_L g4794 ( 
.A(n_4078),
.Y(n_4794)
);

HB1xp67_ASAP7_75t_L g4795 ( 
.A(n_4448),
.Y(n_4795)
);

NAND3xp33_ASAP7_75t_L g4796 ( 
.A(n_4484),
.B(n_499),
.C(n_498),
.Y(n_4796)
);

INVx4_ASAP7_75t_L g4797 ( 
.A(n_4328),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4156),
.B(n_498),
.Y(n_4798)
);

AOI22xp5_ASAP7_75t_L g4799 ( 
.A1(n_4124),
.A2(n_1066),
.B1(n_1067),
.B2(n_1065),
.Y(n_4799)
);

NOR2xp33_ASAP7_75t_R g4800 ( 
.A(n_4246),
.B(n_1068),
.Y(n_4800)
);

NAND2x1p5_ASAP7_75t_L g4801 ( 
.A(n_4209),
.B(n_499),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4157),
.B(n_499),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4262),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4273),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4164),
.B(n_500),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4174),
.Y(n_4806)
);

HB1xp67_ASAP7_75t_L g4807 ( 
.A(n_4179),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4183),
.B(n_4187),
.Y(n_4808)
);

INVx2_ASAP7_75t_SL g4809 ( 
.A(n_4102),
.Y(n_4809)
);

INVx3_ASAP7_75t_L g4810 ( 
.A(n_4078),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4347),
.Y(n_4811)
);

BUFx3_ASAP7_75t_L g4812 ( 
.A(n_4258),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_4287),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4357),
.Y(n_4814)
);

BUFx3_ASAP7_75t_L g4815 ( 
.A(n_4284),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4358),
.Y(n_4816)
);

CKINVDCx5p33_ASAP7_75t_R g4817 ( 
.A(n_4064),
.Y(n_4817)
);

AND2x4_ASAP7_75t_L g4818 ( 
.A(n_4133),
.B(n_500),
.Y(n_4818)
);

INVx2_ASAP7_75t_L g4819 ( 
.A(n_4317),
.Y(n_4819)
);

HB1xp67_ASAP7_75t_L g4820 ( 
.A(n_4339),
.Y(n_4820)
);

INVx2_ASAP7_75t_L g4821 ( 
.A(n_4330),
.Y(n_4821)
);

BUFx6f_ASAP7_75t_L g4822 ( 
.A(n_4133),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_SL g4823 ( 
.A(n_4353),
.B(n_501),
.Y(n_4823)
);

INVx4_ASAP7_75t_L g4824 ( 
.A(n_4208),
.Y(n_4824)
);

HB1xp67_ASAP7_75t_L g4825 ( 
.A(n_4405),
.Y(n_4825)
);

OAI21xp5_ASAP7_75t_L g4826 ( 
.A1(n_4552),
.A2(n_502),
.B(n_501),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4095),
.B(n_502),
.Y(n_4827)
);

INVx2_ASAP7_75t_L g4828 ( 
.A(n_4368),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_SL g4829 ( 
.A(n_4361),
.B(n_503),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4360),
.Y(n_4830)
);

INVx3_ASAP7_75t_L g4831 ( 
.A(n_4208),
.Y(n_4831)
);

INVx2_ASAP7_75t_L g4832 ( 
.A(n_4369),
.Y(n_4832)
);

BUFx6f_ASAP7_75t_L g4833 ( 
.A(n_4113),
.Y(n_4833)
);

INVx2_ASAP7_75t_L g4834 ( 
.A(n_4390),
.Y(n_4834)
);

AOI22xp5_ASAP7_75t_SL g4835 ( 
.A1(n_4431),
.A2(n_1058),
.B1(n_1048),
.B2(n_504),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4363),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4434),
.B(n_503),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_L g4838 ( 
.A(n_4435),
.B(n_503),
.Y(n_4838)
);

NOR2x1_ASAP7_75t_L g4839 ( 
.A(n_4049),
.B(n_4056),
.Y(n_4839)
);

OR2x2_ASAP7_75t_L g4840 ( 
.A(n_4228),
.B(n_505),
.Y(n_4840)
);

INVx4_ASAP7_75t_L g4841 ( 
.A(n_4510),
.Y(n_4841)
);

OR2x6_ASAP7_75t_L g4842 ( 
.A(n_4128),
.B(n_505),
.Y(n_4842)
);

INVx2_ASAP7_75t_SL g4843 ( 
.A(n_4376),
.Y(n_4843)
);

AO21x2_ASAP7_75t_L g4844 ( 
.A1(n_4110),
.A2(n_506),
.B(n_505),
.Y(n_4844)
);

INVx2_ASAP7_75t_L g4845 ( 
.A(n_4411),
.Y(n_4845)
);

NAND2xp5_ASAP7_75t_L g4846 ( 
.A(n_4438),
.B(n_506),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_SL g4847 ( 
.A(n_4375),
.B(n_506),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4370),
.Y(n_4848)
);

NOR2xp33_ASAP7_75t_L g4849 ( 
.A(n_4054),
.B(n_507),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4441),
.B(n_507),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4378),
.Y(n_4851)
);

A2O1A1Ixp33_ASAP7_75t_L g4852 ( 
.A1(n_4472),
.A2(n_508),
.B(n_509),
.C(n_507),
.Y(n_4852)
);

AND2x4_ASAP7_75t_L g4853 ( 
.A(n_4386),
.B(n_508),
.Y(n_4853)
);

INVx3_ASAP7_75t_L g4854 ( 
.A(n_4299),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4387),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4031),
.B(n_508),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4437),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4096),
.B(n_509),
.Y(n_4858)
);

BUFx6f_ASAP7_75t_L g4859 ( 
.A(n_4113),
.Y(n_4859)
);

INVx2_ASAP7_75t_L g4860 ( 
.A(n_4469),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4401),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4571),
.B(n_509),
.Y(n_4862)
);

AOI22xp5_ASAP7_75t_L g4863 ( 
.A1(n_4226),
.A2(n_1058),
.B1(n_1059),
.B2(n_1056),
.Y(n_4863)
);

OR2x2_ASAP7_75t_L g4864 ( 
.A(n_4112),
.B(n_510),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4406),
.Y(n_4865)
);

BUFx3_ASAP7_75t_L g4866 ( 
.A(n_4166),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4417),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_SL g4868 ( 
.A(n_4375),
.B(n_510),
.Y(n_4868)
);

HB1xp67_ASAP7_75t_L g4869 ( 
.A(n_4487),
.Y(n_4869)
);

NOR3xp33_ASAP7_75t_SL g4870 ( 
.A(n_4200),
.B(n_511),
.C(n_510),
.Y(n_4870)
);

HB1xp67_ASAP7_75t_L g4871 ( 
.A(n_4492),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4423),
.Y(n_4872)
);

INVx2_ASAP7_75t_L g4873 ( 
.A(n_4462),
.Y(n_4873)
);

AND2x2_ASAP7_75t_L g4874 ( 
.A(n_4366),
.B(n_511),
.Y(n_4874)
);

INVx2_ASAP7_75t_L g4875 ( 
.A(n_4584),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_SL g4876 ( 
.A(n_4151),
.B(n_511),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_SL g4877 ( 
.A(n_4130),
.B(n_512),
.Y(n_4877)
);

BUFx10_ASAP7_75t_L g4878 ( 
.A(n_4440),
.Y(n_4878)
);

NOR2xp33_ASAP7_75t_L g4879 ( 
.A(n_4061),
.B(n_512),
.Y(n_4879)
);

CKINVDCx5p33_ASAP7_75t_R g4880 ( 
.A(n_4181),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4389),
.B(n_512),
.Y(n_4881)
);

CKINVDCx20_ASAP7_75t_R g4882 ( 
.A(n_4540),
.Y(n_4882)
);

CKINVDCx5p33_ASAP7_75t_R g4883 ( 
.A(n_4440),
.Y(n_4883)
);

AOI22xp33_ASAP7_75t_L g4884 ( 
.A1(n_4521),
.A2(n_514),
.B1(n_515),
.B2(n_513),
.Y(n_4884)
);

INVx3_ASAP7_75t_L g4885 ( 
.A(n_4518),
.Y(n_4885)
);

AOI22xp33_ASAP7_75t_L g4886 ( 
.A1(n_4241),
.A2(n_514),
.B1(n_515),
.B2(n_513),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4272),
.Y(n_4887)
);

INVx2_ASAP7_75t_L g4888 ( 
.A(n_4329),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4052),
.B(n_513),
.Y(n_4889)
);

AOI221xp5_ASAP7_75t_L g4890 ( 
.A1(n_4513),
.A2(n_516),
.B1(n_517),
.B2(n_515),
.C(n_514),
.Y(n_4890)
);

CKINVDCx16_ASAP7_75t_R g4891 ( 
.A(n_4146),
.Y(n_4891)
);

INVx4_ASAP7_75t_L g4892 ( 
.A(n_4510),
.Y(n_4892)
);

AND2x4_ASAP7_75t_L g4893 ( 
.A(n_4386),
.B(n_516),
.Y(n_4893)
);

INVx2_ASAP7_75t_L g4894 ( 
.A(n_4333),
.Y(n_4894)
);

OR2x6_ASAP7_75t_L g4895 ( 
.A(n_4020),
.B(n_516),
.Y(n_4895)
);

INVx5_ASAP7_75t_L g4896 ( 
.A(n_4563),
.Y(n_4896)
);

CKINVDCx5p33_ASAP7_75t_R g4897 ( 
.A(n_4507),
.Y(n_4897)
);

AND2x4_ASAP7_75t_L g4898 ( 
.A(n_4447),
.B(n_517),
.Y(n_4898)
);

AOI22xp33_ASAP7_75t_L g4899 ( 
.A1(n_4244),
.A2(n_518),
.B1(n_519),
.B2(n_517),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4213),
.Y(n_4900)
);

NOR3xp33_ASAP7_75t_SL g4901 ( 
.A(n_4373),
.B(n_519),
.C(n_518),
.Y(n_4901)
);

NOR2xp33_ASAP7_75t_L g4902 ( 
.A(n_4062),
.B(n_518),
.Y(n_4902)
);

BUFx3_ASAP7_75t_L g4903 ( 
.A(n_4335),
.Y(n_4903)
);

BUFx3_ASAP7_75t_L g4904 ( 
.A(n_4123),
.Y(n_4904)
);

NAND3xp33_ASAP7_75t_SL g4905 ( 
.A(n_4267),
.B(n_2),
.C(n_3),
.Y(n_4905)
);

OR2x6_ASAP7_75t_L g4906 ( 
.A(n_4445),
.B(n_520),
.Y(n_4906)
);

OAI22xp5_ASAP7_75t_L g4907 ( 
.A1(n_4446),
.A2(n_521),
.B1(n_522),
.B2(n_520),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4333),
.Y(n_4908)
);

BUFx3_ASAP7_75t_L g4909 ( 
.A(n_4534),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4218),
.Y(n_4910)
);

INVx5_ASAP7_75t_L g4911 ( 
.A(n_4563),
.Y(n_4911)
);

HB1xp67_ASAP7_75t_L g4912 ( 
.A(n_4567),
.Y(n_4912)
);

OAI22xp5_ASAP7_75t_L g4913 ( 
.A1(n_4443),
.A2(n_522),
.B1(n_523),
.B2(n_521),
.Y(n_4913)
);

INVx2_ASAP7_75t_L g4914 ( 
.A(n_4511),
.Y(n_4914)
);

AND2x6_ASAP7_75t_L g4915 ( 
.A(n_4380),
.B(n_521),
.Y(n_4915)
);

INVx3_ASAP7_75t_L g4916 ( 
.A(n_4285),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4119),
.B(n_523),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4219),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_4022),
.B(n_524),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_4280),
.B(n_524),
.Y(n_4920)
);

NOR2xp33_ASAP7_75t_L g4921 ( 
.A(n_4063),
.B(n_524),
.Y(n_4921)
);

AOI22xp33_ASAP7_75t_L g4922 ( 
.A1(n_4428),
.A2(n_526),
.B1(n_527),
.B2(n_525),
.Y(n_4922)
);

CKINVDCx5p33_ASAP7_75t_R g4923 ( 
.A(n_4137),
.Y(n_4923)
);

INVx4_ASAP7_75t_R g4924 ( 
.A(n_4532),
.Y(n_4924)
);

NOR3xp33_ASAP7_75t_SL g4925 ( 
.A(n_4352),
.B(n_526),
.C(n_525),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_4195),
.B(n_525),
.Y(n_4926)
);

HB1xp67_ASAP7_75t_L g4927 ( 
.A(n_4520),
.Y(n_4927)
);

INVx6_ASAP7_75t_L g4928 ( 
.A(n_4447),
.Y(n_4928)
);

BUFx6f_ASAP7_75t_L g4929 ( 
.A(n_4113),
.Y(n_4929)
);

BUFx2_ASAP7_75t_SL g4930 ( 
.A(n_4563),
.Y(n_4930)
);

INVx1_ASAP7_75t_SL g4931 ( 
.A(n_4145),
.Y(n_4931)
);

AOI22xp5_ASAP7_75t_L g4932 ( 
.A1(n_4129),
.A2(n_1061),
.B1(n_1070),
.B2(n_1060),
.Y(n_4932)
);

INVx4_ASAP7_75t_L g4933 ( 
.A(n_4563),
.Y(n_4933)
);

AND2x6_ASAP7_75t_L g4934 ( 
.A(n_4227),
.B(n_527),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4225),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4229),
.Y(n_4936)
);

BUFx2_ASAP7_75t_L g4937 ( 
.A(n_4121),
.Y(n_4937)
);

HB1xp67_ASAP7_75t_L g4938 ( 
.A(n_4343),
.Y(n_4938)
);

BUFx2_ASAP7_75t_L g4939 ( 
.A(n_4121),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4279),
.B(n_527),
.Y(n_4940)
);

NOR2xp67_ASAP7_75t_L g4941 ( 
.A(n_4132),
.B(n_532),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_L g4942 ( 
.A(n_4165),
.B(n_528),
.Y(n_4942)
);

NOR3xp33_ASAP7_75t_SL g4943 ( 
.A(n_4173),
.B(n_529),
.C(n_528),
.Y(n_4943)
);

NAND2xp33_ASAP7_75t_R g4944 ( 
.A(n_4568),
.B(n_1071),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_SL g4945 ( 
.A(n_4110),
.B(n_528),
.Y(n_4945)
);

NOR3xp33_ASAP7_75t_SL g4946 ( 
.A(n_4359),
.B(n_530),
.C(n_529),
.Y(n_4946)
);

BUFx6f_ASAP7_75t_L g4947 ( 
.A(n_4121),
.Y(n_4947)
);

BUFx3_ASAP7_75t_L g4948 ( 
.A(n_4424),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_4517),
.Y(n_4949)
);

AND2x6_ASAP7_75t_L g4950 ( 
.A(n_4126),
.B(n_529),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4167),
.B(n_530),
.Y(n_4951)
);

INVx3_ASAP7_75t_L g4952 ( 
.A(n_4285),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4201),
.B(n_530),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4204),
.B(n_531),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_SL g4955 ( 
.A(n_4572),
.B(n_531),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4249),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4205),
.B(n_532),
.Y(n_4957)
);

INVxp67_ASAP7_75t_L g4958 ( 
.A(n_4114),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4250),
.Y(n_4959)
);

INVx2_ASAP7_75t_L g4960 ( 
.A(n_4529),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4551),
.B(n_532),
.Y(n_4961)
);

NOR2x1_ASAP7_75t_L g4962 ( 
.A(n_4217),
.B(n_533),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_L g4963 ( 
.A(n_4079),
.B(n_533),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4263),
.Y(n_4964)
);

BUFx2_ASAP7_75t_L g4965 ( 
.A(n_4143),
.Y(n_4965)
);

NOR2xp33_ASAP7_75t_R g4966 ( 
.A(n_4099),
.B(n_1047),
.Y(n_4966)
);

OR2x2_ASAP7_75t_L g4967 ( 
.A(n_4127),
.B(n_533),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4264),
.Y(n_4968)
);

INVx2_ASAP7_75t_L g4969 ( 
.A(n_4545),
.Y(n_4969)
);

NAND3xp33_ASAP7_75t_SL g4970 ( 
.A(n_4163),
.B(n_2),
.C(n_4),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4283),
.Y(n_4971)
);

NOR2xp33_ASAP7_75t_L g4972 ( 
.A(n_4073),
.B(n_534),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4040),
.Y(n_4973)
);

INVx1_ASAP7_75t_SL g4974 ( 
.A(n_4168),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4251),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4547),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4574),
.B(n_4578),
.Y(n_4977)
);

CKINVDCx20_ASAP7_75t_R g4978 ( 
.A(n_4231),
.Y(n_4978)
);

INVx4_ASAP7_75t_L g4979 ( 
.A(n_4445),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4120),
.B(n_534),
.Y(n_4980)
);

BUFx4f_ASAP7_75t_L g4981 ( 
.A(n_4560),
.Y(n_4981)
);

BUFx2_ASAP7_75t_L g4982 ( 
.A(n_4143),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4252),
.Y(n_4983)
);

HB1xp67_ASAP7_75t_L g4984 ( 
.A(n_4259),
.Y(n_4984)
);

INVx2_ASAP7_75t_SL g4985 ( 
.A(n_4185),
.Y(n_4985)
);

BUFx8_ASAP7_75t_L g4986 ( 
.A(n_4422),
.Y(n_4986)
);

AOI22xp5_ASAP7_75t_L g4987 ( 
.A1(n_4439),
.A2(n_1050),
.B1(n_1052),
.B2(n_1049),
.Y(n_4987)
);

NAND2xp5_ASAP7_75t_L g4988 ( 
.A(n_4403),
.B(n_534),
.Y(n_4988)
);

BUFx3_ASAP7_75t_L g4989 ( 
.A(n_4176),
.Y(n_4989)
);

INVx5_ASAP7_75t_L g4990 ( 
.A(n_4143),
.Y(n_4990)
);

INVx5_ASAP7_75t_L g4991 ( 
.A(n_4158),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4286),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4048),
.B(n_535),
.Y(n_4993)
);

INVx4_ASAP7_75t_L g4994 ( 
.A(n_4158),
.Y(n_4994)
);

BUFx12f_ASAP7_75t_L g4995 ( 
.A(n_4158),
.Y(n_4995)
);

INVxp67_ASAP7_75t_L g4996 ( 
.A(n_4042),
.Y(n_4996)
);

CKINVDCx20_ASAP7_75t_R g4997 ( 
.A(n_4235),
.Y(n_4997)
);

BUFx2_ASAP7_75t_L g4998 ( 
.A(n_4232),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4558),
.Y(n_4999)
);

OR2x4_ASAP7_75t_L g5000 ( 
.A(n_4180),
.B(n_535),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4291),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4297),
.Y(n_5002)
);

NOR2xp33_ASAP7_75t_L g5003 ( 
.A(n_4233),
.B(n_536),
.Y(n_5003)
);

INVx2_ASAP7_75t_L g5004 ( 
.A(n_4232),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_L g5005 ( 
.A(n_4138),
.B(n_536),
.Y(n_5005)
);

INVx4_ASAP7_75t_L g5006 ( 
.A(n_4232),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4139),
.B(n_537),
.Y(n_5007)
);

NOR2xp33_ASAP7_75t_L g5008 ( 
.A(n_4191),
.B(n_537),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4302),
.Y(n_5009)
);

INVx2_ASAP7_75t_SL g5010 ( 
.A(n_4188),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4314),
.Y(n_5011)
);

BUFx6f_ASAP7_75t_L g5012 ( 
.A(n_4364),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_4111),
.B(n_4533),
.Y(n_5013)
);

CKINVDCx5p33_ASAP7_75t_R g5014 ( 
.A(n_4142),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_SL g5015 ( 
.A(n_4260),
.B(n_537),
.Y(n_5015)
);

AO22x1_ASAP7_75t_L g5016 ( 
.A1(n_4239),
.A2(n_539),
.B1(n_540),
.B2(n_538),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4400),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_SL g5018 ( 
.A(n_4260),
.B(n_538),
.Y(n_5018)
);

INVx4_ASAP7_75t_L g5019 ( 
.A(n_4364),
.Y(n_5019)
);

INVx3_ASAP7_75t_L g5020 ( 
.A(n_4364),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4573),
.B(n_538),
.Y(n_5021)
);

AND2x2_ASAP7_75t_L g5022 ( 
.A(n_4106),
.B(n_539),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4404),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4395),
.Y(n_5024)
);

NOR2xp33_ASAP7_75t_L g5025 ( 
.A(n_4327),
.B(n_539),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_SL g5026 ( 
.A(n_4338),
.B(n_540),
.Y(n_5026)
);

NAND2x1p5_ASAP7_75t_L g5027 ( 
.A(n_4407),
.B(n_4306),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4365),
.B(n_540),
.Y(n_5028)
);

INVx5_ASAP7_75t_L g5029 ( 
.A(n_4490),
.Y(n_5029)
);

NOR2xp33_ASAP7_75t_L g5030 ( 
.A(n_4178),
.B(n_541),
.Y(n_5030)
);

CKINVDCx5p33_ASAP7_75t_R g5031 ( 
.A(n_4160),
.Y(n_5031)
);

INVxp67_ASAP7_75t_L g5032 ( 
.A(n_4115),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_4381),
.B(n_541),
.Y(n_5033)
);

INVx2_ASAP7_75t_SL g5034 ( 
.A(n_4222),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4135),
.Y(n_5035)
);

BUFx4f_ASAP7_75t_L g5036 ( 
.A(n_4497),
.Y(n_5036)
);

NOR3xp33_ASAP7_75t_SL g5037 ( 
.A(n_4295),
.B(n_542),
.C(n_541),
.Y(n_5037)
);

BUFx2_ASAP7_75t_L g5038 ( 
.A(n_4490),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_4555),
.B(n_542),
.Y(n_5039)
);

INVx2_ASAP7_75t_SL g5040 ( 
.A(n_4223),
.Y(n_5040)
);

BUFx2_ASAP7_75t_L g5041 ( 
.A(n_4490),
.Y(n_5041)
);

INVx2_ASAP7_75t_L g5042 ( 
.A(n_4549),
.Y(n_5042)
);

BUFx2_ASAP7_75t_L g5043 ( 
.A(n_4349),
.Y(n_5043)
);

BUFx2_ASAP7_75t_L g5044 ( 
.A(n_4491),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4409),
.Y(n_5045)
);

INVx3_ASAP7_75t_L g5046 ( 
.A(n_4491),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4414),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4415),
.Y(n_5048)
);

NOR2xp33_ASAP7_75t_L g5049 ( 
.A(n_4310),
.B(n_542),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_4416),
.Y(n_5050)
);

INVx2_ASAP7_75t_SL g5051 ( 
.A(n_4531),
.Y(n_5051)
);

INVx2_ASAP7_75t_L g5052 ( 
.A(n_4549),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4576),
.B(n_543),
.Y(n_5053)
);

HB1xp67_ASAP7_75t_L g5054 ( 
.A(n_4265),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4097),
.B(n_543),
.Y(n_5055)
);

INVx2_ASAP7_75t_SL g5056 ( 
.A(n_4531),
.Y(n_5056)
);

AND2x2_ASAP7_75t_L g5057 ( 
.A(n_4396),
.B(n_544),
.Y(n_5057)
);

INVx2_ASAP7_75t_L g5058 ( 
.A(n_4549),
.Y(n_5058)
);

BUFx6f_ASAP7_75t_L g5059 ( 
.A(n_4565),
.Y(n_5059)
);

BUFx2_ASAP7_75t_L g5060 ( 
.A(n_4565),
.Y(n_5060)
);

INVxp67_ASAP7_75t_SL g5061 ( 
.A(n_4294),
.Y(n_5061)
);

BUFx2_ASAP7_75t_L g5062 ( 
.A(n_4549),
.Y(n_5062)
);

AND2x2_ASAP7_75t_L g5063 ( 
.A(n_4458),
.B(n_544),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_4418),
.Y(n_5064)
);

INVx4_ASAP7_75t_L g5065 ( 
.A(n_4549),
.Y(n_5065)
);

NOR2xp33_ASAP7_75t_R g5066 ( 
.A(n_4105),
.B(n_544),
.Y(n_5066)
);

AOI21xp5_ASAP7_75t_L g5067 ( 
.A1(n_4895),
.A2(n_4345),
.B(n_4331),
.Y(n_5067)
);

AOI21xp5_ASAP7_75t_L g5068 ( 
.A1(n_4895),
.A2(n_4298),
.B(n_4350),
.Y(n_5068)
);

AOI21xp5_ASAP7_75t_L g5069 ( 
.A1(n_4600),
.A2(n_4043),
.B(n_4356),
.Y(n_5069)
);

NOR2xp33_ASAP7_75t_L g5070 ( 
.A(n_4897),
.B(n_4254),
.Y(n_5070)
);

INVx2_ASAP7_75t_L g5071 ( 
.A(n_4795),
.Y(n_5071)
);

A2O1A1Ixp33_ASAP7_75t_L g5072 ( 
.A1(n_4981),
.A2(n_4443),
.B(n_4579),
.C(n_4450),
.Y(n_5072)
);

AO21x1_ASAP7_75t_L g5073 ( 
.A1(n_4944),
.A2(n_4682),
.B(n_4702),
.Y(n_5073)
);

AOI21xp5_ASAP7_75t_L g5074 ( 
.A1(n_4733),
.A2(n_4479),
.B(n_4542),
.Y(n_5074)
);

HB1xp67_ASAP7_75t_L g5075 ( 
.A(n_4607),
.Y(n_5075)
);

INVxp67_ASAP7_75t_L g5076 ( 
.A(n_4601),
.Y(n_5076)
);

OAI21xp5_ASAP7_75t_L g5077 ( 
.A1(n_4941),
.A2(n_4421),
.B(n_4430),
.Y(n_5077)
);

BUFx2_ASAP7_75t_SL g5078 ( 
.A(n_4620),
.Y(n_5078)
);

OR2x6_ASAP7_75t_L g5079 ( 
.A(n_4930),
.B(n_4463),
.Y(n_5079)
);

NOR2xp33_ASAP7_75t_L g5080 ( 
.A(n_4891),
.B(n_4257),
.Y(n_5080)
);

AND2x4_ASAP7_75t_L g5081 ( 
.A(n_4608),
.B(n_4050),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_SL g5082 ( 
.A(n_4723),
.B(n_4338),
.Y(n_5082)
);

INVx2_ASAP7_75t_L g5083 ( 
.A(n_4869),
.Y(n_5083)
);

AOI21xp5_ASAP7_75t_L g5084 ( 
.A1(n_4723),
.A2(n_4896),
.B(n_4788),
.Y(n_5084)
);

AND2x2_ASAP7_75t_L g5085 ( 
.A(n_4661),
.B(n_4581),
.Y(n_5085)
);

INVx2_ASAP7_75t_L g5086 ( 
.A(n_4871),
.Y(n_5086)
);

AOI22xp5_ASAP7_75t_L g5087 ( 
.A1(n_4662),
.A2(n_4503),
.B1(n_4450),
.B2(n_4103),
.Y(n_5087)
);

AOI21xp5_ASAP7_75t_L g5088 ( 
.A1(n_4723),
.A2(n_4277),
.B(n_4354),
.Y(n_5088)
);

NOR2xp33_ASAP7_75t_L g5089 ( 
.A(n_4882),
.B(n_4271),
.Y(n_5089)
);

OAI21x1_ASAP7_75t_L g5090 ( 
.A1(n_4839),
.A2(n_4362),
.B(n_4384),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_L g5091 ( 
.A(n_4973),
.B(n_4992),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_4788),
.A2(n_4429),
.B(n_4481),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_5001),
.B(n_4539),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_4807),
.Y(n_5094)
);

BUFx3_ASAP7_75t_L g5095 ( 
.A(n_4596),
.Y(n_5095)
);

BUFx12f_ASAP7_75t_L g5096 ( 
.A(n_4618),
.Y(n_5096)
);

OAI22xp5_ASAP7_75t_L g5097 ( 
.A1(n_4906),
.A2(n_5036),
.B1(n_4608),
.B2(n_5000),
.Y(n_5097)
);

O2A1O1Ixp33_ASAP7_75t_L g5098 ( 
.A1(n_4906),
.A2(n_4342),
.B(n_4583),
.C(n_4582),
.Y(n_5098)
);

INVx2_ASAP7_75t_SL g5099 ( 
.A(n_4601),
.Y(n_5099)
);

INVxp67_ASAP7_75t_L g5100 ( 
.A(n_4715),
.Y(n_5100)
);

OR2x2_ASAP7_75t_L g5101 ( 
.A(n_4820),
.B(n_4351),
.Y(n_5101)
);

NOR2xp33_ASAP7_75t_L g5102 ( 
.A(n_5031),
.B(n_4296),
.Y(n_5102)
);

A2O1A1Ixp33_ASAP7_75t_L g5103 ( 
.A1(n_4835),
.A2(n_4122),
.B(n_4311),
.C(n_4131),
.Y(n_5103)
);

AO21x1_ASAP7_75t_L g5104 ( 
.A1(n_4792),
.A2(n_4467),
.B(n_4402),
.Y(n_5104)
);

OAI22xp5_ASAP7_75t_L g5105 ( 
.A1(n_4842),
.A2(n_4304),
.B1(n_4466),
.B2(n_4144),
.Y(n_5105)
);

OAI21xp5_ASAP7_75t_L g5106 ( 
.A1(n_4752),
.A2(n_4388),
.B(n_4410),
.Y(n_5106)
);

AOI21x1_ASAP7_75t_L g5107 ( 
.A1(n_4670),
.A2(n_4456),
.B(n_4514),
.Y(n_5107)
);

NOR2xp33_ASAP7_75t_L g5108 ( 
.A(n_4923),
.B(n_4695),
.Y(n_5108)
);

NAND2xp5_ASAP7_75t_L g5109 ( 
.A(n_5002),
.B(n_4557),
.Y(n_5109)
);

INVx2_ASAP7_75t_L g5110 ( 
.A(n_4589),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_4587),
.Y(n_5111)
);

INVx4_ASAP7_75t_L g5112 ( 
.A(n_4636),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4590),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_5009),
.B(n_4459),
.Y(n_5114)
);

CKINVDCx6p67_ASAP7_75t_R g5115 ( 
.A(n_4660),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4597),
.Y(n_5116)
);

OAI22xp5_ASAP7_75t_L g5117 ( 
.A1(n_4842),
.A2(n_4141),
.B1(n_4253),
.B2(n_4216),
.Y(n_5117)
);

AND3x4_ASAP7_75t_L g5118 ( 
.A(n_4866),
.B(n_4050),
.C(n_4412),
.Y(n_5118)
);

INVx4_ASAP7_75t_L g5119 ( 
.A(n_4645),
.Y(n_5119)
);

INVx2_ASAP7_75t_L g5120 ( 
.A(n_4598),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_4762),
.B(n_4524),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4614),
.Y(n_5122)
);

BUFx6f_ASAP7_75t_L g5123 ( 
.A(n_4629),
.Y(n_5123)
);

INVx4_ASAP7_75t_L g5124 ( 
.A(n_4657),
.Y(n_5124)
);

NAND2xp33_ASAP7_75t_L g5125 ( 
.A(n_4605),
.B(n_4408),
.Y(n_5125)
);

OR2x6_ASAP7_75t_L g5126 ( 
.A(n_4684),
.B(n_4525),
.Y(n_5126)
);

INVx8_ASAP7_75t_L g5127 ( 
.A(n_4684),
.Y(n_5127)
);

NAND2xp5_ASAP7_75t_L g5128 ( 
.A(n_5011),
.B(n_4433),
.Y(n_5128)
);

NAND2xp5_ASAP7_75t_L g5129 ( 
.A(n_4975),
.B(n_4318),
.Y(n_5129)
);

OR2x6_ASAP7_75t_SL g5130 ( 
.A(n_4817),
.B(n_4346),
.Y(n_5130)
);

BUFx4f_ASAP7_75t_L g5131 ( 
.A(n_4790),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_4983),
.B(n_4320),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_4624),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_4635),
.Y(n_5134)
);

INVxp67_ASAP7_75t_L g5135 ( 
.A(n_4717),
.Y(n_5135)
);

NAND2xp5_ASAP7_75t_SL g5136 ( 
.A(n_4788),
.B(n_4896),
.Y(n_5136)
);

AOI21xp5_ASAP7_75t_L g5137 ( 
.A1(n_4896),
.A2(n_4214),
.B(n_4355),
.Y(n_5137)
);

AND2x4_ASAP7_75t_L g5138 ( 
.A(n_4824),
.B(n_4242),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_4782),
.B(n_4325),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_4887),
.B(n_4374),
.Y(n_5140)
);

INVx5_ASAP7_75t_L g5141 ( 
.A(n_4934),
.Y(n_5141)
);

BUFx6f_ASAP7_75t_L g5142 ( 
.A(n_4629),
.Y(n_5142)
);

AOI22xp5_ASAP7_75t_L g5143 ( 
.A1(n_4970),
.A2(n_4212),
.B1(n_4506),
.B2(n_4505),
.Y(n_5143)
);

AND2x6_ASAP7_75t_L g5144 ( 
.A(n_4712),
.B(n_4385),
.Y(n_5144)
);

NAND2xp5_ASAP7_75t_L g5145 ( 
.A(n_4971),
.B(n_4377),
.Y(n_5145)
);

NAND2xp5_ASAP7_75t_SL g5146 ( 
.A(n_4911),
.B(n_4341),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_4938),
.B(n_4382),
.Y(n_5147)
);

OAI21x1_ASAP7_75t_L g5148 ( 
.A1(n_4724),
.A2(n_4055),
.B(n_4372),
.Y(n_5148)
);

NOR3xp33_ASAP7_75t_L g5149 ( 
.A(n_4905),
.B(n_4577),
.C(n_4575),
.Y(n_5149)
);

O2A1O1Ixp33_ASAP7_75t_SL g5150 ( 
.A1(n_4713),
.A2(n_4550),
.B(n_4570),
.C(n_4546),
.Y(n_5150)
);

AOI21xp5_ASAP7_75t_L g5151 ( 
.A1(n_4911),
.A2(n_4504),
.B(n_4482),
.Y(n_5151)
);

INVx2_ASAP7_75t_L g5152 ( 
.A(n_4611),
.Y(n_5152)
);

O2A1O1Ixp33_ASAP7_75t_L g5153 ( 
.A1(n_4617),
.A2(n_4149),
.B(n_4147),
.C(n_4538),
.Y(n_5153)
);

A2O1A1Ixp33_ASAP7_75t_L g5154 ( 
.A1(n_4870),
.A2(n_4305),
.B(n_4425),
.C(n_4477),
.Y(n_5154)
);

INVx2_ASAP7_75t_L g5155 ( 
.A(n_4616),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_SL g5156 ( 
.A(n_4911),
.B(n_4483),
.Y(n_5156)
);

AND2x6_ASAP7_75t_L g5157 ( 
.A(n_4853),
.B(n_4485),
.Y(n_5157)
);

AOI22xp5_ASAP7_75t_L g5158 ( 
.A1(n_5008),
.A2(n_4326),
.B1(n_4528),
.B2(n_4098),
.Y(n_5158)
);

OAI22xp5_ASAP7_75t_L g5159 ( 
.A1(n_4599),
.A2(n_4098),
.B1(n_4455),
.B2(n_4452),
.Y(n_5159)
);

NOR3xp33_ASAP7_75t_SL g5160 ( 
.A(n_4623),
.B(n_4427),
.C(n_4420),
.Y(n_5160)
);

BUFx6f_ASAP7_75t_L g5161 ( 
.A(n_4632),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4643),
.Y(n_5162)
);

O2A1O1Ixp33_ASAP7_75t_L g5163 ( 
.A1(n_4626),
.A2(n_4548),
.B(n_4553),
.C(n_4530),
.Y(n_5163)
);

INVx2_ASAP7_75t_L g5164 ( 
.A(n_4633),
.Y(n_5164)
);

BUFx2_ASAP7_75t_L g5165 ( 
.A(n_4610),
.Y(n_5165)
);

OAI22xp5_ASAP7_75t_L g5166 ( 
.A1(n_4668),
.A2(n_4465),
.B1(n_4086),
.B2(n_4436),
.Y(n_5166)
);

A2O1A1Ixp33_ASAP7_75t_L g5167 ( 
.A1(n_4901),
.A2(n_4535),
.B(n_4556),
.C(n_4544),
.Y(n_5167)
);

NAND2xp5_ASAP7_75t_SL g5168 ( 
.A(n_4765),
.B(n_4841),
.Y(n_5168)
);

INVx2_ASAP7_75t_L g5169 ( 
.A(n_4646),
.Y(n_5169)
);

AOI21xp5_ASAP7_75t_L g5170 ( 
.A1(n_4610),
.A2(n_4486),
.B(n_4580),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_4912),
.B(n_4927),
.Y(n_5171)
);

NAND2xp5_ASAP7_75t_SL g5172 ( 
.A(n_4892),
.B(n_4432),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_4640),
.B(n_4413),
.Y(n_5173)
);

BUFx6f_ASAP7_75t_L g5174 ( 
.A(n_4632),
.Y(n_5174)
);

AOI21xp5_ASAP7_75t_L g5175 ( 
.A1(n_4823),
.A2(n_4829),
.B(n_4594),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4647),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_4649),
.Y(n_5177)
);

OAI22xp5_ASAP7_75t_L g5178 ( 
.A1(n_4979),
.A2(n_4426),
.B1(n_4478),
.B2(n_4495),
.Y(n_5178)
);

OAI22xp5_ASAP7_75t_L g5179 ( 
.A1(n_4665),
.A2(n_4526),
.B1(n_4125),
.B2(n_4444),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_SL g5180 ( 
.A(n_4933),
.B(n_4966),
.Y(n_5180)
);

AOI21xp5_ASAP7_75t_L g5181 ( 
.A1(n_5062),
.A2(n_4500),
.B(n_4522),
.Y(n_5181)
);

AO22x1_ASAP7_75t_L g5182 ( 
.A1(n_4634),
.A2(n_4449),
.B1(n_4451),
.B2(n_4442),
.Y(n_5182)
);

OAI22xp33_ASAP7_75t_L g5183 ( 
.A1(n_4708),
.A2(n_4454),
.B1(n_4468),
.B2(n_4453),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_4648),
.Y(n_5184)
);

AND2x2_ASAP7_75t_L g5185 ( 
.A(n_4985),
.B(n_4),
.Y(n_5185)
);

INVx3_ASAP7_75t_L g5186 ( 
.A(n_4622),
.Y(n_5186)
);

AND2x4_ASAP7_75t_L g5187 ( 
.A(n_4822),
.B(n_4470),
.Y(n_5187)
);

AOI21xp5_ASAP7_75t_L g5188 ( 
.A1(n_5062),
.A2(n_4523),
.B(n_4475),
.Y(n_5188)
);

NOR2xp33_ASAP7_75t_L g5189 ( 
.A(n_5014),
.B(n_4474),
.Y(n_5189)
);

OAI221xp5_ASAP7_75t_L g5190 ( 
.A1(n_4630),
.A2(n_4494),
.B1(n_4496),
.B2(n_4489),
.C(n_4488),
.Y(n_5190)
);

INVx4_ASAP7_75t_L g5191 ( 
.A(n_4618),
.Y(n_5191)
);

BUFx3_ASAP7_75t_L g5192 ( 
.A(n_4731),
.Y(n_5192)
);

NAND2xp5_ASAP7_75t_L g5193 ( 
.A(n_4783),
.B(n_4791),
.Y(n_5193)
);

NOR2xp33_ASAP7_75t_R g5194 ( 
.A(n_4776),
.B(n_545),
.Y(n_5194)
);

BUFx6f_ASAP7_75t_L g5195 ( 
.A(n_4731),
.Y(n_5195)
);

AOI21xp5_ASAP7_75t_L g5196 ( 
.A1(n_5043),
.A2(n_4508),
.B(n_4502),
.Y(n_5196)
);

INVx1_ASAP7_75t_SL g5197 ( 
.A(n_4754),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_L g5198 ( 
.A(n_4806),
.B(n_4515),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_L g5199 ( 
.A(n_4900),
.B(n_4519),
.Y(n_5199)
);

OAI21x1_ASAP7_75t_L g5200 ( 
.A1(n_4694),
.A2(n_4559),
.B(n_4554),
.Y(n_5200)
);

HB1xp67_ASAP7_75t_L g5201 ( 
.A(n_4688),
.Y(n_5201)
);

OR2x6_ASAP7_75t_L g5202 ( 
.A(n_4676),
.B(n_4509),
.Y(n_5202)
);

OAI22xp5_ASAP7_75t_L g5203 ( 
.A1(n_4697),
.A2(n_4562),
.B1(n_4566),
.B2(n_4512),
.Y(n_5203)
);

AOI21xp5_ASAP7_75t_L g5204 ( 
.A1(n_5043),
.A2(n_4569),
.B(n_546),
.Y(n_5204)
);

AOI21xp5_ASAP7_75t_L g5205 ( 
.A1(n_5015),
.A2(n_546),
.B(n_545),
.Y(n_5205)
);

INVx3_ASAP7_75t_L g5206 ( 
.A(n_4586),
.Y(n_5206)
);

NOR3xp33_ASAP7_75t_L g5207 ( 
.A(n_5016),
.B(n_5),
.C(n_6),
.Y(n_5207)
);

AND2x4_ASAP7_75t_L g5208 ( 
.A(n_4822),
.B(n_545),
.Y(n_5208)
);

AOI21xp33_ASAP7_75t_L g5209 ( 
.A1(n_4679),
.A2(n_548),
.B(n_547),
.Y(n_5209)
);

NOR2xp33_ASAP7_75t_R g5210 ( 
.A(n_4883),
.B(n_547),
.Y(n_5210)
);

NOR2xp33_ASAP7_75t_L g5211 ( 
.A(n_4989),
.B(n_5),
.Y(n_5211)
);

AND2x2_ASAP7_75t_L g5212 ( 
.A(n_5010),
.B(n_5),
.Y(n_5212)
);

NOR2xp33_ASAP7_75t_L g5213 ( 
.A(n_4797),
.B(n_5),
.Y(n_5213)
);

OR2x6_ASAP7_75t_L g5214 ( 
.A(n_4676),
.B(n_547),
.Y(n_5214)
);

NOR2xp33_ASAP7_75t_R g5215 ( 
.A(n_4689),
.B(n_548),
.Y(n_5215)
);

AOI21xp5_ASAP7_75t_L g5216 ( 
.A1(n_5018),
.A2(n_550),
.B(n_549),
.Y(n_5216)
);

AOI22xp5_ASAP7_75t_L g5217 ( 
.A1(n_4593),
.A2(n_550),
.B1(n_551),
.B2(n_549),
.Y(n_5217)
);

AOI22xp5_ASAP7_75t_L g5218 ( 
.A1(n_5049),
.A2(n_550),
.B1(n_551),
.B2(n_549),
.Y(n_5218)
);

NOR2x1_ASAP7_75t_L g5219 ( 
.A(n_4658),
.B(n_551),
.Y(n_5219)
);

A2O1A1Ixp33_ASAP7_75t_L g5220 ( 
.A1(n_4615),
.A2(n_553),
.B(n_554),
.C(n_552),
.Y(n_5220)
);

OAI21xp5_ASAP7_75t_L g5221 ( 
.A1(n_4663),
.A2(n_553),
.B(n_552),
.Y(n_5221)
);

A2O1A1Ixp33_ASAP7_75t_SL g5222 ( 
.A1(n_4748),
.A2(n_554),
.B(n_555),
.C(n_553),
.Y(n_5222)
);

NOR2xp33_ASAP7_75t_L g5223 ( 
.A(n_4978),
.B(n_6),
.Y(n_5223)
);

INVx2_ASAP7_75t_L g5224 ( 
.A(n_4681),
.Y(n_5224)
);

NOR2xp33_ASAP7_75t_SL g5225 ( 
.A(n_4696),
.B(n_555),
.Y(n_5225)
);

OAI21xp33_ASAP7_75t_SL g5226 ( 
.A1(n_4692),
.A2(n_556),
.B(n_555),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_SL g5227 ( 
.A(n_5066),
.B(n_556),
.Y(n_5227)
);

AOI22xp33_ASAP7_75t_L g5228 ( 
.A1(n_4915),
.A2(n_557),
.B1(n_558),
.B2(n_556),
.Y(n_5228)
);

OAI21x1_ASAP7_75t_L g5229 ( 
.A1(n_5004),
.A2(n_558),
.B(n_557),
.Y(n_5229)
);

AOI21xp5_ASAP7_75t_L g5230 ( 
.A1(n_5026),
.A2(n_559),
.B(n_557),
.Y(n_5230)
);

AND2x2_ASAP7_75t_SL g5231 ( 
.A(n_4721),
.B(n_559),
.Y(n_5231)
);

INVx2_ASAP7_75t_L g5232 ( 
.A(n_4685),
.Y(n_5232)
);

OAI22xp5_ASAP7_75t_L g5233 ( 
.A1(n_4997),
.A2(n_561),
.B1(n_562),
.B2(n_560),
.Y(n_5233)
);

INVx2_ASAP7_75t_L g5234 ( 
.A(n_4687),
.Y(n_5234)
);

INVx2_ASAP7_75t_SL g5235 ( 
.A(n_4754),
.Y(n_5235)
);

A2O1A1Ixp33_ASAP7_75t_SL g5236 ( 
.A1(n_5003),
.A2(n_561),
.B(n_562),
.C(n_560),
.Y(n_5236)
);

AOI21xp5_ASAP7_75t_L g5237 ( 
.A1(n_5061),
.A2(n_562),
.B(n_560),
.Y(n_5237)
);

BUFx3_ASAP7_75t_L g5238 ( 
.A(n_4812),
.Y(n_5238)
);

OAI21xp5_ASAP7_75t_L g5239 ( 
.A1(n_4796),
.A2(n_564),
.B(n_563),
.Y(n_5239)
);

O2A1O1Ixp5_ASAP7_75t_SL g5240 ( 
.A1(n_4945),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_5240)
);

AND2x2_ASAP7_75t_L g5241 ( 
.A(n_5035),
.B(n_7),
.Y(n_5241)
);

O2A1O1Ixp33_ASAP7_75t_L g5242 ( 
.A1(n_4638),
.A2(n_564),
.B(n_565),
.C(n_563),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_4654),
.Y(n_5243)
);

NAND2xp5_ASAP7_75t_SL g5244 ( 
.A(n_4800),
.B(n_563),
.Y(n_5244)
);

NOR2xp33_ASAP7_75t_L g5245 ( 
.A(n_4931),
.B(n_7),
.Y(n_5245)
);

INVx2_ASAP7_75t_L g5246 ( 
.A(n_4699),
.Y(n_5246)
);

OAI22xp5_ASAP7_75t_SL g5247 ( 
.A1(n_4880),
.A2(n_566),
.B1(n_567),
.B2(n_565),
.Y(n_5247)
);

BUFx2_ASAP7_75t_L g5248 ( 
.A(n_4995),
.Y(n_5248)
);

OAI21xp5_ASAP7_75t_L g5249 ( 
.A1(n_5037),
.A2(n_567),
.B(n_566),
.Y(n_5249)
);

AOI21xp5_ASAP7_75t_L g5250 ( 
.A1(n_4652),
.A2(n_567),
.B(n_566),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_4910),
.B(n_568),
.Y(n_5251)
);

AOI21xp5_ASAP7_75t_L g5252 ( 
.A1(n_4621),
.A2(n_569),
.B(n_568),
.Y(n_5252)
);

NOR2xp33_ASAP7_75t_L g5253 ( 
.A(n_4974),
.B(n_8),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_L g5254 ( 
.A(n_4918),
.B(n_569),
.Y(n_5254)
);

BUFx6f_ASAP7_75t_L g5255 ( 
.A(n_4651),
.Y(n_5255)
);

OAI22xp5_ASAP7_75t_L g5256 ( 
.A1(n_4943),
.A2(n_4946),
.B1(n_4925),
.B2(n_4758),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_4655),
.Y(n_5257)
);

NAND2xp5_ASAP7_75t_L g5258 ( 
.A(n_4935),
.B(n_570),
.Y(n_5258)
);

CKINVDCx20_ASAP7_75t_R g5259 ( 
.A(n_4737),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_SL g5260 ( 
.A(n_4786),
.B(n_570),
.Y(n_5260)
);

NOR2xp33_ASAP7_75t_L g5261 ( 
.A(n_4986),
.B(n_8),
.Y(n_5261)
);

O2A1O1Ixp33_ASAP7_75t_L g5262 ( 
.A1(n_4988),
.A2(n_571),
.B(n_572),
.C(n_570),
.Y(n_5262)
);

AOI21xp5_ASAP7_75t_L g5263 ( 
.A1(n_4621),
.A2(n_4680),
.B(n_4664),
.Y(n_5263)
);

NOR2xp33_ASAP7_75t_L g5264 ( 
.A(n_4986),
.B(n_9),
.Y(n_5264)
);

NOR2xp33_ASAP7_75t_SL g5265 ( 
.A(n_4744),
.B(n_571),
.Y(n_5265)
);

NOR2xp33_ASAP7_75t_L g5266 ( 
.A(n_4659),
.B(n_9),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_L g5267 ( 
.A(n_4936),
.B(n_571),
.Y(n_5267)
);

NAND2xp5_ASAP7_75t_L g5268 ( 
.A(n_4956),
.B(n_573),
.Y(n_5268)
);

INVx2_ASAP7_75t_L g5269 ( 
.A(n_4706),
.Y(n_5269)
);

AND2x4_ASAP7_75t_L g5270 ( 
.A(n_4810),
.B(n_4831),
.Y(n_5270)
);

AOI21xp5_ASAP7_75t_L g5271 ( 
.A1(n_4664),
.A2(n_574),
.B(n_573),
.Y(n_5271)
);

AOI21xp5_ASAP7_75t_L g5272 ( 
.A1(n_4680),
.A2(n_574),
.B(n_573),
.Y(n_5272)
);

OAI22xp5_ASAP7_75t_L g5273 ( 
.A1(n_4612),
.A2(n_575),
.B1(n_577),
.B2(n_574),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_4959),
.B(n_575),
.Y(n_5274)
);

AOI21xp5_ASAP7_75t_L g5275 ( 
.A1(n_4743),
.A2(n_577),
.B(n_575),
.Y(n_5275)
);

NAND2xp5_ASAP7_75t_L g5276 ( 
.A(n_4964),
.B(n_577),
.Y(n_5276)
);

AO32x1_ASAP7_75t_L g5277 ( 
.A1(n_5065),
.A2(n_580),
.A3(n_581),
.B1(n_579),
.B2(n_578),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_SL g5278 ( 
.A(n_4786),
.B(n_578),
.Y(n_5278)
);

INVx3_ASAP7_75t_L g5279 ( 
.A(n_4606),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_4968),
.B(n_579),
.Y(n_5280)
);

AOI22xp5_ASAP7_75t_L g5281 ( 
.A1(n_4955),
.A2(n_580),
.B1(n_581),
.B2(n_579),
.Y(n_5281)
);

AOI21xp5_ASAP7_75t_L g5282 ( 
.A1(n_4743),
.A2(n_583),
.B(n_582),
.Y(n_5282)
);

OAI22xp5_ASAP7_75t_L g5283 ( 
.A1(n_4718),
.A2(n_585),
.B1(n_586),
.B2(n_584),
.Y(n_5283)
);

OAI22xp5_ASAP7_75t_L g5284 ( 
.A1(n_4666),
.A2(n_585),
.B1(n_586),
.B2(n_584),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_L g5285 ( 
.A(n_4811),
.B(n_4814),
.Y(n_5285)
);

OAI21xp33_ASAP7_75t_L g5286 ( 
.A1(n_4736),
.A2(n_5025),
.B(n_4879),
.Y(n_5286)
);

NOR2x1_ASAP7_75t_L g5287 ( 
.A(n_4769),
.B(n_584),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_4745),
.A2(n_586),
.B(n_585),
.Y(n_5288)
);

O2A1O1Ixp33_ASAP7_75t_L g5289 ( 
.A1(n_4980),
.A2(n_588),
.B(n_589),
.C(n_587),
.Y(n_5289)
);

BUFx8_ASAP7_75t_L g5290 ( 
.A(n_4651),
.Y(n_5290)
);

INVx1_ASAP7_75t_SL g5291 ( 
.A(n_4653),
.Y(n_5291)
);

AOI21xp5_ASAP7_75t_L g5292 ( 
.A1(n_4745),
.A2(n_588),
.B(n_587),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_4674),
.Y(n_5293)
);

NAND2xp5_ASAP7_75t_L g5294 ( 
.A(n_4816),
.B(n_4830),
.Y(n_5294)
);

INVx2_ASAP7_75t_L g5295 ( 
.A(n_4707),
.Y(n_5295)
);

NAND2xp5_ASAP7_75t_L g5296 ( 
.A(n_4836),
.B(n_589),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_4848),
.B(n_590),
.Y(n_5297)
);

OAI22xp5_ASAP7_75t_L g5298 ( 
.A1(n_4666),
.A2(n_591),
.B1(n_592),
.B2(n_590),
.Y(n_5298)
);

AOI21xp5_ASAP7_75t_L g5299 ( 
.A1(n_4751),
.A2(n_592),
.B(n_591),
.Y(n_5299)
);

OAI22xp5_ASAP7_75t_L g5300 ( 
.A1(n_4698),
.A2(n_592),
.B1(n_593),
.B2(n_591),
.Y(n_5300)
);

AOI21x1_ASAP7_75t_L g5301 ( 
.A1(n_4669),
.A2(n_594),
.B(n_593),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_4851),
.B(n_593),
.Y(n_5302)
);

OAI21x1_ASAP7_75t_L g5303 ( 
.A1(n_5027),
.A2(n_595),
.B(n_594),
.Y(n_5303)
);

INVx1_ASAP7_75t_L g5304 ( 
.A(n_4675),
.Y(n_5304)
);

INVx1_ASAP7_75t_L g5305 ( 
.A(n_4678),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_4855),
.B(n_594),
.Y(n_5306)
);

AND2x2_ASAP7_75t_SL g5307 ( 
.A(n_4700),
.B(n_595),
.Y(n_5307)
);

INVxp67_ASAP7_75t_SL g5308 ( 
.A(n_4716),
.Y(n_5308)
);

NAND2x1p5_ASAP7_75t_L g5309 ( 
.A(n_4779),
.B(n_595),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_4861),
.B(n_596),
.Y(n_5310)
);

OAI22xp5_ASAP7_75t_L g5311 ( 
.A1(n_4698),
.A2(n_597),
.B1(n_598),
.B2(n_596),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_4693),
.B(n_596),
.Y(n_5312)
);

BUFx2_ASAP7_75t_L g5313 ( 
.A(n_4909),
.Y(n_5313)
);

INVx2_ASAP7_75t_SL g5314 ( 
.A(n_4924),
.Y(n_5314)
);

BUFx6f_ASAP7_75t_L g5315 ( 
.A(n_4653),
.Y(n_5315)
);

OR2x2_ASAP7_75t_L g5316 ( 
.A(n_4726),
.B(n_597),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_4703),
.Y(n_5317)
);

NAND2xp5_ASAP7_75t_L g5318 ( 
.A(n_4705),
.B(n_598),
.Y(n_5318)
);

O2A1O1Ixp33_ASAP7_75t_L g5319 ( 
.A1(n_4942),
.A2(n_600),
.B(n_601),
.C(n_599),
.Y(n_5319)
);

AOI21xp5_ASAP7_75t_L g5320 ( 
.A1(n_4751),
.A2(n_600),
.B(n_599),
.Y(n_5320)
);

AOI21xp5_ASAP7_75t_L g5321 ( 
.A1(n_4937),
.A2(n_601),
.B(n_599),
.Y(n_5321)
);

NOR2xp33_ASAP7_75t_L g5322 ( 
.A(n_4667),
.B(n_9),
.Y(n_5322)
);

A2O1A1Ixp33_ASAP7_75t_L g5323 ( 
.A1(n_4714),
.A2(n_602),
.B(n_603),
.C(n_601),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_4709),
.B(n_602),
.Y(n_5324)
);

INVx4_ASAP7_75t_L g5325 ( 
.A(n_4948),
.Y(n_5325)
);

A2O1A1Ixp33_ASAP7_75t_L g5326 ( 
.A1(n_4677),
.A2(n_603),
.B(n_604),
.C(n_602),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_4729),
.Y(n_5327)
);

NOR2xp33_ASAP7_75t_L g5328 ( 
.A(n_4958),
.B(n_9),
.Y(n_5328)
);

BUFx6f_ASAP7_75t_L g5329 ( 
.A(n_4815),
.Y(n_5329)
);

NOR2xp33_ASAP7_75t_L g5330 ( 
.A(n_5032),
.B(n_4977),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_4741),
.B(n_4746),
.Y(n_5331)
);

INVx3_ASAP7_75t_L g5332 ( 
.A(n_4928),
.Y(n_5332)
);

BUFx2_ASAP7_75t_L g5333 ( 
.A(n_4928),
.Y(n_5333)
);

OAI22xp5_ASAP7_75t_L g5334 ( 
.A1(n_4672),
.A2(n_4757),
.B1(n_4722),
.B2(n_4720),
.Y(n_5334)
);

O2A1O1Ixp33_ASAP7_75t_L g5335 ( 
.A1(n_4951),
.A2(n_604),
.B(n_605),
.C(n_603),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_4747),
.B(n_604),
.Y(n_5336)
);

INVx2_ASAP7_75t_L g5337 ( 
.A(n_4740),
.Y(n_5337)
);

A2O1A1Ixp33_ASAP7_75t_SL g5338 ( 
.A1(n_4849),
.A2(n_606),
.B(n_607),
.C(n_605),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_L g5339 ( 
.A(n_4760),
.B(n_606),
.Y(n_5339)
);

AND2x6_ASAP7_75t_L g5340 ( 
.A(n_4853),
.B(n_606),
.Y(n_5340)
);

AOI21xp5_ASAP7_75t_L g5341 ( 
.A1(n_4937),
.A2(n_609),
.B(n_608),
.Y(n_5341)
);

BUFx2_ASAP7_75t_L g5342 ( 
.A(n_4885),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_L g5343 ( 
.A(n_4764),
.B(n_608),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_L g5344 ( 
.A(n_4766),
.B(n_608),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_4865),
.B(n_609),
.Y(n_5345)
);

INVx3_ASAP7_75t_L g5346 ( 
.A(n_4742),
.Y(n_5346)
);

OAI21xp33_ASAP7_75t_L g5347 ( 
.A1(n_4902),
.A2(n_610),
.B(n_609),
.Y(n_5347)
);

NOR2xp33_ASAP7_75t_L g5348 ( 
.A(n_4701),
.B(n_10),
.Y(n_5348)
);

INVx2_ASAP7_75t_L g5349 ( 
.A(n_4756),
.Y(n_5349)
);

NAND2xp5_ASAP7_75t_L g5350 ( 
.A(n_4867),
.B(n_610),
.Y(n_5350)
);

NAND2xp5_ASAP7_75t_SL g5351 ( 
.A(n_4700),
.B(n_610),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_4872),
.Y(n_5352)
);

BUFx2_ASAP7_75t_SL g5353 ( 
.A(n_4878),
.Y(n_5353)
);

AND2x4_ASAP7_75t_L g5354 ( 
.A(n_4904),
.B(n_611),
.Y(n_5354)
);

AOI22xp5_ASAP7_75t_L g5355 ( 
.A1(n_4642),
.A2(n_612),
.B1(n_613),
.B2(n_611),
.Y(n_5355)
);

NAND2xp5_ASAP7_75t_L g5356 ( 
.A(n_5017),
.B(n_611),
.Y(n_5356)
);

NOR2xp33_ASAP7_75t_L g5357 ( 
.A(n_4996),
.B(n_10),
.Y(n_5357)
);

INVx4_ASAP7_75t_L g5358 ( 
.A(n_4775),
.Y(n_5358)
);

HB1xp67_ASAP7_75t_L g5359 ( 
.A(n_4749),
.Y(n_5359)
);

O2A1O1Ixp33_ASAP7_75t_L g5360 ( 
.A1(n_5039),
.A2(n_613),
.B(n_614),
.C(n_612),
.Y(n_5360)
);

INVx2_ASAP7_75t_SL g5361 ( 
.A(n_4793),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_4778),
.Y(n_5362)
);

INVx2_ASAP7_75t_SL g5363 ( 
.A(n_4903),
.Y(n_5363)
);

AOI21xp5_ASAP7_75t_L g5364 ( 
.A1(n_4939),
.A2(n_616),
.B(n_615),
.Y(n_5364)
);

AOI21xp5_ASAP7_75t_L g5365 ( 
.A1(n_4939),
.A2(n_616),
.B(n_615),
.Y(n_5365)
);

NAND2xp5_ASAP7_75t_SL g5366 ( 
.A(n_4757),
.B(n_4704),
.Y(n_5366)
);

OAI21x1_ASAP7_75t_L g5367 ( 
.A1(n_4962),
.A2(n_5020),
.B(n_4801),
.Y(n_5367)
);

HB1xp67_ASAP7_75t_L g5368 ( 
.A(n_4825),
.Y(n_5368)
);

OAI21xp33_ASAP7_75t_L g5369 ( 
.A1(n_4921),
.A2(n_616),
.B(n_615),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_4808),
.Y(n_5370)
);

AND2x4_ASAP7_75t_SL g5371 ( 
.A(n_4779),
.B(n_617),
.Y(n_5371)
);

CKINVDCx14_ASAP7_75t_R g5372 ( 
.A(n_4710),
.Y(n_5372)
);

NOR2xp33_ASAP7_75t_L g5373 ( 
.A(n_4739),
.B(n_10),
.Y(n_5373)
);

NAND2xp5_ASAP7_75t_L g5374 ( 
.A(n_5023),
.B(n_617),
.Y(n_5374)
);

AOI21xp5_ASAP7_75t_L g5375 ( 
.A1(n_4965),
.A2(n_618),
.B(n_617),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_5013),
.B(n_618),
.Y(n_5376)
);

OAI22xp33_ASAP7_75t_L g5377 ( 
.A1(n_4628),
.A2(n_619),
.B1(n_620),
.B2(n_618),
.Y(n_5377)
);

O2A1O1Ixp5_ASAP7_75t_L g5378 ( 
.A1(n_4876),
.A2(n_621),
.B(n_622),
.C(n_619),
.Y(n_5378)
);

BUFx6f_ASAP7_75t_L g5379 ( 
.A(n_4833),
.Y(n_5379)
);

OAI21x1_ASAP7_75t_L g5380 ( 
.A1(n_5042),
.A2(n_621),
.B(n_619),
.Y(n_5380)
);

BUFx12f_ASAP7_75t_L g5381 ( 
.A(n_4809),
.Y(n_5381)
);

INVx4_ASAP7_75t_L g5382 ( 
.A(n_4656),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_4772),
.Y(n_5383)
);

BUFx3_ASAP7_75t_L g5384 ( 
.A(n_4843),
.Y(n_5384)
);

OAI21x1_ASAP7_75t_L g5385 ( 
.A1(n_5052),
.A2(n_622),
.B(n_621),
.Y(n_5385)
);

INVx2_ASAP7_75t_L g5386 ( 
.A(n_4773),
.Y(n_5386)
);

BUFx2_ASAP7_75t_L g5387 ( 
.A(n_4994),
.Y(n_5387)
);

HB1xp67_ASAP7_75t_L g5388 ( 
.A(n_4755),
.Y(n_5388)
);

INVx2_ASAP7_75t_L g5389 ( 
.A(n_4777),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_5071),
.B(n_5024),
.Y(n_5390)
);

A2O1A1Ixp33_ASAP7_75t_L g5391 ( 
.A1(n_5127),
.A2(n_4637),
.B(n_4625),
.C(n_4818),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_5094),
.Y(n_5392)
);

OAI21x1_ASAP7_75t_L g5393 ( 
.A1(n_5090),
.A2(n_5058),
.B(n_4952),
.Y(n_5393)
);

BUFx10_ASAP7_75t_L g5394 ( 
.A(n_5231),
.Y(n_5394)
);

NOR4xp25_ASAP7_75t_L g5395 ( 
.A(n_5097),
.B(n_5047),
.C(n_5048),
.D(n_5045),
.Y(n_5395)
);

NAND2x1p5_ASAP7_75t_L g5396 ( 
.A(n_5124),
.B(n_5112),
.Y(n_5396)
);

NOR3xp33_ASAP7_75t_SL g5397 ( 
.A(n_5168),
.B(n_4770),
.C(n_4913),
.Y(n_5397)
);

NAND3xp33_ASAP7_75t_L g5398 ( 
.A(n_5160),
.B(n_4972),
.C(n_4856),
.Y(n_5398)
);

AOI21xp5_ASAP7_75t_L g5399 ( 
.A1(n_5092),
.A2(n_4784),
.B(n_4728),
.Y(n_5399)
);

INVxp67_ASAP7_75t_SL g5400 ( 
.A(n_5165),
.Y(n_5400)
);

NAND2xp5_ASAP7_75t_L g5401 ( 
.A(n_5083),
.B(n_5050),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5193),
.Y(n_5402)
);

AOI221x1_ASAP7_75t_L g5403 ( 
.A1(n_5261),
.A2(n_5064),
.B1(n_4961),
.B2(n_4704),
.C(n_4730),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_L g5404 ( 
.A(n_5086),
.B(n_5022),
.Y(n_5404)
);

NAND2xp5_ASAP7_75t_L g5405 ( 
.A(n_5362),
.B(n_4888),
.Y(n_5405)
);

OAI21x1_ASAP7_75t_L g5406 ( 
.A1(n_5084),
.A2(n_5069),
.B(n_5148),
.Y(n_5406)
);

BUFx2_ASAP7_75t_L g5407 ( 
.A(n_5387),
.Y(n_5407)
);

INVxp67_ASAP7_75t_L g5408 ( 
.A(n_5313),
.Y(n_5408)
);

O2A1O1Ixp5_ASAP7_75t_L g5409 ( 
.A1(n_5073),
.A2(n_4787),
.B(n_4898),
.C(n_4818),
.Y(n_5409)
);

NAND2xp5_ASAP7_75t_L g5410 ( 
.A(n_5370),
.B(n_4631),
.Y(n_5410)
);

INVx1_ASAP7_75t_SL g5411 ( 
.A(n_5095),
.Y(n_5411)
);

AOI21xp5_ASAP7_75t_L g5412 ( 
.A1(n_5136),
.A2(n_4686),
.B(n_4847),
.Y(n_5412)
);

INVx2_ASAP7_75t_L g5413 ( 
.A(n_5110),
.Y(n_5413)
);

AO21x1_ASAP7_75t_L g5414 ( 
.A1(n_5244),
.A2(n_4787),
.B(n_4898),
.Y(n_5414)
);

BUFx12f_ASAP7_75t_L g5415 ( 
.A(n_5096),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5111),
.Y(n_5416)
);

NAND2xp5_ASAP7_75t_L g5417 ( 
.A(n_5075),
.B(n_4595),
.Y(n_5417)
);

NOR2xp67_ASAP7_75t_L g5418 ( 
.A(n_5314),
.B(n_4759),
.Y(n_5418)
);

AOI21x1_ASAP7_75t_L g5419 ( 
.A1(n_5182),
.A2(n_4877),
.B(n_4868),
.Y(n_5419)
);

NAND2x1p5_ASAP7_75t_L g5420 ( 
.A(n_5119),
.B(n_4720),
.Y(n_5420)
);

AO31x2_ASAP7_75t_L g5421 ( 
.A1(n_5263),
.A2(n_5060),
.A3(n_5044),
.B(n_4982),
.Y(n_5421)
);

OAI22xp5_ASAP7_75t_L g5422 ( 
.A1(n_5079),
.A2(n_4893),
.B1(n_4722),
.B2(n_4628),
.Y(n_5422)
);

AO21x2_ASAP7_75t_L g5423 ( 
.A1(n_5196),
.A2(n_4725),
.B(n_4711),
.Y(n_5423)
);

NAND3x1_ASAP7_75t_L g5424 ( 
.A(n_5264),
.B(n_4881),
.C(n_4874),
.Y(n_5424)
);

AOI22xp33_ASAP7_75t_L g5425 ( 
.A1(n_5207),
.A2(n_4915),
.B1(n_4619),
.B2(n_4934),
.Y(n_5425)
);

AO22x2_ASAP7_75t_L g5426 ( 
.A1(n_5308),
.A2(n_4893),
.B1(n_4763),
.B2(n_4840),
.Y(n_5426)
);

CKINVDCx20_ASAP7_75t_R g5427 ( 
.A(n_5290),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_SL g5428 ( 
.A(n_5141),
.B(n_4990),
.Y(n_5428)
);

AOI21xp5_ASAP7_75t_L g5429 ( 
.A1(n_5137),
.A2(n_4619),
.B(n_4965),
.Y(n_5429)
);

CKINVDCx14_ASAP7_75t_R g5430 ( 
.A(n_5372),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_5113),
.Y(n_5431)
);

NAND2x1p5_ASAP7_75t_L g5432 ( 
.A(n_5191),
.B(n_4990),
.Y(n_5432)
);

NAND3x1_ASAP7_75t_L g5433 ( 
.A(n_5108),
.B(n_5030),
.C(n_4753),
.Y(n_5433)
);

INVxp67_ASAP7_75t_SL g5434 ( 
.A(n_5359),
.Y(n_5434)
);

NAND2x1p5_ASAP7_75t_L g5435 ( 
.A(n_5325),
.B(n_4990),
.Y(n_5435)
);

OAI22xp5_ASAP7_75t_L g5436 ( 
.A1(n_5079),
.A2(n_4886),
.B1(n_4899),
.B2(n_4794),
.Y(n_5436)
);

OAI21xp5_ASAP7_75t_L g5437 ( 
.A1(n_5226),
.A2(n_4934),
.B(n_4950),
.Y(n_5437)
);

OAI21x1_ASAP7_75t_L g5438 ( 
.A1(n_5088),
.A2(n_4916),
.B(n_5046),
.Y(n_5438)
);

OAI21x1_ASAP7_75t_L g5439 ( 
.A1(n_5068),
.A2(n_5054),
.B(n_4984),
.Y(n_5439)
);

NAND2xp33_ASAP7_75t_L g5440 ( 
.A(n_5127),
.B(n_4950),
.Y(n_5440)
);

AOI21xp5_ASAP7_75t_SL g5441 ( 
.A1(n_5180),
.A2(n_4844),
.B(n_5034),
.Y(n_5441)
);

NAND2xp5_ASAP7_75t_L g5442 ( 
.A(n_5201),
.B(n_4875),
.Y(n_5442)
);

NOR2x1_ASAP7_75t_L g5443 ( 
.A(n_5358),
.B(n_5006),
.Y(n_5443)
);

A2O1A1Ixp33_ASAP7_75t_L g5444 ( 
.A1(n_5227),
.A2(n_4644),
.B(n_4863),
.C(n_4789),
.Y(n_5444)
);

OAI21x1_ASAP7_75t_SL g5445 ( 
.A1(n_5104),
.A2(n_5067),
.B(n_5334),
.Y(n_5445)
);

INVxp67_ASAP7_75t_SL g5446 ( 
.A(n_5368),
.Y(n_5446)
);

NAND2xp5_ASAP7_75t_L g5447 ( 
.A(n_5388),
.B(n_4780),
.Y(n_5447)
);

OAI21xp5_ASAP7_75t_L g5448 ( 
.A1(n_5098),
.A2(n_4950),
.B(n_4852),
.Y(n_5448)
);

CKINVDCx20_ASAP7_75t_R g5449 ( 
.A(n_5259),
.Y(n_5449)
);

AOI21xp5_ASAP7_75t_L g5450 ( 
.A1(n_5146),
.A2(n_5082),
.B(n_5172),
.Y(n_5450)
);

NAND2xp5_ASAP7_75t_L g5451 ( 
.A(n_5091),
.B(n_5171),
.Y(n_5451)
);

OR2x2_ASAP7_75t_L g5452 ( 
.A(n_5285),
.B(n_4781),
.Y(n_5452)
);

INVx3_ASAP7_75t_L g5453 ( 
.A(n_5238),
.Y(n_5453)
);

NAND2xp5_ASAP7_75t_L g5454 ( 
.A(n_5116),
.B(n_4803),
.Y(n_5454)
);

OAI21x1_ASAP7_75t_L g5455 ( 
.A1(n_5367),
.A2(n_4854),
.B(n_4914),
.Y(n_5455)
);

OA21x2_ASAP7_75t_L g5456 ( 
.A1(n_5074),
.A2(n_5060),
.B(n_5044),
.Y(n_5456)
);

INVx2_ASAP7_75t_L g5457 ( 
.A(n_5120),
.Y(n_5457)
);

OAI21x1_ASAP7_75t_L g5458 ( 
.A1(n_5151),
.A2(n_4960),
.B(n_4949),
.Y(n_5458)
);

OAI21x1_ASAP7_75t_L g5459 ( 
.A1(n_5170),
.A2(n_4976),
.B(n_4969),
.Y(n_5459)
);

AOI21x1_ASAP7_75t_L g5460 ( 
.A1(n_5366),
.A2(n_4998),
.B(n_4982),
.Y(n_5460)
);

AOI21xp5_ASAP7_75t_L g5461 ( 
.A1(n_5156),
.A2(n_5038),
.B(n_4998),
.Y(n_5461)
);

AOI21xp5_ASAP7_75t_L g5462 ( 
.A1(n_5141),
.A2(n_5041),
.B(n_5038),
.Y(n_5462)
);

AOI21xp5_ASAP7_75t_L g5463 ( 
.A1(n_5141),
.A2(n_5041),
.B(n_5051),
.Y(n_5463)
);

NAND2xp5_ASAP7_75t_L g5464 ( 
.A(n_5122),
.B(n_5133),
.Y(n_5464)
);

INVxp67_ASAP7_75t_SL g5465 ( 
.A(n_5152),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5134),
.Y(n_5466)
);

NOR2xp33_ASAP7_75t_L g5467 ( 
.A(n_5291),
.B(n_4967),
.Y(n_5467)
);

NAND2xp5_ASAP7_75t_SL g5468 ( 
.A(n_5329),
.B(n_4991),
.Y(n_5468)
);

O2A1O1Ixp5_ASAP7_75t_L g5469 ( 
.A1(n_5213),
.A2(n_5053),
.B(n_5007),
.C(n_5005),
.Y(n_5469)
);

CKINVDCx5p33_ASAP7_75t_R g5470 ( 
.A(n_5115),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5162),
.Y(n_5471)
);

NAND2xp5_ASAP7_75t_L g5472 ( 
.A(n_5176),
.B(n_4804),
.Y(n_5472)
);

NAND2xp5_ASAP7_75t_L g5473 ( 
.A(n_5184),
.B(n_4813),
.Y(n_5473)
);

AOI21xp5_ASAP7_75t_L g5474 ( 
.A1(n_5181),
.A2(n_5056),
.B(n_5040),
.Y(n_5474)
);

BUFx2_ASAP7_75t_L g5475 ( 
.A(n_5333),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_5243),
.B(n_4819),
.Y(n_5476)
);

NAND2x1p5_ASAP7_75t_L g5477 ( 
.A(n_5248),
.B(n_4991),
.Y(n_5477)
);

NAND2xp5_ASAP7_75t_L g5478 ( 
.A(n_5257),
.B(n_4821),
.Y(n_5478)
);

NOR4xp25_ASAP7_75t_L g5479 ( 
.A(n_5183),
.B(n_4993),
.C(n_4727),
.D(n_4735),
.Y(n_5479)
);

OA21x2_ASAP7_75t_L g5480 ( 
.A1(n_5200),
.A2(n_4832),
.B(n_4828),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5293),
.Y(n_5481)
);

OAI21x1_ASAP7_75t_L g5482 ( 
.A1(n_5188),
.A2(n_4999),
.B(n_4845),
.Y(n_5482)
);

INVxp67_ASAP7_75t_L g5483 ( 
.A(n_5342),
.Y(n_5483)
);

OAI21x1_ASAP7_75t_L g5484 ( 
.A1(n_5301),
.A2(n_4857),
.B(n_4834),
.Y(n_5484)
);

AOI21x1_ASAP7_75t_L g5485 ( 
.A1(n_5287),
.A2(n_4604),
.B(n_5055),
.Y(n_5485)
);

AOI21xp5_ASAP7_75t_L g5486 ( 
.A1(n_5103),
.A2(n_4627),
.B(n_4826),
.Y(n_5486)
);

NAND2xp5_ASAP7_75t_L g5487 ( 
.A(n_5304),
.B(n_4860),
.Y(n_5487)
);

OAI21xp5_ASAP7_75t_L g5488 ( 
.A1(n_5220),
.A2(n_4915),
.B(n_4932),
.Y(n_5488)
);

BUFx6f_ASAP7_75t_L g5489 ( 
.A(n_5255),
.Y(n_5489)
);

INVx2_ASAP7_75t_SL g5490 ( 
.A(n_5255),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5305),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_L g5492 ( 
.A(n_5317),
.B(n_4873),
.Y(n_5492)
);

AO31x2_ASAP7_75t_L g5493 ( 
.A1(n_5117),
.A2(n_4894),
.A3(n_4908),
.B(n_5019),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_5327),
.Y(n_5494)
);

AO31x2_ASAP7_75t_L g5495 ( 
.A1(n_5105),
.A2(n_4602),
.A3(n_4603),
.B(n_4609),
.Y(n_5495)
);

AND2x2_ASAP7_75t_L g5496 ( 
.A(n_5085),
.B(n_4719),
.Y(n_5496)
);

AND2x2_ASAP7_75t_L g5497 ( 
.A(n_5121),
.B(n_4761),
.Y(n_5497)
);

OAI21xp5_ASAP7_75t_L g5498 ( 
.A1(n_5307),
.A2(n_4987),
.B(n_5057),
.Y(n_5498)
);

OAI21x1_ASAP7_75t_L g5499 ( 
.A1(n_5175),
.A2(n_4734),
.B(n_4785),
.Y(n_5499)
);

OAI21x1_ASAP7_75t_L g5500 ( 
.A1(n_5107),
.A2(n_4802),
.B(n_4798),
.Y(n_5500)
);

AND2x6_ASAP7_75t_SL g5501 ( 
.A(n_5089),
.B(n_5063),
.Y(n_5501)
);

OAI21xp5_ASAP7_75t_L g5502 ( 
.A1(n_5323),
.A2(n_4907),
.B(n_4919),
.Y(n_5502)
);

OAI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_5326),
.A2(n_4889),
.B(n_4799),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_5352),
.B(n_4771),
.Y(n_5504)
);

AOI21xp5_ASAP7_75t_L g5505 ( 
.A1(n_5150),
.A2(n_4627),
.B(n_4604),
.Y(n_5505)
);

AOI21xp5_ASAP7_75t_L g5506 ( 
.A1(n_5072),
.A2(n_5029),
.B(n_4991),
.Y(n_5506)
);

OA22x2_ASAP7_75t_L g5507 ( 
.A1(n_5081),
.A2(n_4774),
.B1(n_4588),
.B2(n_4641),
.Y(n_5507)
);

NOR3xp33_ASAP7_75t_SL g5508 ( 
.A(n_5247),
.B(n_4890),
.C(n_5021),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5294),
.Y(n_5509)
);

BUFx2_ASAP7_75t_L g5510 ( 
.A(n_5100),
.Y(n_5510)
);

NAND2xp5_ASAP7_75t_L g5511 ( 
.A(n_5101),
.B(n_4864),
.Y(n_5511)
);

NOR2xp33_ASAP7_75t_SL g5512 ( 
.A(n_5131),
.B(n_4794),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5155),
.Y(n_5513)
);

NOR2x1_ASAP7_75t_SL g5514 ( 
.A(n_5078),
.B(n_5029),
.Y(n_5514)
);

BUFx3_ASAP7_75t_L g5515 ( 
.A(n_5329),
.Y(n_5515)
);

AOI21xp5_ASAP7_75t_L g5516 ( 
.A1(n_5138),
.A2(n_5135),
.B(n_5077),
.Y(n_5516)
);

BUFx2_ASAP7_75t_L g5517 ( 
.A(n_5382),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_5331),
.Y(n_5518)
);

OAI21x1_ASAP7_75t_L g5519 ( 
.A1(n_5380),
.A2(n_4805),
.B(n_4738),
.Y(n_5519)
);

O2A1O1Ixp5_ASAP7_75t_SL g5520 ( 
.A1(n_5076),
.A2(n_4926),
.B(n_4750),
.C(n_4732),
.Y(n_5520)
);

OAI21x1_ASAP7_75t_SL g5521 ( 
.A1(n_5219),
.A2(n_4768),
.B(n_4862),
.Y(n_5521)
);

AOI21xp5_ASAP7_75t_L g5522 ( 
.A1(n_5125),
.A2(n_5029),
.B(n_4641),
.Y(n_5522)
);

AOI21xp5_ASAP7_75t_L g5523 ( 
.A1(n_5236),
.A2(n_4650),
.B(n_4639),
.Y(n_5523)
);

OAI21x1_ASAP7_75t_L g5524 ( 
.A1(n_5385),
.A2(n_5229),
.B(n_5303),
.Y(n_5524)
);

INVx3_ASAP7_75t_L g5525 ( 
.A(n_5315),
.Y(n_5525)
);

CKINVDCx11_ASAP7_75t_R g5526 ( 
.A(n_5381),
.Y(n_5526)
);

AOI21xp5_ASAP7_75t_L g5527 ( 
.A1(n_5338),
.A2(n_4650),
.B(n_4639),
.Y(n_5527)
);

INVx2_ASAP7_75t_SL g5528 ( 
.A(n_5315),
.Y(n_5528)
);

OAI22xp5_ASAP7_75t_L g5529 ( 
.A1(n_5118),
.A2(n_4884),
.B1(n_4767),
.B2(n_4613),
.Y(n_5529)
);

OAI22xp5_ASAP7_75t_L g5530 ( 
.A1(n_5228),
.A2(n_4922),
.B1(n_4588),
.B2(n_4592),
.Y(n_5530)
);

AOI21xp5_ASAP7_75t_L g5531 ( 
.A1(n_5126),
.A2(n_4940),
.B(n_4917),
.Y(n_5531)
);

AOI21xp5_ASAP7_75t_L g5532 ( 
.A1(n_5126),
.A2(n_4691),
.B(n_4833),
.Y(n_5532)
);

AOI21xp5_ASAP7_75t_L g5533 ( 
.A1(n_5256),
.A2(n_4929),
.B(n_4859),
.Y(n_5533)
);

OAI21x1_ASAP7_75t_L g5534 ( 
.A1(n_5204),
.A2(n_4591),
.B(n_4671),
.Y(n_5534)
);

NAND2xp5_ASAP7_75t_L g5535 ( 
.A(n_5383),
.B(n_4858),
.Y(n_5535)
);

OR2x2_ASAP7_75t_L g5536 ( 
.A(n_5164),
.B(n_5169),
.Y(n_5536)
);

OAI21x1_ASAP7_75t_L g5537 ( 
.A1(n_5332),
.A2(n_4683),
.B(n_4673),
.Y(n_5537)
);

OA21x2_ASAP7_75t_L g5538 ( 
.A1(n_5128),
.A2(n_4690),
.B(n_4837),
.Y(n_5538)
);

INVx2_ASAP7_75t_L g5539 ( 
.A(n_5177),
.Y(n_5539)
);

OAI21x1_ASAP7_75t_L g5540 ( 
.A1(n_5309),
.A2(n_4846),
.B(n_4838),
.Y(n_5540)
);

A2O1A1Ixp33_ASAP7_75t_L g5541 ( 
.A1(n_5347),
.A2(n_4963),
.B(n_4827),
.C(n_5028),
.Y(n_5541)
);

AOI21x1_ASAP7_75t_L g5542 ( 
.A1(n_5260),
.A2(n_4850),
.B(n_4953),
.Y(n_5542)
);

AO31x2_ASAP7_75t_L g5543 ( 
.A1(n_5224),
.A2(n_4920),
.A3(n_4957),
.B(n_4954),
.Y(n_5543)
);

OAI21x1_ASAP7_75t_SL g5544 ( 
.A1(n_5363),
.A2(n_5033),
.B(n_623),
.Y(n_5544)
);

OAI21x1_ASAP7_75t_SL g5545 ( 
.A1(n_5361),
.A2(n_623),
.B(n_622),
.Y(n_5545)
);

NAND2x1_ASAP7_75t_L g5546 ( 
.A(n_5340),
.B(n_4859),
.Y(n_5546)
);

OAI21xp5_ASAP7_75t_L g5547 ( 
.A1(n_5242),
.A2(n_625),
.B(n_624),
.Y(n_5547)
);

BUFx24_ASAP7_75t_L g5548 ( 
.A(n_5354),
.Y(n_5548)
);

OAI21xp33_ASAP7_75t_L g5549 ( 
.A1(n_5194),
.A2(n_5059),
.B(n_4947),
.Y(n_5549)
);

AOI21xp5_ASAP7_75t_L g5550 ( 
.A1(n_5222),
.A2(n_4947),
.B(n_4929),
.Y(n_5550)
);

OAI21xp5_ASAP7_75t_L g5551 ( 
.A1(n_5265),
.A2(n_625),
.B(n_624),
.Y(n_5551)
);

NAND2xp5_ASAP7_75t_L g5552 ( 
.A(n_5139),
.B(n_5059),
.Y(n_5552)
);

A2O1A1Ixp33_ASAP7_75t_L g5553 ( 
.A1(n_5369),
.A2(n_5012),
.B(n_626),
.C(n_627),
.Y(n_5553)
);

OA21x2_ASAP7_75t_L g5554 ( 
.A1(n_5198),
.A2(n_5012),
.B(n_1050),
.Y(n_5554)
);

NOR2xp67_ASAP7_75t_SL g5555 ( 
.A(n_5353),
.B(n_5195),
.Y(n_5555)
);

AOI21xp5_ASAP7_75t_L g5556 ( 
.A1(n_5202),
.A2(n_5159),
.B(n_5239),
.Y(n_5556)
);

NAND2xp5_ASAP7_75t_L g5557 ( 
.A(n_5129),
.B(n_625),
.Y(n_5557)
);

AOI21xp5_ASAP7_75t_L g5558 ( 
.A1(n_5202),
.A2(n_627),
.B(n_626),
.Y(n_5558)
);

HB1xp67_ASAP7_75t_L g5559 ( 
.A(n_5232),
.Y(n_5559)
);

OR2x2_ASAP7_75t_L g5560 ( 
.A(n_5234),
.B(n_626),
.Y(n_5560)
);

AOI21x1_ASAP7_75t_L g5561 ( 
.A1(n_5278),
.A2(n_628),
.B(n_627),
.Y(n_5561)
);

O2A1O1Ixp5_ASAP7_75t_L g5562 ( 
.A1(n_5233),
.A2(n_629),
.B(n_630),
.C(n_628),
.Y(n_5562)
);

NAND2xp5_ASAP7_75t_L g5563 ( 
.A(n_5132),
.B(n_628),
.Y(n_5563)
);

AND2x2_ASAP7_75t_L g5564 ( 
.A(n_5246),
.B(n_629),
.Y(n_5564)
);

OAI21xp5_ASAP7_75t_L g5565 ( 
.A1(n_5221),
.A2(n_631),
.B(n_630),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_L g5566 ( 
.A(n_5147),
.B(n_631),
.Y(n_5566)
);

AOI221xp5_ASAP7_75t_SL g5567 ( 
.A1(n_5286),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.C(n_13),
.Y(n_5567)
);

OAI21xp5_ASAP7_75t_L g5568 ( 
.A1(n_5378),
.A2(n_632),
.B(n_631),
.Y(n_5568)
);

OAI21x1_ASAP7_75t_L g5569 ( 
.A1(n_5240),
.A2(n_633),
.B(n_632),
.Y(n_5569)
);

INVx2_ASAP7_75t_L g5570 ( 
.A(n_5269),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_SL g5571 ( 
.A(n_5195),
.B(n_632),
.Y(n_5571)
);

AO31x2_ASAP7_75t_L g5572 ( 
.A1(n_5295),
.A2(n_5337),
.A3(n_5386),
.B(n_5349),
.Y(n_5572)
);

NAND2xp5_ASAP7_75t_L g5573 ( 
.A(n_5145),
.B(n_633),
.Y(n_5573)
);

OAI21xp5_ASAP7_75t_L g5574 ( 
.A1(n_5289),
.A2(n_635),
.B(n_634),
.Y(n_5574)
);

OAI21xp5_ASAP7_75t_L g5575 ( 
.A1(n_5262),
.A2(n_636),
.B(n_634),
.Y(n_5575)
);

AOI21xp5_ASAP7_75t_L g5576 ( 
.A1(n_5106),
.A2(n_637),
.B(n_636),
.Y(n_5576)
);

OAI21x1_ASAP7_75t_SL g5577 ( 
.A1(n_5099),
.A2(n_637),
.B(n_636),
.Y(n_5577)
);

INVxp67_ASAP7_75t_SL g5578 ( 
.A(n_5389),
.Y(n_5578)
);

AO21x2_ASAP7_75t_L g5579 ( 
.A1(n_5296),
.A2(n_639),
.B(n_638),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5316),
.Y(n_5580)
);

BUFx10_ASAP7_75t_L g5581 ( 
.A(n_5371),
.Y(n_5581)
);

OAI21x1_ASAP7_75t_L g5582 ( 
.A1(n_5250),
.A2(n_639),
.B(n_638),
.Y(n_5582)
);

NOR2xp33_ASAP7_75t_R g5583 ( 
.A(n_5225),
.B(n_11),
.Y(n_5583)
);

O2A1O1Ixp5_ASAP7_75t_SL g5584 ( 
.A1(n_5346),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_5584)
);

OAI21x1_ASAP7_75t_L g5585 ( 
.A1(n_5237),
.A2(n_639),
.B(n_638),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_L g5586 ( 
.A(n_5199),
.B(n_640),
.Y(n_5586)
);

OAI22xp33_ASAP7_75t_L g5587 ( 
.A1(n_5507),
.A2(n_5214),
.B1(n_5130),
.B2(n_5087),
.Y(n_5587)
);

AOI21xp5_ASAP7_75t_L g5588 ( 
.A1(n_5440),
.A2(n_5277),
.B(n_5214),
.Y(n_5588)
);

A2O1A1Ixp33_ASAP7_75t_L g5589 ( 
.A1(n_5409),
.A2(n_5211),
.B(n_5080),
.C(n_5245),
.Y(n_5589)
);

NAND2xp5_ASAP7_75t_L g5590 ( 
.A(n_5495),
.B(n_5241),
.Y(n_5590)
);

A2O1A1Ixp33_ASAP7_75t_L g5591 ( 
.A1(n_5549),
.A2(n_5253),
.B(n_5223),
.C(n_5266),
.Y(n_5591)
);

OAI21x1_ASAP7_75t_L g5592 ( 
.A1(n_5460),
.A2(n_5206),
.B(n_5297),
.Y(n_5592)
);

CKINVDCx5p33_ASAP7_75t_R g5593 ( 
.A(n_5427),
.Y(n_5593)
);

AND2x2_ASAP7_75t_L g5594 ( 
.A(n_5407),
.B(n_5384),
.Y(n_5594)
);

NOR2xp33_ASAP7_75t_L g5595 ( 
.A(n_5430),
.B(n_5197),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5572),
.Y(n_5596)
);

NAND3xp33_ASAP7_75t_SL g5597 ( 
.A(n_5583),
.B(n_5215),
.C(n_5210),
.Y(n_5597)
);

AND2x2_ASAP7_75t_L g5598 ( 
.A(n_5434),
.B(n_5446),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5572),
.Y(n_5599)
);

AOI21xp5_ASAP7_75t_L g5600 ( 
.A1(n_5437),
.A2(n_5277),
.B(n_5319),
.Y(n_5600)
);

AOI22xp33_ASAP7_75t_L g5601 ( 
.A1(n_5445),
.A2(n_5157),
.B1(n_5340),
.B2(n_5144),
.Y(n_5601)
);

CKINVDCx16_ASAP7_75t_R g5602 ( 
.A(n_5415),
.Y(n_5602)
);

INVx2_ASAP7_75t_L g5603 ( 
.A(n_5572),
.Y(n_5603)
);

A2O1A1Ixp33_ASAP7_75t_L g5604 ( 
.A1(n_5391),
.A2(n_5322),
.B(n_5348),
.C(n_5102),
.Y(n_5604)
);

NAND2xp5_ASAP7_75t_L g5605 ( 
.A(n_5495),
.B(n_5140),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5464),
.Y(n_5606)
);

NAND2xp5_ASAP7_75t_L g5607 ( 
.A(n_5495),
.B(n_5330),
.Y(n_5607)
);

NAND2xp5_ASAP7_75t_L g5608 ( 
.A(n_5402),
.B(n_5093),
.Y(n_5608)
);

BUFx10_ASAP7_75t_L g5609 ( 
.A(n_5470),
.Y(n_5609)
);

BUFx4_ASAP7_75t_SL g5610 ( 
.A(n_5449),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5416),
.Y(n_5611)
);

AOI21xp5_ASAP7_75t_L g5612 ( 
.A1(n_5546),
.A2(n_5335),
.B(n_5360),
.Y(n_5612)
);

A2O1A1Ixp33_ASAP7_75t_SL g5613 ( 
.A1(n_5551),
.A2(n_5328),
.B(n_5357),
.C(n_5373),
.Y(n_5613)
);

OAI21xp5_ASAP7_75t_L g5614 ( 
.A1(n_5424),
.A2(n_5340),
.B(n_5273),
.Y(n_5614)
);

BUFx2_ASAP7_75t_L g5615 ( 
.A(n_5517),
.Y(n_5615)
);

OAI211xp5_ASAP7_75t_SL g5616 ( 
.A1(n_5556),
.A2(n_5469),
.B(n_5444),
.C(n_5448),
.Y(n_5616)
);

OAI21xp5_ASAP7_75t_L g5617 ( 
.A1(n_5433),
.A2(n_5249),
.B(n_5284),
.Y(n_5617)
);

AOI22xp33_ASAP7_75t_L g5618 ( 
.A1(n_5414),
.A2(n_5157),
.B1(n_5144),
.B2(n_5149),
.Y(n_5618)
);

INVxp67_ASAP7_75t_SL g5619 ( 
.A(n_5559),
.Y(n_5619)
);

NOR2xp33_ASAP7_75t_L g5620 ( 
.A(n_5515),
.B(n_5192),
.Y(n_5620)
);

AOI21xp5_ASAP7_75t_L g5621 ( 
.A1(n_5441),
.A2(n_5428),
.B(n_5506),
.Y(n_5621)
);

O2A1O1Ixp33_ASAP7_75t_L g5622 ( 
.A1(n_5541),
.A2(n_5154),
.B(n_5351),
.C(n_5283),
.Y(n_5622)
);

AOI21xp5_ASAP7_75t_L g5623 ( 
.A1(n_5474),
.A2(n_5377),
.B(n_5209),
.Y(n_5623)
);

OAI21x1_ASAP7_75t_L g5624 ( 
.A1(n_5406),
.A2(n_5306),
.B(n_5302),
.Y(n_5624)
);

OR2x2_ASAP7_75t_L g5625 ( 
.A(n_5536),
.B(n_5109),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5431),
.Y(n_5626)
);

HB1xp67_ASAP7_75t_L g5627 ( 
.A(n_5465),
.Y(n_5627)
);

O2A1O1Ixp33_ASAP7_75t_SL g5628 ( 
.A1(n_5548),
.A2(n_5235),
.B(n_5186),
.C(n_5298),
.Y(n_5628)
);

O2A1O1Ixp33_ASAP7_75t_SL g5629 ( 
.A1(n_5411),
.A2(n_5300),
.B(n_5311),
.C(n_5070),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_L g5630 ( 
.A(n_5509),
.B(n_5114),
.Y(n_5630)
);

NAND2x1p5_ASAP7_75t_L g5631 ( 
.A(n_5555),
.B(n_5123),
.Y(n_5631)
);

NOR3xp33_ASAP7_75t_L g5632 ( 
.A(n_5398),
.B(n_5190),
.C(n_5163),
.Y(n_5632)
);

INVx1_ASAP7_75t_SL g5633 ( 
.A(n_5396),
.Y(n_5633)
);

AO21x2_ASAP7_75t_L g5634 ( 
.A1(n_5395),
.A2(n_5312),
.B(n_5310),
.Y(n_5634)
);

A2O1A1Ixp33_ASAP7_75t_L g5635 ( 
.A1(n_5418),
.A2(n_5143),
.B(n_5212),
.C(n_5185),
.Y(n_5635)
);

O2A1O1Ixp33_ASAP7_75t_SL g5636 ( 
.A1(n_5408),
.A2(n_5376),
.B(n_5189),
.C(n_5218),
.Y(n_5636)
);

AO31x2_ASAP7_75t_L g5637 ( 
.A1(n_5450),
.A2(n_5324),
.A3(n_5336),
.B(n_5318),
.Y(n_5637)
);

AOI22xp5_ASAP7_75t_L g5638 ( 
.A1(n_5529),
.A2(n_5144),
.B1(n_5157),
.B2(n_5178),
.Y(n_5638)
);

BUFx12f_ASAP7_75t_L g5639 ( 
.A(n_5526),
.Y(n_5639)
);

AOI21xp5_ASAP7_75t_L g5640 ( 
.A1(n_5505),
.A2(n_5271),
.B(n_5252),
.Y(n_5640)
);

INVx2_ASAP7_75t_L g5641 ( 
.A(n_5413),
.Y(n_5641)
);

OAI22xp5_ASAP7_75t_L g5642 ( 
.A1(n_5425),
.A2(n_5158),
.B1(n_5270),
.B2(n_5208),
.Y(n_5642)
);

AOI21xp5_ASAP7_75t_L g5643 ( 
.A1(n_5522),
.A2(n_5275),
.B(n_5272),
.Y(n_5643)
);

AO22x1_ASAP7_75t_L g5644 ( 
.A1(n_5400),
.A2(n_5142),
.B1(n_5161),
.B2(n_5123),
.Y(n_5644)
);

AOI21xp5_ASAP7_75t_L g5645 ( 
.A1(n_5422),
.A2(n_5288),
.B(n_5282),
.Y(n_5645)
);

A2O1A1Ixp33_ASAP7_75t_L g5646 ( 
.A1(n_5516),
.A2(n_5532),
.B(n_5443),
.C(n_5567),
.Y(n_5646)
);

AND2x4_ASAP7_75t_L g5647 ( 
.A(n_5578),
.B(n_5379),
.Y(n_5647)
);

A2O1A1Ixp33_ASAP7_75t_L g5648 ( 
.A1(n_5558),
.A2(n_5292),
.B(n_5320),
.C(n_5299),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_5518),
.B(n_5580),
.Y(n_5649)
);

AOI22xp33_ASAP7_75t_L g5650 ( 
.A1(n_5488),
.A2(n_5179),
.B1(n_5187),
.B2(n_5166),
.Y(n_5650)
);

O2A1O1Ixp33_ASAP7_75t_L g5651 ( 
.A1(n_5521),
.A2(n_5153),
.B(n_5374),
.C(n_5356),
.Y(n_5651)
);

AOI221x1_ASAP7_75t_L g5652 ( 
.A1(n_5453),
.A2(n_5279),
.B1(n_5343),
.B2(n_5344),
.C(n_5339),
.Y(n_5652)
);

NAND2x1p5_ASAP7_75t_L g5653 ( 
.A(n_5468),
.B(n_5142),
.Y(n_5653)
);

INVx6_ASAP7_75t_SL g5654 ( 
.A(n_5581),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_5457),
.Y(n_5655)
);

O2A1O1Ixp5_ASAP7_75t_L g5656 ( 
.A1(n_5419),
.A2(n_5254),
.B(n_5258),
.C(n_5251),
.Y(n_5656)
);

O2A1O1Ixp33_ASAP7_75t_SL g5657 ( 
.A1(n_5483),
.A2(n_5167),
.B(n_5268),
.C(n_5267),
.Y(n_5657)
);

INVx2_ASAP7_75t_L g5658 ( 
.A(n_5513),
.Y(n_5658)
);

AOI221x1_ASAP7_75t_L g5659 ( 
.A1(n_5531),
.A2(n_5426),
.B1(n_5533),
.B2(n_5486),
.C(n_5525),
.Y(n_5659)
);

BUFx6f_ASAP7_75t_L g5660 ( 
.A(n_5489),
.Y(n_5660)
);

A2O1A1Ixp33_ASAP7_75t_L g5661 ( 
.A1(n_5498),
.A2(n_5341),
.B(n_5364),
.C(n_5321),
.Y(n_5661)
);

OAI21xp5_ASAP7_75t_L g5662 ( 
.A1(n_5562),
.A2(n_5375),
.B(n_5365),
.Y(n_5662)
);

O2A1O1Ixp33_ASAP7_75t_L g5663 ( 
.A1(n_5545),
.A2(n_5544),
.B(n_5553),
.C(n_5479),
.Y(n_5663)
);

O2A1O1Ixp33_ASAP7_75t_L g5664 ( 
.A1(n_5577),
.A2(n_5575),
.B(n_5574),
.C(n_5571),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_5466),
.Y(n_5665)
);

NOR2xp33_ASAP7_75t_L g5666 ( 
.A(n_5501),
.B(n_5161),
.Y(n_5666)
);

AOI21xp5_ASAP7_75t_L g5667 ( 
.A1(n_5463),
.A2(n_5514),
.B(n_5429),
.Y(n_5667)
);

BUFx12f_ASAP7_75t_L g5668 ( 
.A(n_5394),
.Y(n_5668)
);

AOI21xp5_ASAP7_75t_L g5669 ( 
.A1(n_5462),
.A2(n_5216),
.B(n_5205),
.Y(n_5669)
);

OR2x2_ASAP7_75t_SL g5670 ( 
.A(n_5456),
.B(n_5174),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_5471),
.Y(n_5671)
);

A2O1A1Ixp33_ASAP7_75t_L g5672 ( 
.A1(n_5512),
.A2(n_5230),
.B(n_5217),
.C(n_5281),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_5481),
.Y(n_5673)
);

OAI21xp5_ASAP7_75t_L g5674 ( 
.A1(n_5403),
.A2(n_5355),
.B(n_5276),
.Y(n_5674)
);

A2O1A1Ixp33_ASAP7_75t_L g5675 ( 
.A1(n_5576),
.A2(n_5280),
.B(n_5274),
.C(n_5174),
.Y(n_5675)
);

NOR2xp33_ASAP7_75t_L g5676 ( 
.A(n_5510),
.B(n_5345),
.Y(n_5676)
);

INVx1_ASAP7_75t_SL g5677 ( 
.A(n_5475),
.Y(n_5677)
);

AOI21xp5_ASAP7_75t_L g5678 ( 
.A1(n_5461),
.A2(n_5350),
.B(n_5173),
.Y(n_5678)
);

INVx2_ASAP7_75t_L g5679 ( 
.A(n_5539),
.Y(n_5679)
);

OAI222xp33_ASAP7_75t_L g5680 ( 
.A1(n_5420),
.A2(n_5203),
.B1(n_5379),
.B2(n_643),
.C1(n_641),
.C2(n_644),
.Y(n_5680)
);

O2A1O1Ixp33_ASAP7_75t_L g5681 ( 
.A1(n_5547),
.A2(n_642),
.B(n_643),
.C(n_640),
.Y(n_5681)
);

AOI21xp5_ASAP7_75t_L g5682 ( 
.A1(n_5399),
.A2(n_643),
.B(n_642),
.Y(n_5682)
);

AOI21xp5_ASAP7_75t_L g5683 ( 
.A1(n_5550),
.A2(n_644),
.B(n_642),
.Y(n_5683)
);

OAI21xp5_ASAP7_75t_L g5684 ( 
.A1(n_5520),
.A2(n_11),
.B(n_12),
.Y(n_5684)
);

NOR2xp33_ASAP7_75t_SL g5685 ( 
.A(n_5435),
.B(n_645),
.Y(n_5685)
);

AOI21xp5_ASAP7_75t_L g5686 ( 
.A1(n_5554),
.A2(n_646),
.B(n_645),
.Y(n_5686)
);

AOI221xp5_ASAP7_75t_L g5687 ( 
.A1(n_5426),
.A2(n_5392),
.B1(n_5566),
.B2(n_5586),
.C(n_5573),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_5491),
.Y(n_5688)
);

OAI21x1_ASAP7_75t_L g5689 ( 
.A1(n_5439),
.A2(n_646),
.B(n_645),
.Y(n_5689)
);

NAND2xp5_ASAP7_75t_L g5690 ( 
.A(n_5451),
.B(n_647),
.Y(n_5690)
);

BUFx8_ASAP7_75t_L g5691 ( 
.A(n_5489),
.Y(n_5691)
);

OAI21x1_ASAP7_75t_L g5692 ( 
.A1(n_5393),
.A2(n_648),
.B(n_647),
.Y(n_5692)
);

AND2x4_ASAP7_75t_L g5693 ( 
.A(n_5421),
.B(n_5493),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_5494),
.Y(n_5694)
);

O2A1O1Ixp33_ASAP7_75t_SL g5695 ( 
.A1(n_5565),
.A2(n_648),
.B(n_649),
.C(n_647),
.Y(n_5695)
);

A2O1A1Ixp33_ASAP7_75t_L g5696 ( 
.A1(n_5397),
.A2(n_650),
.B(n_651),
.C(n_649),
.Y(n_5696)
);

AND2x4_ASAP7_75t_L g5697 ( 
.A(n_5421),
.B(n_649),
.Y(n_5697)
);

AOI21xp5_ASAP7_75t_L g5698 ( 
.A1(n_5554),
.A2(n_651),
.B(n_650),
.Y(n_5698)
);

NAND2xp5_ASAP7_75t_L g5699 ( 
.A(n_5390),
.B(n_651),
.Y(n_5699)
);

NOR2xp33_ASAP7_75t_L g5700 ( 
.A(n_5417),
.B(n_652),
.Y(n_5700)
);

INVx3_ASAP7_75t_L g5701 ( 
.A(n_5477),
.Y(n_5701)
);

OAI22xp33_ASAP7_75t_L g5702 ( 
.A1(n_5485),
.A2(n_653),
.B1(n_654),
.B2(n_652),
.Y(n_5702)
);

INVx1_ASAP7_75t_SL g5703 ( 
.A(n_5432),
.Y(n_5703)
);

AOI21xp5_ASAP7_75t_L g5704 ( 
.A1(n_5412),
.A2(n_653),
.B(n_652),
.Y(n_5704)
);

OAI21xp5_ASAP7_75t_L g5705 ( 
.A1(n_5499),
.A2(n_5500),
.B(n_5568),
.Y(n_5705)
);

INVx2_ASAP7_75t_L g5706 ( 
.A(n_5570),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5401),
.Y(n_5707)
);

AOI22xp33_ASAP7_75t_L g5708 ( 
.A1(n_5423),
.A2(n_5436),
.B1(n_5538),
.B2(n_5502),
.Y(n_5708)
);

INVx2_ASAP7_75t_L g5709 ( 
.A(n_5452),
.Y(n_5709)
);

BUFx2_ASAP7_75t_L g5710 ( 
.A(n_5490),
.Y(n_5710)
);

NAND2xp5_ASAP7_75t_L g5711 ( 
.A(n_5405),
.B(n_654),
.Y(n_5711)
);

AOI22xp33_ASAP7_75t_L g5712 ( 
.A1(n_5538),
.A2(n_655),
.B1(n_656),
.B2(n_654),
.Y(n_5712)
);

AO31x2_ASAP7_75t_L g5713 ( 
.A1(n_5442),
.A2(n_656),
.A3(n_657),
.B(n_655),
.Y(n_5713)
);

OAI21xp5_ASAP7_75t_L g5714 ( 
.A1(n_5523),
.A2(n_5527),
.B(n_5582),
.Y(n_5714)
);

NAND2xp5_ASAP7_75t_L g5715 ( 
.A(n_5447),
.B(n_655),
.Y(n_5715)
);

AOI221x1_ASAP7_75t_L g5716 ( 
.A1(n_5467),
.A2(n_659),
.B1(n_660),
.B2(n_658),
.C(n_657),
.Y(n_5716)
);

O2A1O1Ixp33_ASAP7_75t_SL g5717 ( 
.A1(n_5528),
.A2(n_658),
.B(n_659),
.C(n_657),
.Y(n_5717)
);

NAND2xp5_ASAP7_75t_L g5718 ( 
.A(n_5504),
.B(n_658),
.Y(n_5718)
);

AOI22xp5_ASAP7_75t_L g5719 ( 
.A1(n_5530),
.A2(n_660),
.B1(n_661),
.B2(n_659),
.Y(n_5719)
);

A2O1A1Ixp33_ASAP7_75t_L g5720 ( 
.A1(n_5438),
.A2(n_662),
.B(n_663),
.C(n_661),
.Y(n_5720)
);

O2A1O1Ixp33_ASAP7_75t_L g5721 ( 
.A1(n_5503),
.A2(n_663),
.B(n_664),
.C(n_662),
.Y(n_5721)
);

OR2x2_ASAP7_75t_L g5722 ( 
.A(n_5404),
.B(n_662),
.Y(n_5722)
);

O2A1O1Ixp33_ASAP7_75t_L g5723 ( 
.A1(n_5557),
.A2(n_664),
.B(n_665),
.C(n_663),
.Y(n_5723)
);

INVx2_ASAP7_75t_L g5724 ( 
.A(n_5421),
.Y(n_5724)
);

AOI21xp5_ASAP7_75t_L g5725 ( 
.A1(n_5456),
.A2(n_665),
.B(n_664),
.Y(n_5725)
);

INVx2_ASAP7_75t_SL g5726 ( 
.A(n_5496),
.Y(n_5726)
);

AOI21xp5_ASAP7_75t_L g5727 ( 
.A1(n_5484),
.A2(n_667),
.B(n_666),
.Y(n_5727)
);

AOI22xp5_ASAP7_75t_L g5728 ( 
.A1(n_5508),
.A2(n_667),
.B1(n_668),
.B2(n_666),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_5454),
.Y(n_5729)
);

INVx2_ASAP7_75t_L g5730 ( 
.A(n_5627),
.Y(n_5730)
);

NAND2xp5_ASAP7_75t_L g5731 ( 
.A(n_5605),
.B(n_5590),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5619),
.Y(n_5732)
);

OR2x2_ASAP7_75t_L g5733 ( 
.A(n_5709),
.B(n_5511),
.Y(n_5733)
);

OAI21x1_ASAP7_75t_L g5734 ( 
.A1(n_5667),
.A2(n_5482),
.B(n_5459),
.Y(n_5734)
);

INVx4_ASAP7_75t_L g5735 ( 
.A(n_5602),
.Y(n_5735)
);

NAND2xp5_ASAP7_75t_L g5736 ( 
.A(n_5607),
.B(n_5543),
.Y(n_5736)
);

INVx3_ASAP7_75t_L g5737 ( 
.A(n_5654),
.Y(n_5737)
);

NAND3xp33_ASAP7_75t_SL g5738 ( 
.A(n_5618),
.B(n_5560),
.C(n_5563),
.Y(n_5738)
);

NAND2xp5_ASAP7_75t_L g5739 ( 
.A(n_5606),
.B(n_5543),
.Y(n_5739)
);

NOR2xp67_ASAP7_75t_L g5740 ( 
.A(n_5621),
.B(n_5561),
.Y(n_5740)
);

OA21x2_ASAP7_75t_L g5741 ( 
.A1(n_5659),
.A2(n_5455),
.B(n_5458),
.Y(n_5741)
);

AOI21x1_ASAP7_75t_L g5742 ( 
.A1(n_5644),
.A2(n_5542),
.B(n_5480),
.Y(n_5742)
);

AOI21xp5_ASAP7_75t_L g5743 ( 
.A1(n_5628),
.A2(n_5480),
.B(n_5579),
.Y(n_5743)
);

OAI21xp5_ASAP7_75t_L g5744 ( 
.A1(n_5616),
.A2(n_5534),
.B(n_5537),
.Y(n_5744)
);

INVx1_ASAP7_75t_L g5745 ( 
.A(n_5611),
.Y(n_5745)
);

NOR2x1_ASAP7_75t_R g5746 ( 
.A(n_5639),
.B(n_5564),
.Y(n_5746)
);

OAI21x1_ASAP7_75t_L g5747 ( 
.A1(n_5592),
.A2(n_5473),
.B(n_5472),
.Y(n_5747)
);

INVx1_ASAP7_75t_SL g5748 ( 
.A(n_5610),
.Y(n_5748)
);

OAI21x1_ASAP7_75t_L g5749 ( 
.A1(n_5724),
.A2(n_5599),
.B(n_5596),
.Y(n_5749)
);

OAI21xp5_ASAP7_75t_L g5750 ( 
.A1(n_5646),
.A2(n_5540),
.B(n_5585),
.Y(n_5750)
);

INVx3_ASAP7_75t_L g5751 ( 
.A(n_5654),
.Y(n_5751)
);

OA21x2_ASAP7_75t_L g5752 ( 
.A1(n_5708),
.A2(n_5410),
.B(n_5535),
.Y(n_5752)
);

NOR2x1_ASAP7_75t_SL g5753 ( 
.A(n_5597),
.B(n_5497),
.Y(n_5753)
);

CKINVDCx5p33_ASAP7_75t_R g5754 ( 
.A(n_5593),
.Y(n_5754)
);

OAI21x1_ASAP7_75t_SL g5755 ( 
.A1(n_5614),
.A2(n_5478),
.B(n_5476),
.Y(n_5755)
);

OAI21x1_ASAP7_75t_L g5756 ( 
.A1(n_5603),
.A2(n_5492),
.B(n_5487),
.Y(n_5756)
);

AOI22xp33_ASAP7_75t_L g5757 ( 
.A1(n_5587),
.A2(n_5552),
.B1(n_5519),
.B2(n_5524),
.Y(n_5757)
);

AO21x2_ASAP7_75t_L g5758 ( 
.A1(n_5705),
.A2(n_5725),
.B(n_5714),
.Y(n_5758)
);

AND2x2_ASAP7_75t_L g5759 ( 
.A(n_5598),
.B(n_5493),
.Y(n_5759)
);

OAI21xp33_ASAP7_75t_SL g5760 ( 
.A1(n_5677),
.A2(n_5493),
.B(n_5584),
.Y(n_5760)
);

NOR2xp33_ASAP7_75t_SL g5761 ( 
.A(n_5633),
.B(n_5543),
.Y(n_5761)
);

OAI21x1_ASAP7_75t_L g5762 ( 
.A1(n_5624),
.A2(n_5569),
.B(n_668),
.Y(n_5762)
);

OAI21x1_ASAP7_75t_SL g5763 ( 
.A1(n_5601),
.A2(n_669),
.B(n_666),
.Y(n_5763)
);

OAI21x1_ASAP7_75t_L g5764 ( 
.A1(n_5701),
.A2(n_670),
.B(n_669),
.Y(n_5764)
);

INVx2_ASAP7_75t_L g5765 ( 
.A(n_5615),
.Y(n_5765)
);

OAI21x1_ASAP7_75t_L g5766 ( 
.A1(n_5653),
.A2(n_671),
.B(n_670),
.Y(n_5766)
);

INVx3_ASAP7_75t_L g5767 ( 
.A(n_5691),
.Y(n_5767)
);

OAI21x1_ASAP7_75t_L g5768 ( 
.A1(n_5588),
.A2(n_5631),
.B(n_5594),
.Y(n_5768)
);

INVx1_ASAP7_75t_L g5769 ( 
.A(n_5626),
.Y(n_5769)
);

INVx2_ASAP7_75t_L g5770 ( 
.A(n_5647),
.Y(n_5770)
);

NAND2x1p5_ASAP7_75t_L g5771 ( 
.A(n_5703),
.B(n_675),
.Y(n_5771)
);

OAI21x1_ASAP7_75t_L g5772 ( 
.A1(n_5686),
.A2(n_671),
.B(n_670),
.Y(n_5772)
);

OAI21x1_ASAP7_75t_L g5773 ( 
.A1(n_5698),
.A2(n_672),
.B(n_671),
.Y(n_5773)
);

NOR2xp33_ASAP7_75t_L g5774 ( 
.A(n_5668),
.B(n_5666),
.Y(n_5774)
);

CKINVDCx5p33_ASAP7_75t_R g5775 ( 
.A(n_5609),
.Y(n_5775)
);

AO21x1_ASAP7_75t_L g5776 ( 
.A1(n_5697),
.A2(n_12),
.B(n_13),
.Y(n_5776)
);

INVx2_ASAP7_75t_L g5777 ( 
.A(n_5647),
.Y(n_5777)
);

OAI21x1_ASAP7_75t_L g5778 ( 
.A1(n_5689),
.A2(n_5656),
.B(n_5663),
.Y(n_5778)
);

OAI21x1_ASAP7_75t_SL g5779 ( 
.A1(n_5726),
.A2(n_673),
.B(n_672),
.Y(n_5779)
);

AO21x2_ASAP7_75t_L g5780 ( 
.A1(n_5693),
.A2(n_674),
.B(n_672),
.Y(n_5780)
);

AND2x4_ASAP7_75t_L g5781 ( 
.A(n_5710),
.B(n_674),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5665),
.Y(n_5782)
);

OR2x2_ASAP7_75t_L g5783 ( 
.A(n_5625),
.B(n_674),
.Y(n_5783)
);

OR2x2_ASAP7_75t_L g5784 ( 
.A(n_5649),
.B(n_675),
.Y(n_5784)
);

BUFx3_ASAP7_75t_L g5785 ( 
.A(n_5595),
.Y(n_5785)
);

AND2x4_ASAP7_75t_L g5786 ( 
.A(n_5729),
.B(n_675),
.Y(n_5786)
);

NAND2xp5_ASAP7_75t_L g5787 ( 
.A(n_5707),
.B(n_1056),
.Y(n_5787)
);

HB1xp67_ASAP7_75t_L g5788 ( 
.A(n_5641),
.Y(n_5788)
);

AOI21xp5_ASAP7_75t_L g5789 ( 
.A1(n_5629),
.A2(n_677),
.B(n_676),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_5671),
.Y(n_5790)
);

AND2x4_ASAP7_75t_L g5791 ( 
.A(n_5660),
.B(n_677),
.Y(n_5791)
);

OAI21x1_ASAP7_75t_L g5792 ( 
.A1(n_5678),
.A2(n_678),
.B(n_677),
.Y(n_5792)
);

OR2x2_ASAP7_75t_L g5793 ( 
.A(n_5630),
.B(n_678),
.Y(n_5793)
);

OAI21x1_ASAP7_75t_L g5794 ( 
.A1(n_5655),
.A2(n_5679),
.B(n_5658),
.Y(n_5794)
);

OAI22xp5_ASAP7_75t_L g5795 ( 
.A1(n_5638),
.A2(n_679),
.B1(n_680),
.B2(n_678),
.Y(n_5795)
);

OAI22xp5_ASAP7_75t_L g5796 ( 
.A1(n_5635),
.A2(n_680),
.B1(n_681),
.B2(n_679),
.Y(n_5796)
);

OR2x2_ASAP7_75t_L g5797 ( 
.A(n_5706),
.B(n_681),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5673),
.Y(n_5798)
);

AND2x2_ASAP7_75t_L g5799 ( 
.A(n_5688),
.B(n_681),
.Y(n_5799)
);

INVx2_ASAP7_75t_L g5800 ( 
.A(n_5694),
.Y(n_5800)
);

OAI21x1_ASAP7_75t_L g5801 ( 
.A1(n_5670),
.A2(n_683),
.B(n_682),
.Y(n_5801)
);

INVx3_ASAP7_75t_L g5802 ( 
.A(n_5660),
.Y(n_5802)
);

OA21x2_ASAP7_75t_L g5803 ( 
.A1(n_5687),
.A2(n_13),
.B(n_14),
.Y(n_5803)
);

INVx1_ASAP7_75t_L g5804 ( 
.A(n_5608),
.Y(n_5804)
);

OAI21x1_ASAP7_75t_L g5805 ( 
.A1(n_5692),
.A2(n_684),
.B(n_683),
.Y(n_5805)
);

NOR2xp33_ASAP7_75t_L g5806 ( 
.A(n_5620),
.B(n_14),
.Y(n_5806)
);

INVx1_ASAP7_75t_SL g5807 ( 
.A(n_5685),
.Y(n_5807)
);

A2O1A1Ixp33_ASAP7_75t_L g5808 ( 
.A1(n_5664),
.A2(n_685),
.B(n_686),
.C(n_683),
.Y(n_5808)
);

OAI21x1_ASAP7_75t_L g5809 ( 
.A1(n_5669),
.A2(n_686),
.B(n_685),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_5637),
.Y(n_5810)
);

NAND2xp5_ASAP7_75t_L g5811 ( 
.A(n_5637),
.B(n_1050),
.Y(n_5811)
);

OA21x2_ASAP7_75t_L g5812 ( 
.A1(n_5693),
.A2(n_14),
.B(n_15),
.Y(n_5812)
);

AO21x2_ASAP7_75t_L g5813 ( 
.A1(n_5697),
.A2(n_687),
.B(n_685),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5637),
.Y(n_5814)
);

OAI21x1_ASAP7_75t_L g5815 ( 
.A1(n_5640),
.A2(n_688),
.B(n_687),
.Y(n_5815)
);

OA21x2_ASAP7_75t_L g5816 ( 
.A1(n_5652),
.A2(n_14),
.B(n_16),
.Y(n_5816)
);

AOI21xp5_ASAP7_75t_L g5817 ( 
.A1(n_5657),
.A2(n_688),
.B(n_687),
.Y(n_5817)
);

CKINVDCx20_ASAP7_75t_R g5818 ( 
.A(n_5676),
.Y(n_5818)
);

OAI21x1_ASAP7_75t_SL g5819 ( 
.A1(n_5617),
.A2(n_5600),
.B(n_5612),
.Y(n_5819)
);

OAI21x1_ASAP7_75t_SL g5820 ( 
.A1(n_5642),
.A2(n_690),
.B(n_689),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5715),
.Y(n_5821)
);

OAI21x1_ASAP7_75t_L g5822 ( 
.A1(n_5643),
.A2(n_690),
.B(n_689),
.Y(n_5822)
);

OAI21x1_ASAP7_75t_L g5823 ( 
.A1(n_5651),
.A2(n_691),
.B(n_689),
.Y(n_5823)
);

NOR2xp67_ASAP7_75t_L g5824 ( 
.A(n_5683),
.B(n_691),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5722),
.Y(n_5825)
);

AO31x2_ASAP7_75t_L g5826 ( 
.A1(n_5589),
.A2(n_692),
.A3(n_693),
.B(n_691),
.Y(n_5826)
);

OAI21x1_ASAP7_75t_L g5827 ( 
.A1(n_5727),
.A2(n_693),
.B(n_692),
.Y(n_5827)
);

NOR2x1_ASAP7_75t_L g5828 ( 
.A(n_5680),
.B(n_16),
.Y(n_5828)
);

OA21x2_ASAP7_75t_L g5829 ( 
.A1(n_5650),
.A2(n_16),
.B(n_17),
.Y(n_5829)
);

INVx8_ASAP7_75t_L g5830 ( 
.A(n_5660),
.Y(n_5830)
);

OAI21x1_ASAP7_75t_L g5831 ( 
.A1(n_5645),
.A2(n_693),
.B(n_692),
.Y(n_5831)
);

HB1xp67_ASAP7_75t_L g5832 ( 
.A(n_5713),
.Y(n_5832)
);

INVx6_ASAP7_75t_L g5833 ( 
.A(n_5636),
.Y(n_5833)
);

AOI21xp5_ASAP7_75t_L g5834 ( 
.A1(n_5720),
.A2(n_695),
.B(n_694),
.Y(n_5834)
);

OAI21x1_ASAP7_75t_L g5835 ( 
.A1(n_5623),
.A2(n_695),
.B(n_694),
.Y(n_5835)
);

AO21x2_ASAP7_75t_L g5836 ( 
.A1(n_5632),
.A2(n_697),
.B(n_696),
.Y(n_5836)
);

AOI21xp5_ASAP7_75t_L g5837 ( 
.A1(n_5717),
.A2(n_698),
.B(n_696),
.Y(n_5837)
);

AO21x2_ASAP7_75t_L g5838 ( 
.A1(n_5702),
.A2(n_698),
.B(n_696),
.Y(n_5838)
);

AOI22xp33_ASAP7_75t_L g5839 ( 
.A1(n_5634),
.A2(n_700),
.B1(n_701),
.B2(n_699),
.Y(n_5839)
);

INVx3_ASAP7_75t_L g5840 ( 
.A(n_5713),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5699),
.Y(n_5841)
);

OAI21x1_ASAP7_75t_SL g5842 ( 
.A1(n_5622),
.A2(n_701),
.B(n_699),
.Y(n_5842)
);

AO21x2_ASAP7_75t_L g5843 ( 
.A1(n_5690),
.A2(n_5674),
.B(n_5684),
.Y(n_5843)
);

BUFx2_ASAP7_75t_L g5844 ( 
.A(n_5713),
.Y(n_5844)
);

AND2x2_ASAP7_75t_SL g5845 ( 
.A(n_5712),
.B(n_699),
.Y(n_5845)
);

AOI21xp5_ASAP7_75t_L g5846 ( 
.A1(n_5695),
.A2(n_702),
.B(n_701),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_5711),
.Y(n_5847)
);

OR2x2_ASAP7_75t_L g5848 ( 
.A(n_5718),
.B(n_702),
.Y(n_5848)
);

AND2x2_ASAP7_75t_L g5849 ( 
.A(n_5700),
.B(n_703),
.Y(n_5849)
);

OAI21x1_ASAP7_75t_SL g5850 ( 
.A1(n_5704),
.A2(n_5682),
.B(n_5721),
.Y(n_5850)
);

OAI21x1_ASAP7_75t_L g5851 ( 
.A1(n_5662),
.A2(n_704),
.B(n_703),
.Y(n_5851)
);

NOR2xp33_ASAP7_75t_L g5852 ( 
.A(n_5604),
.B(n_16),
.Y(n_5852)
);

OR2x6_ASAP7_75t_L g5853 ( 
.A(n_5681),
.B(n_705),
.Y(n_5853)
);

INVxp33_ASAP7_75t_L g5854 ( 
.A(n_5719),
.Y(n_5854)
);

INVx3_ASAP7_75t_L g5855 ( 
.A(n_5591),
.Y(n_5855)
);

OAI21xp5_ASAP7_75t_L g5856 ( 
.A1(n_5696),
.A2(n_17),
.B(n_18),
.Y(n_5856)
);

BUFx6f_ASAP7_75t_L g5857 ( 
.A(n_5723),
.Y(n_5857)
);

INVx5_ASAP7_75t_L g5858 ( 
.A(n_5716),
.Y(n_5858)
);

INVx2_ASAP7_75t_SL g5859 ( 
.A(n_5728),
.Y(n_5859)
);

OAI21x1_ASAP7_75t_L g5860 ( 
.A1(n_5675),
.A2(n_706),
.B(n_705),
.Y(n_5860)
);

OA21x2_ASAP7_75t_L g5861 ( 
.A1(n_5661),
.A2(n_17),
.B(n_18),
.Y(n_5861)
);

INVx1_ASAP7_75t_L g5862 ( 
.A(n_5672),
.Y(n_5862)
);

AOI22xp33_ASAP7_75t_L g5863 ( 
.A1(n_5862),
.A2(n_5613),
.B1(n_5648),
.B2(n_706),
.Y(n_5863)
);

OR2x2_ASAP7_75t_L g5864 ( 
.A(n_5731),
.B(n_18),
.Y(n_5864)
);

NAND2xp5_ASAP7_75t_L g5865 ( 
.A(n_5844),
.B(n_705),
.Y(n_5865)
);

NAND2xp5_ASAP7_75t_L g5866 ( 
.A(n_5844),
.B(n_707),
.Y(n_5866)
);

AOI21xp5_ASAP7_75t_L g5867 ( 
.A1(n_5753),
.A2(n_18),
.B(n_19),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5800),
.Y(n_5868)
);

AOI21xp5_ASAP7_75t_L g5869 ( 
.A1(n_5789),
.A2(n_19),
.B(n_20),
.Y(n_5869)
);

NAND2xp5_ASAP7_75t_L g5870 ( 
.A(n_5832),
.B(n_707),
.Y(n_5870)
);

AND2x2_ASAP7_75t_L g5871 ( 
.A(n_5759),
.B(n_19),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_5732),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_5739),
.Y(n_5873)
);

INVx2_ASAP7_75t_L g5874 ( 
.A(n_5788),
.Y(n_5874)
);

OAI22xp5_ASAP7_75t_L g5875 ( 
.A1(n_5833),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_5875)
);

OR2x2_ASAP7_75t_L g5876 ( 
.A(n_5730),
.B(n_20),
.Y(n_5876)
);

INVx2_ASAP7_75t_L g5877 ( 
.A(n_5794),
.Y(n_5877)
);

AND2x4_ASAP7_75t_L g5878 ( 
.A(n_5737),
.B(n_1046),
.Y(n_5878)
);

NAND2xp5_ASAP7_75t_L g5879 ( 
.A(n_5736),
.B(n_707),
.Y(n_5879)
);

A2O1A1Ixp33_ASAP7_75t_L g5880 ( 
.A1(n_5740),
.A2(n_709),
.B(n_710),
.C(n_708),
.Y(n_5880)
);

OR2x2_ASAP7_75t_L g5881 ( 
.A(n_5733),
.B(n_21),
.Y(n_5881)
);

AOI21xp5_ASAP7_75t_L g5882 ( 
.A1(n_5743),
.A2(n_21),
.B(n_22),
.Y(n_5882)
);

AOI21xp5_ASAP7_75t_SL g5883 ( 
.A1(n_5812),
.A2(n_22),
.B(n_23),
.Y(n_5883)
);

OA21x2_ASAP7_75t_L g5884 ( 
.A1(n_5768),
.A2(n_22),
.B(n_23),
.Y(n_5884)
);

AO31x2_ASAP7_75t_L g5885 ( 
.A1(n_5810),
.A2(n_25),
.A3(n_22),
.B(n_24),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5745),
.Y(n_5886)
);

BUFx6f_ASAP7_75t_L g5887 ( 
.A(n_5767),
.Y(n_5887)
);

INVx3_ASAP7_75t_L g5888 ( 
.A(n_5735),
.Y(n_5888)
);

OA21x2_ASAP7_75t_L g5889 ( 
.A1(n_5755),
.A2(n_24),
.B(n_25),
.Y(n_5889)
);

CKINVDCx6p67_ASAP7_75t_R g5890 ( 
.A(n_5748),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5769),
.Y(n_5891)
);

AND2x2_ASAP7_75t_L g5892 ( 
.A(n_5770),
.B(n_24),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5782),
.Y(n_5893)
);

AO21x2_ASAP7_75t_L g5894 ( 
.A1(n_5819),
.A2(n_710),
.B(n_708),
.Y(n_5894)
);

NOR2xp67_ASAP7_75t_L g5895 ( 
.A(n_5855),
.B(n_26),
.Y(n_5895)
);

OR2x2_ASAP7_75t_L g5896 ( 
.A(n_5804),
.B(n_26),
.Y(n_5896)
);

AOI21xp5_ASAP7_75t_L g5897 ( 
.A1(n_5812),
.A2(n_27),
.B(n_28),
.Y(n_5897)
);

BUFx3_ASAP7_75t_L g5898 ( 
.A(n_5754),
.Y(n_5898)
);

A2O1A1Ixp33_ASAP7_75t_L g5899 ( 
.A1(n_5778),
.A2(n_710),
.B(n_711),
.C(n_708),
.Y(n_5899)
);

AOI22xp33_ASAP7_75t_L g5900 ( 
.A1(n_5857),
.A2(n_712),
.B1(n_713),
.B2(n_711),
.Y(n_5900)
);

OR2x6_ASAP7_75t_L g5901 ( 
.A(n_5771),
.B(n_711),
.Y(n_5901)
);

NAND2xp5_ASAP7_75t_L g5902 ( 
.A(n_5814),
.B(n_712),
.Y(n_5902)
);

BUFx3_ASAP7_75t_L g5903 ( 
.A(n_5775),
.Y(n_5903)
);

A2O1A1Ixp33_ASAP7_75t_L g5904 ( 
.A1(n_5828),
.A2(n_713),
.B(n_714),
.C(n_712),
.Y(n_5904)
);

INVx2_ASAP7_75t_L g5905 ( 
.A(n_5756),
.Y(n_5905)
);

BUFx10_ASAP7_75t_L g5906 ( 
.A(n_5781),
.Y(n_5906)
);

CKINVDCx5p33_ASAP7_75t_R g5907 ( 
.A(n_5751),
.Y(n_5907)
);

OAI21xp5_ASAP7_75t_L g5908 ( 
.A1(n_5817),
.A2(n_27),
.B(n_28),
.Y(n_5908)
);

AOI21xp5_ASAP7_75t_L g5909 ( 
.A1(n_5746),
.A2(n_27),
.B(n_28),
.Y(n_5909)
);

OA21x2_ASAP7_75t_L g5910 ( 
.A1(n_5757),
.A2(n_5744),
.B(n_5747),
.Y(n_5910)
);

AO21x1_ASAP7_75t_L g5911 ( 
.A1(n_5761),
.A2(n_28),
.B(n_29),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5790),
.Y(n_5912)
);

INVx4_ASAP7_75t_L g5913 ( 
.A(n_5830),
.Y(n_5913)
);

AOI21xp5_ASAP7_75t_L g5914 ( 
.A1(n_5750),
.A2(n_29),
.B(n_30),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_5749),
.Y(n_5915)
);

AO21x2_ASAP7_75t_L g5916 ( 
.A1(n_5811),
.A2(n_715),
.B(n_714),
.Y(n_5916)
);

OR2x6_ASAP7_75t_L g5917 ( 
.A(n_5833),
.B(n_5779),
.Y(n_5917)
);

OR2x2_ASAP7_75t_L g5918 ( 
.A(n_5765),
.B(n_29),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_5798),
.Y(n_5919)
);

INVx2_ASAP7_75t_L g5920 ( 
.A(n_5742),
.Y(n_5920)
);

AOI21xp5_ASAP7_75t_L g5921 ( 
.A1(n_5780),
.A2(n_30),
.B(n_31),
.Y(n_5921)
);

BUFx2_ASAP7_75t_L g5922 ( 
.A(n_5785),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_5847),
.Y(n_5923)
);

OAI21xp33_ASAP7_75t_L g5924 ( 
.A1(n_5854),
.A2(n_5852),
.B(n_5760),
.Y(n_5924)
);

AO31x2_ASAP7_75t_L g5925 ( 
.A1(n_5774),
.A2(n_32),
.A3(n_30),
.B(n_31),
.Y(n_5925)
);

AO31x2_ASAP7_75t_L g5926 ( 
.A1(n_5776),
.A2(n_33),
.A3(n_31),
.B(n_32),
.Y(n_5926)
);

A2O1A1Ixp33_ASAP7_75t_L g5927 ( 
.A1(n_5807),
.A2(n_716),
.B(n_717),
.C(n_715),
.Y(n_5927)
);

OAI21x1_ASAP7_75t_L g5928 ( 
.A1(n_5734),
.A2(n_716),
.B(n_715),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_5841),
.Y(n_5929)
);

OA21x2_ASAP7_75t_L g5930 ( 
.A1(n_5801),
.A2(n_31),
.B(n_32),
.Y(n_5930)
);

AOI21x1_ASAP7_75t_L g5931 ( 
.A1(n_5816),
.A2(n_32),
.B(n_33),
.Y(n_5931)
);

INVx1_ASAP7_75t_L g5932 ( 
.A(n_5825),
.Y(n_5932)
);

INVx2_ASAP7_75t_L g5933 ( 
.A(n_5840),
.Y(n_5933)
);

AND2x4_ASAP7_75t_L g5934 ( 
.A(n_5777),
.B(n_5791),
.Y(n_5934)
);

OAI21x1_ASAP7_75t_L g5935 ( 
.A1(n_5752),
.A2(n_717),
.B(n_716),
.Y(n_5935)
);

OA21x2_ASAP7_75t_L g5936 ( 
.A1(n_5821),
.A2(n_34),
.B(n_35),
.Y(n_5936)
);

NOR2xp33_ASAP7_75t_L g5937 ( 
.A(n_5857),
.B(n_34),
.Y(n_5937)
);

NAND2xp5_ASAP7_75t_L g5938 ( 
.A(n_5752),
.B(n_718),
.Y(n_5938)
);

NOR2x1_ASAP7_75t_R g5939 ( 
.A(n_5858),
.B(n_34),
.Y(n_5939)
);

AOI221xp5_ASAP7_75t_L g5940 ( 
.A1(n_5839),
.A2(n_720),
.B1(n_721),
.B2(n_719),
.C(n_718),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5797),
.Y(n_5941)
);

INVx2_ASAP7_75t_L g5942 ( 
.A(n_5813),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5787),
.Y(n_5943)
);

INVx1_ASAP7_75t_L g5944 ( 
.A(n_5799),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5784),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5802),
.B(n_34),
.Y(n_5946)
);

OR2x2_ASAP7_75t_L g5947 ( 
.A(n_5783),
.B(n_35),
.Y(n_5947)
);

NAND2xp5_ASAP7_75t_SL g5948 ( 
.A(n_5818),
.B(n_35),
.Y(n_5948)
);

OAI221xp5_ASAP7_75t_L g5949 ( 
.A1(n_5808),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.C(n_38),
.Y(n_5949)
);

OAI21x1_ASAP7_75t_L g5950 ( 
.A1(n_5741),
.A2(n_5792),
.B(n_5815),
.Y(n_5950)
);

NAND2xp5_ASAP7_75t_L g5951 ( 
.A(n_5758),
.B(n_719),
.Y(n_5951)
);

OR2x6_ASAP7_75t_L g5952 ( 
.A(n_5830),
.B(n_719),
.Y(n_5952)
);

AOI21xp5_ASAP7_75t_L g5953 ( 
.A1(n_5816),
.A2(n_5861),
.B(n_5803),
.Y(n_5953)
);

BUFx10_ASAP7_75t_L g5954 ( 
.A(n_5786),
.Y(n_5954)
);

AOI21xp5_ASAP7_75t_L g5955 ( 
.A1(n_5861),
.A2(n_36),
.B(n_37),
.Y(n_5955)
);

AND2x2_ASAP7_75t_L g5956 ( 
.A(n_5741),
.B(n_36),
.Y(n_5956)
);

NAND2xp5_ASAP7_75t_L g5957 ( 
.A(n_5803),
.B(n_720),
.Y(n_5957)
);

AO31x2_ASAP7_75t_L g5958 ( 
.A1(n_5806),
.A2(n_5796),
.A3(n_5795),
.B(n_5846),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5793),
.Y(n_5959)
);

A2O1A1Ixp33_ASAP7_75t_L g5960 ( 
.A1(n_5831),
.A2(n_721),
.B(n_722),
.C(n_720),
.Y(n_5960)
);

AND2x2_ASAP7_75t_L g5961 ( 
.A(n_5859),
.B(n_36),
.Y(n_5961)
);

NAND2x1p5_ASAP7_75t_L g5962 ( 
.A(n_5764),
.B(n_721),
.Y(n_5962)
);

AOI21x1_ASAP7_75t_L g5963 ( 
.A1(n_5829),
.A2(n_37),
.B(n_38),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5848),
.Y(n_5964)
);

OR2x2_ASAP7_75t_SL g5965 ( 
.A(n_5829),
.B(n_38),
.Y(n_5965)
);

OAI21x1_ASAP7_75t_L g5966 ( 
.A1(n_5809),
.A2(n_723),
.B(n_722),
.Y(n_5966)
);

AOI21xp5_ASAP7_75t_L g5967 ( 
.A1(n_5738),
.A2(n_38),
.B(n_39),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5843),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5835),
.Y(n_5969)
);

AOI22xp33_ASAP7_75t_L g5970 ( 
.A1(n_5853),
.A2(n_723),
.B1(n_724),
.B2(n_722),
.Y(n_5970)
);

NAND2xp5_ASAP7_75t_SL g5971 ( 
.A(n_5858),
.B(n_39),
.Y(n_5971)
);

A2O1A1Ixp33_ASAP7_75t_L g5972 ( 
.A1(n_5822),
.A2(n_724),
.B(n_725),
.C(n_723),
.Y(n_5972)
);

INVx1_ASAP7_75t_L g5973 ( 
.A(n_5851),
.Y(n_5973)
);

AOI21xp5_ASAP7_75t_L g5974 ( 
.A1(n_5820),
.A2(n_39),
.B(n_40),
.Y(n_5974)
);

AND2x4_ASAP7_75t_L g5975 ( 
.A(n_5853),
.B(n_1049),
.Y(n_5975)
);

OAI22xp33_ASAP7_75t_L g5976 ( 
.A1(n_5858),
.A2(n_1052),
.B1(n_1053),
.B2(n_1049),
.Y(n_5976)
);

A2O1A1Ixp33_ASAP7_75t_L g5977 ( 
.A1(n_5824),
.A2(n_5823),
.B(n_5856),
.C(n_5860),
.Y(n_5977)
);

AOI22xp33_ASAP7_75t_L g5978 ( 
.A1(n_5845),
.A2(n_725),
.B1(n_726),
.B2(n_724),
.Y(n_5978)
);

AND2x2_ASAP7_75t_L g5979 ( 
.A(n_5849),
.B(n_39),
.Y(n_5979)
);

AOI22xp33_ASAP7_75t_L g5980 ( 
.A1(n_5850),
.A2(n_726),
.B1(n_727),
.B2(n_725),
.Y(n_5980)
);

INVx1_ASAP7_75t_L g5981 ( 
.A(n_5762),
.Y(n_5981)
);

BUFx2_ASAP7_75t_L g5982 ( 
.A(n_5826),
.Y(n_5982)
);

INVx2_ASAP7_75t_L g5983 ( 
.A(n_5836),
.Y(n_5983)
);

INVx2_ASAP7_75t_L g5984 ( 
.A(n_5826),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5805),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5766),
.Y(n_5986)
);

AND2x2_ASAP7_75t_L g5987 ( 
.A(n_5922),
.B(n_5838),
.Y(n_5987)
);

OAI21xp5_ASAP7_75t_SL g5988 ( 
.A1(n_5867),
.A2(n_5837),
.B(n_5834),
.Y(n_5988)
);

INVx3_ASAP7_75t_L g5989 ( 
.A(n_5887),
.Y(n_5989)
);

AO21x2_ASAP7_75t_L g5990 ( 
.A1(n_5968),
.A2(n_5842),
.B(n_5763),
.Y(n_5990)
);

BUFx12f_ASAP7_75t_L g5991 ( 
.A(n_5887),
.Y(n_5991)
);

BUFx12f_ASAP7_75t_L g5992 ( 
.A(n_5907),
.Y(n_5992)
);

BUFx2_ASAP7_75t_L g5993 ( 
.A(n_5917),
.Y(n_5993)
);

INVx2_ASAP7_75t_SL g5994 ( 
.A(n_5888),
.Y(n_5994)
);

AO32x2_ASAP7_75t_L g5995 ( 
.A1(n_5875),
.A2(n_5773),
.A3(n_5772),
.B1(n_5827),
.B2(n_729),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5923),
.Y(n_5996)
);

CKINVDCx16_ASAP7_75t_R g5997 ( 
.A(n_5901),
.Y(n_5997)
);

BUFx2_ASAP7_75t_L g5998 ( 
.A(n_5917),
.Y(n_5998)
);

INVx1_ASAP7_75t_L g5999 ( 
.A(n_5929),
.Y(n_5999)
);

OAI21xp5_ASAP7_75t_SL g6000 ( 
.A1(n_5863),
.A2(n_40),
.B(n_41),
.Y(n_6000)
);

AOI22xp33_ASAP7_75t_L g6001 ( 
.A1(n_5924),
.A2(n_727),
.B1(n_729),
.B2(n_726),
.Y(n_6001)
);

AOI22xp33_ASAP7_75t_L g6002 ( 
.A1(n_5894),
.A2(n_730),
.B1(n_731),
.B2(n_729),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_5981),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5985),
.Y(n_6004)
);

OR2x2_ASAP7_75t_L g6005 ( 
.A(n_5873),
.B(n_40),
.Y(n_6005)
);

AND2x2_ASAP7_75t_L g6006 ( 
.A(n_5874),
.B(n_40),
.Y(n_6006)
);

HB1xp67_ASAP7_75t_L g6007 ( 
.A(n_5956),
.Y(n_6007)
);

NAND2xp5_ASAP7_75t_L g6008 ( 
.A(n_5973),
.B(n_41),
.Y(n_6008)
);

INVx2_ASAP7_75t_L g6009 ( 
.A(n_5868),
.Y(n_6009)
);

AND2x4_ASAP7_75t_L g6010 ( 
.A(n_5913),
.B(n_730),
.Y(n_6010)
);

AOI22xp33_ASAP7_75t_L g6011 ( 
.A1(n_5975),
.A2(n_732),
.B1(n_733),
.B2(n_731),
.Y(n_6011)
);

NOR2xp33_ASAP7_75t_R g6012 ( 
.A(n_5890),
.B(n_42),
.Y(n_6012)
);

AND2x2_ASAP7_75t_L g6013 ( 
.A(n_5871),
.B(n_42),
.Y(n_6013)
);

AND2x2_ASAP7_75t_L g6014 ( 
.A(n_5934),
.B(n_42),
.Y(n_6014)
);

CKINVDCx5p33_ASAP7_75t_R g6015 ( 
.A(n_5903),
.Y(n_6015)
);

CKINVDCx14_ASAP7_75t_R g6016 ( 
.A(n_5906),
.Y(n_6016)
);

AND2x2_ASAP7_75t_L g6017 ( 
.A(n_5959),
.B(n_42),
.Y(n_6017)
);

OAI21xp5_ASAP7_75t_SL g6018 ( 
.A1(n_5909),
.A2(n_43),
.B(n_44),
.Y(n_6018)
);

XOR2x2_ASAP7_75t_SL g6019 ( 
.A(n_5962),
.B(n_43),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_5872),
.Y(n_6020)
);

NAND2xp33_ASAP7_75t_R g6021 ( 
.A(n_5884),
.B(n_44),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_5886),
.Y(n_6022)
);

AND2x2_ASAP7_75t_L g6023 ( 
.A(n_5943),
.B(n_44),
.Y(n_6023)
);

AOI22xp5_ASAP7_75t_L g6024 ( 
.A1(n_5911),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_6024)
);

AOI22xp33_ASAP7_75t_SL g6025 ( 
.A1(n_5910),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_6025)
);

AND2x2_ASAP7_75t_L g6026 ( 
.A(n_5945),
.B(n_45),
.Y(n_6026)
);

HB1xp67_ASAP7_75t_L g6027 ( 
.A(n_5936),
.Y(n_6027)
);

CKINVDCx5p33_ASAP7_75t_R g6028 ( 
.A(n_5898),
.Y(n_6028)
);

INVx1_ASAP7_75t_L g6029 ( 
.A(n_5891),
.Y(n_6029)
);

AOI22xp33_ASAP7_75t_SL g6030 ( 
.A1(n_5982),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_6030)
);

AOI22xp33_ASAP7_75t_SL g6031 ( 
.A1(n_5920),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_6031)
);

AND2x4_ASAP7_75t_L g6032 ( 
.A(n_5952),
.B(n_731),
.Y(n_6032)
);

NOR2xp33_ASAP7_75t_L g6033 ( 
.A(n_5937),
.B(n_732),
.Y(n_6033)
);

INVx3_ASAP7_75t_L g6034 ( 
.A(n_5952),
.Y(n_6034)
);

CKINVDCx16_ASAP7_75t_R g6035 ( 
.A(n_5901),
.Y(n_6035)
);

AOI22xp33_ASAP7_75t_L g6036 ( 
.A1(n_5942),
.A2(n_733),
.B1(n_734),
.B2(n_732),
.Y(n_6036)
);

AND3x2_ASAP7_75t_L g6037 ( 
.A(n_5883),
.B(n_5908),
.C(n_5878),
.Y(n_6037)
);

OR2x2_ASAP7_75t_L g6038 ( 
.A(n_5879),
.B(n_47),
.Y(n_6038)
);

AO31x2_ASAP7_75t_L g6039 ( 
.A1(n_5983),
.A2(n_50),
.A3(n_48),
.B(n_49),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5893),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5912),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5919),
.Y(n_6042)
);

NAND2xp5_ASAP7_75t_L g6043 ( 
.A(n_5969),
.B(n_49),
.Y(n_6043)
);

CKINVDCx16_ASAP7_75t_R g6044 ( 
.A(n_5954),
.Y(n_6044)
);

INVx2_ASAP7_75t_L g6045 ( 
.A(n_5946),
.Y(n_6045)
);

CKINVDCx5p33_ASAP7_75t_R g6046 ( 
.A(n_5979),
.Y(n_6046)
);

AOI21xp5_ASAP7_75t_L g6047 ( 
.A1(n_5914),
.A2(n_49),
.B(n_50),
.Y(n_6047)
);

OR2x2_ASAP7_75t_L g6048 ( 
.A(n_5932),
.B(n_49),
.Y(n_6048)
);

INVx1_ASAP7_75t_L g6049 ( 
.A(n_5865),
.Y(n_6049)
);

OAI21xp5_ASAP7_75t_L g6050 ( 
.A1(n_5882),
.A2(n_50),
.B(n_51),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_5866),
.Y(n_6051)
);

OAI22xp5_ASAP7_75t_L g6052 ( 
.A1(n_5965),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_6052)
);

INVx1_ASAP7_75t_L g6053 ( 
.A(n_5986),
.Y(n_6053)
);

AND2x2_ASAP7_75t_L g6054 ( 
.A(n_5964),
.B(n_51),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5870),
.Y(n_6055)
);

CKINVDCx5p33_ASAP7_75t_R g6056 ( 
.A(n_5961),
.Y(n_6056)
);

INVx2_ASAP7_75t_L g6057 ( 
.A(n_5933),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5941),
.Y(n_6058)
);

INVx2_ASAP7_75t_L g6059 ( 
.A(n_5877),
.Y(n_6059)
);

AO31x2_ASAP7_75t_L g6060 ( 
.A1(n_5951),
.A2(n_5938),
.A3(n_5915),
.B(n_5984),
.Y(n_6060)
);

AOI22xp33_ASAP7_75t_SL g6061 ( 
.A1(n_5889),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_6061)
);

NOR2xp33_ASAP7_75t_R g6062 ( 
.A(n_5963),
.B(n_52),
.Y(n_6062)
);

INVx1_ASAP7_75t_L g6063 ( 
.A(n_5902),
.Y(n_6063)
);

AND2x2_ASAP7_75t_L g6064 ( 
.A(n_5944),
.B(n_53),
.Y(n_6064)
);

AOI22xp33_ASAP7_75t_L g6065 ( 
.A1(n_5895),
.A2(n_734),
.B1(n_735),
.B2(n_733),
.Y(n_6065)
);

INVx2_ASAP7_75t_L g6066 ( 
.A(n_5928),
.Y(n_6066)
);

OR2x6_ASAP7_75t_L g6067 ( 
.A(n_5967),
.B(n_735),
.Y(n_6067)
);

NOR2x1_ASAP7_75t_L g6068 ( 
.A(n_5971),
.B(n_53),
.Y(n_6068)
);

AND2x2_ASAP7_75t_L g6069 ( 
.A(n_5892),
.B(n_54),
.Y(n_6069)
);

INVx1_ASAP7_75t_L g6070 ( 
.A(n_5950),
.Y(n_6070)
);

NOR2xp33_ASAP7_75t_R g6071 ( 
.A(n_5931),
.B(n_54),
.Y(n_6071)
);

INVx1_ASAP7_75t_SL g6072 ( 
.A(n_5948),
.Y(n_6072)
);

BUFx2_ASAP7_75t_L g6073 ( 
.A(n_5939),
.Y(n_6073)
);

CKINVDCx16_ASAP7_75t_R g6074 ( 
.A(n_5947),
.Y(n_6074)
);

CKINVDCx16_ASAP7_75t_R g6075 ( 
.A(n_5881),
.Y(n_6075)
);

OAI22xp5_ASAP7_75t_L g6076 ( 
.A1(n_5953),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_6076)
);

O2A1O1Ixp33_ASAP7_75t_SL g6077 ( 
.A1(n_5977),
.A2(n_5904),
.B(n_5880),
.C(n_5899),
.Y(n_6077)
);

NOR2xp33_ASAP7_75t_L g6078 ( 
.A(n_5864),
.B(n_735),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_5876),
.Y(n_6079)
);

BUFx2_ASAP7_75t_L g6080 ( 
.A(n_5935),
.Y(n_6080)
);

NOR3xp33_ASAP7_75t_SL g6081 ( 
.A(n_5976),
.B(n_55),
.C(n_56),
.Y(n_6081)
);

AND2x2_ASAP7_75t_L g6082 ( 
.A(n_5918),
.B(n_55),
.Y(n_6082)
);

OAI22xp5_ASAP7_75t_L g6083 ( 
.A1(n_5897),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_6083)
);

AND2x2_ASAP7_75t_L g6084 ( 
.A(n_5905),
.B(n_56),
.Y(n_6084)
);

NAND2xp5_ASAP7_75t_L g6085 ( 
.A(n_5916),
.B(n_58),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5896),
.Y(n_6086)
);

XNOR2xp5_ASAP7_75t_L g6087 ( 
.A(n_5978),
.B(n_5980),
.Y(n_6087)
);

INVx1_ASAP7_75t_L g6088 ( 
.A(n_5885),
.Y(n_6088)
);

AND2x4_ASAP7_75t_L g6089 ( 
.A(n_5958),
.B(n_736),
.Y(n_6089)
);

INVxp67_ASAP7_75t_L g6090 ( 
.A(n_5957),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5885),
.Y(n_6091)
);

NOR2xp33_ASAP7_75t_R g6092 ( 
.A(n_5970),
.B(n_58),
.Y(n_6092)
);

NAND2xp5_ASAP7_75t_L g6093 ( 
.A(n_5925),
.B(n_5921),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_5925),
.Y(n_6094)
);

CKINVDCx5p33_ASAP7_75t_R g6095 ( 
.A(n_5900),
.Y(n_6095)
);

INVx2_ASAP7_75t_L g6096 ( 
.A(n_5926),
.Y(n_6096)
);

INVx1_ASAP7_75t_L g6097 ( 
.A(n_5926),
.Y(n_6097)
);

AOI22xp33_ASAP7_75t_SL g6098 ( 
.A1(n_5930),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_6098)
);

INVx2_ASAP7_75t_L g6099 ( 
.A(n_5966),
.Y(n_6099)
);

NAND3xp33_ASAP7_75t_L g6100 ( 
.A(n_5927),
.B(n_58),
.C(n_59),
.Y(n_6100)
);

NAND2xp33_ASAP7_75t_R g6101 ( 
.A(n_5869),
.B(n_59),
.Y(n_6101)
);

O2A1O1Ixp33_ASAP7_75t_L g6102 ( 
.A1(n_5960),
.A2(n_737),
.B(n_738),
.C(n_736),
.Y(n_6102)
);

OAI22xp5_ASAP7_75t_L g6103 ( 
.A1(n_5955),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_6103)
);

NAND2xp33_ASAP7_75t_R g6104 ( 
.A(n_5974),
.B(n_60),
.Y(n_6104)
);

NAND3xp33_ASAP7_75t_SL g6105 ( 
.A(n_5972),
.B(n_60),
.C(n_61),
.Y(n_6105)
);

NAND2xp33_ASAP7_75t_SL g6106 ( 
.A(n_5958),
.B(n_61),
.Y(n_6106)
);

BUFx4f_ASAP7_75t_SL g6107 ( 
.A(n_5940),
.Y(n_6107)
);

HB1xp67_ASAP7_75t_L g6108 ( 
.A(n_5949),
.Y(n_6108)
);

NOR2xp33_ASAP7_75t_L g6109 ( 
.A(n_5890),
.B(n_736),
.Y(n_6109)
);

BUFx2_ASAP7_75t_L g6110 ( 
.A(n_5922),
.Y(n_6110)
);

CKINVDCx16_ASAP7_75t_R g6111 ( 
.A(n_5901),
.Y(n_6111)
);

AND2x2_ASAP7_75t_L g6112 ( 
.A(n_5922),
.B(n_61),
.Y(n_6112)
);

INVx6_ASAP7_75t_L g6113 ( 
.A(n_5887),
.Y(n_6113)
);

NAND2xp5_ASAP7_75t_L g6114 ( 
.A(n_5956),
.B(n_62),
.Y(n_6114)
);

BUFx3_ASAP7_75t_L g6115 ( 
.A(n_5887),
.Y(n_6115)
);

AO31x2_ASAP7_75t_L g6116 ( 
.A1(n_5968),
.A2(n_65),
.A3(n_63),
.B(n_64),
.Y(n_6116)
);

INVx2_ASAP7_75t_SL g6117 ( 
.A(n_5887),
.Y(n_6117)
);

INVx1_ASAP7_75t_L g6118 ( 
.A(n_5923),
.Y(n_6118)
);

BUFx6f_ASAP7_75t_L g6119 ( 
.A(n_5887),
.Y(n_6119)
);

OAI22xp33_ASAP7_75t_L g6120 ( 
.A1(n_5917),
.A2(n_738),
.B1(n_739),
.B2(n_737),
.Y(n_6120)
);

AOI22xp5_ASAP7_75t_L g6121 ( 
.A1(n_5924),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_6121)
);

INVx2_ASAP7_75t_L g6122 ( 
.A(n_5922),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5923),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_5923),
.Y(n_6124)
);

NAND2xp5_ASAP7_75t_L g6125 ( 
.A(n_5956),
.B(n_63),
.Y(n_6125)
);

CKINVDCx11_ASAP7_75t_R g6126 ( 
.A(n_5890),
.Y(n_6126)
);

CKINVDCx16_ASAP7_75t_R g6127 ( 
.A(n_5901),
.Y(n_6127)
);

AO31x2_ASAP7_75t_L g6128 ( 
.A1(n_5968),
.A2(n_65),
.A3(n_63),
.B(n_64),
.Y(n_6128)
);

INVx2_ASAP7_75t_L g6129 ( 
.A(n_5922),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_5923),
.Y(n_6130)
);

CKINVDCx5p33_ASAP7_75t_R g6131 ( 
.A(n_5890),
.Y(n_6131)
);

NAND2xp5_ASAP7_75t_L g6132 ( 
.A(n_5956),
.B(n_65),
.Y(n_6132)
);

NAND2xp5_ASAP7_75t_L g6133 ( 
.A(n_5956),
.B(n_66),
.Y(n_6133)
);

INVx2_ASAP7_75t_L g6134 ( 
.A(n_5922),
.Y(n_6134)
);

NOR2xp33_ASAP7_75t_R g6135 ( 
.A(n_5890),
.B(n_66),
.Y(n_6135)
);

INVx2_ASAP7_75t_L g6136 ( 
.A(n_5922),
.Y(n_6136)
);

OAI21xp5_ASAP7_75t_L g6137 ( 
.A1(n_5867),
.A2(n_66),
.B(n_67),
.Y(n_6137)
);

INVx8_ASAP7_75t_L g6138 ( 
.A(n_5887),
.Y(n_6138)
);

AND2x4_ASAP7_75t_L g6139 ( 
.A(n_5888),
.B(n_737),
.Y(n_6139)
);

AND2x2_ASAP7_75t_L g6140 ( 
.A(n_5922),
.B(n_67),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_5923),
.Y(n_6141)
);

NOR2xp33_ASAP7_75t_R g6142 ( 
.A(n_5890),
.B(n_67),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5923),
.Y(n_6143)
);

OAI22xp5_ASAP7_75t_L g6144 ( 
.A1(n_5917),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_5923),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_5923),
.Y(n_6146)
);

OR2x2_ASAP7_75t_L g6147 ( 
.A(n_5873),
.B(n_68),
.Y(n_6147)
);

INVx1_ASAP7_75t_L g6148 ( 
.A(n_5923),
.Y(n_6148)
);

NAND2xp33_ASAP7_75t_R g6149 ( 
.A(n_5884),
.B(n_68),
.Y(n_6149)
);

OR2x2_ASAP7_75t_L g6150 ( 
.A(n_5873),
.B(n_69),
.Y(n_6150)
);

INVx1_ASAP7_75t_L g6151 ( 
.A(n_6110),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_6027),
.Y(n_6152)
);

INVx2_ASAP7_75t_L g6153 ( 
.A(n_6122),
.Y(n_6153)
);

OA21x2_ASAP7_75t_L g6154 ( 
.A1(n_6089),
.A2(n_69),
.B(n_70),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_6129),
.Y(n_6155)
);

INVx1_ASAP7_75t_L g6156 ( 
.A(n_6134),
.Y(n_6156)
);

OR2x6_ASAP7_75t_L g6157 ( 
.A(n_6138),
.B(n_738),
.Y(n_6157)
);

AND2x2_ASAP7_75t_L g6158 ( 
.A(n_5993),
.B(n_69),
.Y(n_6158)
);

OR2x6_ASAP7_75t_L g6159 ( 
.A(n_6138),
.B(n_739),
.Y(n_6159)
);

OR2x2_ASAP7_75t_L g6160 ( 
.A(n_6136),
.B(n_70),
.Y(n_6160)
);

INVx2_ASAP7_75t_L g6161 ( 
.A(n_5994),
.Y(n_6161)
);

AND2x2_ASAP7_75t_L g6162 ( 
.A(n_5998),
.B(n_70),
.Y(n_6162)
);

AO21x2_ASAP7_75t_L g6163 ( 
.A1(n_6070),
.A2(n_70),
.B(n_71),
.Y(n_6163)
);

OAI21xp5_ASAP7_75t_L g6164 ( 
.A1(n_6106),
.A2(n_71),
.B(n_72),
.Y(n_6164)
);

AOI211xp5_ASAP7_75t_SL g6165 ( 
.A1(n_6077),
.A2(n_741),
.B(n_742),
.C(n_740),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_6039),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_6039),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_6079),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_6007),
.Y(n_6169)
);

AOI21x1_ASAP7_75t_L g6170 ( 
.A1(n_6073),
.A2(n_71),
.B(n_72),
.Y(n_6170)
);

OR2x6_ASAP7_75t_L g6171 ( 
.A(n_5991),
.B(n_740),
.Y(n_6171)
);

AO21x2_ASAP7_75t_L g6172 ( 
.A1(n_6094),
.A2(n_71),
.B(n_72),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_6096),
.Y(n_6173)
);

AND2x2_ASAP7_75t_L g6174 ( 
.A(n_6044),
.B(n_73),
.Y(n_6174)
);

INVx2_ASAP7_75t_SL g6175 ( 
.A(n_6113),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_6112),
.Y(n_6176)
);

INVxp33_ASAP7_75t_L g6177 ( 
.A(n_6126),
.Y(n_6177)
);

OAI21xp5_ASAP7_75t_L g6178 ( 
.A1(n_6025),
.A2(n_73),
.B(n_74),
.Y(n_6178)
);

INVx3_ASAP7_75t_L g6179 ( 
.A(n_5992),
.Y(n_6179)
);

AND2x2_ASAP7_75t_L g6180 ( 
.A(n_5989),
.B(n_6117),
.Y(n_6180)
);

INVx2_ASAP7_75t_L g6181 ( 
.A(n_6115),
.Y(n_6181)
);

AND2x4_ASAP7_75t_L g6182 ( 
.A(n_6119),
.B(n_740),
.Y(n_6182)
);

HB1xp67_ASAP7_75t_L g6183 ( 
.A(n_6140),
.Y(n_6183)
);

INVx2_ASAP7_75t_L g6184 ( 
.A(n_6009),
.Y(n_6184)
);

INVx2_ASAP7_75t_L g6185 ( 
.A(n_6057),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_6086),
.Y(n_6186)
);

INVx2_ASAP7_75t_SL g6187 ( 
.A(n_6113),
.Y(n_6187)
);

INVx2_ASAP7_75t_L g6188 ( 
.A(n_6034),
.Y(n_6188)
);

HB1xp67_ASAP7_75t_L g6189 ( 
.A(n_6097),
.Y(n_6189)
);

AND2x2_ASAP7_75t_L g6190 ( 
.A(n_6016),
.B(n_73),
.Y(n_6190)
);

AND2x2_ASAP7_75t_L g6191 ( 
.A(n_5987),
.B(n_73),
.Y(n_6191)
);

INVx2_ASAP7_75t_L g6192 ( 
.A(n_6059),
.Y(n_6192)
);

AND2x2_ASAP7_75t_L g6193 ( 
.A(n_6084),
.B(n_74),
.Y(n_6193)
);

INVx2_ASAP7_75t_L g6194 ( 
.A(n_6045),
.Y(n_6194)
);

INVxp67_ASAP7_75t_L g6195 ( 
.A(n_6109),
.Y(n_6195)
);

INVx2_ASAP7_75t_L g6196 ( 
.A(n_6099),
.Y(n_6196)
);

AND2x4_ASAP7_75t_L g6197 ( 
.A(n_6119),
.B(n_741),
.Y(n_6197)
);

AOI22xp33_ASAP7_75t_L g6198 ( 
.A1(n_6107),
.A2(n_742),
.B1(n_743),
.B2(n_741),
.Y(n_6198)
);

OR2x6_ASAP7_75t_L g6199 ( 
.A(n_6032),
.B(n_743),
.Y(n_6199)
);

NAND5xp2_ASAP7_75t_SL g6200 ( 
.A(n_6131),
.B(n_76),
.C(n_74),
.D(n_75),
.E(n_77),
.Y(n_6200)
);

AND2x2_ASAP7_75t_L g6201 ( 
.A(n_6074),
.B(n_75),
.Y(n_6201)
);

NAND2xp5_ASAP7_75t_L g6202 ( 
.A(n_6090),
.B(n_76),
.Y(n_6202)
);

INVx1_ASAP7_75t_L g6203 ( 
.A(n_6048),
.Y(n_6203)
);

OAI211xp5_ASAP7_75t_L g6204 ( 
.A1(n_6121),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_6204)
);

INVx2_ASAP7_75t_L g6205 ( 
.A(n_6066),
.Y(n_6205)
);

INVx2_ASAP7_75t_L g6206 ( 
.A(n_6139),
.Y(n_6206)
);

NAND4xp25_ASAP7_75t_L g6207 ( 
.A(n_6001),
.B(n_78),
.C(n_76),
.D(n_77),
.Y(n_6207)
);

AOI22xp33_ASAP7_75t_L g6208 ( 
.A1(n_6108),
.A2(n_744),
.B1(n_745),
.B2(n_743),
.Y(n_6208)
);

BUFx2_ASAP7_75t_L g6209 ( 
.A(n_5997),
.Y(n_6209)
);

AND2x2_ASAP7_75t_L g6210 ( 
.A(n_6035),
.B(n_78),
.Y(n_6210)
);

HB1xp67_ASAP7_75t_L g6211 ( 
.A(n_6116),
.Y(n_6211)
);

OR2x6_ASAP7_75t_L g6212 ( 
.A(n_6010),
.B(n_744),
.Y(n_6212)
);

INVx2_ASAP7_75t_L g6213 ( 
.A(n_6058),
.Y(n_6213)
);

INVx1_ASAP7_75t_L g6214 ( 
.A(n_6043),
.Y(n_6214)
);

BUFx3_ASAP7_75t_L g6215 ( 
.A(n_6015),
.Y(n_6215)
);

AND2x2_ASAP7_75t_L g6216 ( 
.A(n_6111),
.B(n_78),
.Y(n_6216)
);

INVx1_ASAP7_75t_SL g6217 ( 
.A(n_6028),
.Y(n_6217)
);

INVx1_ASAP7_75t_L g6218 ( 
.A(n_6088),
.Y(n_6218)
);

OA21x2_ASAP7_75t_L g6219 ( 
.A1(n_6080),
.A2(n_79),
.B(n_80),
.Y(n_6219)
);

NOR2xp33_ASAP7_75t_L g6220 ( 
.A(n_6127),
.B(n_79),
.Y(n_6220)
);

INVxp67_ASAP7_75t_L g6221 ( 
.A(n_6021),
.Y(n_6221)
);

INVx2_ASAP7_75t_L g6222 ( 
.A(n_6020),
.Y(n_6222)
);

INVx2_ASAP7_75t_SL g6223 ( 
.A(n_6012),
.Y(n_6223)
);

INVx3_ASAP7_75t_L g6224 ( 
.A(n_6037),
.Y(n_6224)
);

AND2x2_ASAP7_75t_L g6225 ( 
.A(n_6075),
.B(n_79),
.Y(n_6225)
);

INVx2_ASAP7_75t_L g6226 ( 
.A(n_6022),
.Y(n_6226)
);

BUFx3_ASAP7_75t_L g6227 ( 
.A(n_6014),
.Y(n_6227)
);

OAI21xp5_ASAP7_75t_L g6228 ( 
.A1(n_6144),
.A2(n_80),
.B(n_81),
.Y(n_6228)
);

OR2x6_ASAP7_75t_L g6229 ( 
.A(n_6067),
.B(n_6068),
.Y(n_6229)
);

AND2x6_ASAP7_75t_L g6230 ( 
.A(n_6024),
.B(n_745),
.Y(n_6230)
);

OR2x6_ASAP7_75t_L g6231 ( 
.A(n_6067),
.B(n_745),
.Y(n_6231)
);

OAI221xp5_ASAP7_75t_L g6232 ( 
.A1(n_6149),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.C(n_83),
.Y(n_6232)
);

BUFx2_ASAP7_75t_L g6233 ( 
.A(n_6060),
.Y(n_6233)
);

NAND2xp5_ASAP7_75t_L g6234 ( 
.A(n_6055),
.B(n_80),
.Y(n_6234)
);

INVx2_ASAP7_75t_L g6235 ( 
.A(n_6029),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_6091),
.Y(n_6236)
);

OR2x2_ASAP7_75t_L g6237 ( 
.A(n_6008),
.B(n_81),
.Y(n_6237)
);

AOI21x1_ASAP7_75t_L g6238 ( 
.A1(n_6093),
.A2(n_81),
.B(n_82),
.Y(n_6238)
);

AND2x2_ASAP7_75t_L g6239 ( 
.A(n_6072),
.B(n_82),
.Y(n_6239)
);

INVx1_ASAP7_75t_L g6240 ( 
.A(n_6005),
.Y(n_6240)
);

AND2x2_ASAP7_75t_L g6241 ( 
.A(n_6049),
.B(n_83),
.Y(n_6241)
);

OA21x2_ASAP7_75t_L g6242 ( 
.A1(n_6053),
.A2(n_83),
.B(n_84),
.Y(n_6242)
);

INVx2_ASAP7_75t_L g6243 ( 
.A(n_6040),
.Y(n_6243)
);

INVx2_ASAP7_75t_L g6244 ( 
.A(n_6041),
.Y(n_6244)
);

NAND2xp5_ASAP7_75t_L g6245 ( 
.A(n_6051),
.B(n_83),
.Y(n_6245)
);

INVx2_ASAP7_75t_L g6246 ( 
.A(n_6042),
.Y(n_6246)
);

OAI21x1_ASAP7_75t_L g6247 ( 
.A1(n_6004),
.A2(n_747),
.B(n_746),
.Y(n_6247)
);

AND2x2_ASAP7_75t_L g6248 ( 
.A(n_6063),
.B(n_84),
.Y(n_6248)
);

AND2x2_ASAP7_75t_L g6249 ( 
.A(n_6006),
.B(n_84),
.Y(n_6249)
);

OA21x2_ASAP7_75t_L g6250 ( 
.A1(n_6003),
.A2(n_84),
.B(n_85),
.Y(n_6250)
);

INVx1_ASAP7_75t_L g6251 ( 
.A(n_6147),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_6150),
.Y(n_6252)
);

BUFx2_ASAP7_75t_L g6253 ( 
.A(n_6060),
.Y(n_6253)
);

AO21x2_ASAP7_75t_L g6254 ( 
.A1(n_6135),
.A2(n_85),
.B(n_86),
.Y(n_6254)
);

HB1xp67_ASAP7_75t_L g6255 ( 
.A(n_6116),
.Y(n_6255)
);

OA21x2_ASAP7_75t_L g6256 ( 
.A1(n_6114),
.A2(n_86),
.B(n_87),
.Y(n_6256)
);

AND2x2_ASAP7_75t_L g6257 ( 
.A(n_6023),
.B(n_87),
.Y(n_6257)
);

INVx1_ASAP7_75t_SL g6258 ( 
.A(n_6142),
.Y(n_6258)
);

HB1xp67_ASAP7_75t_L g6259 ( 
.A(n_6128),
.Y(n_6259)
);

INVx3_ASAP7_75t_L g6260 ( 
.A(n_6056),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_5996),
.Y(n_6261)
);

INVx2_ASAP7_75t_L g6262 ( 
.A(n_6148),
.Y(n_6262)
);

AND2x4_ASAP7_75t_L g6263 ( 
.A(n_5990),
.B(n_746),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_6128),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5999),
.Y(n_6265)
);

INVx2_ASAP7_75t_L g6266 ( 
.A(n_6146),
.Y(n_6266)
);

INVx2_ASAP7_75t_L g6267 ( 
.A(n_6118),
.Y(n_6267)
);

NAND2xp5_ASAP7_75t_L g6268 ( 
.A(n_6123),
.B(n_87),
.Y(n_6268)
);

AND2x2_ASAP7_75t_L g6269 ( 
.A(n_6017),
.B(n_87),
.Y(n_6269)
);

AND2x2_ASAP7_75t_L g6270 ( 
.A(n_6026),
.B(n_88),
.Y(n_6270)
);

INVx2_ASAP7_75t_L g6271 ( 
.A(n_6124),
.Y(n_6271)
);

INVx1_ASAP7_75t_L g6272 ( 
.A(n_6130),
.Y(n_6272)
);

AND2x2_ASAP7_75t_L g6273 ( 
.A(n_6054),
.B(n_6064),
.Y(n_6273)
);

AND2x2_ASAP7_75t_L g6274 ( 
.A(n_6141),
.B(n_88),
.Y(n_6274)
);

INVxp67_ASAP7_75t_L g6275 ( 
.A(n_6033),
.Y(n_6275)
);

AO21x2_ASAP7_75t_L g6276 ( 
.A1(n_6120),
.A2(n_88),
.B(n_89),
.Y(n_6276)
);

AO21x2_ASAP7_75t_L g6277 ( 
.A1(n_6071),
.A2(n_88),
.B(n_89),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_6143),
.Y(n_6278)
);

OAI21xp5_ASAP7_75t_L g6279 ( 
.A1(n_5988),
.A2(n_89),
.B(n_90),
.Y(n_6279)
);

HB1xp67_ASAP7_75t_L g6280 ( 
.A(n_6145),
.Y(n_6280)
);

AND2x2_ASAP7_75t_L g6281 ( 
.A(n_6013),
.B(n_89),
.Y(n_6281)
);

INVxp67_ASAP7_75t_L g6282 ( 
.A(n_6104),
.Y(n_6282)
);

INVx3_ASAP7_75t_L g6283 ( 
.A(n_6046),
.Y(n_6283)
);

INVx1_ASAP7_75t_L g6284 ( 
.A(n_6125),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_6132),
.Y(n_6285)
);

AOI22xp33_ASAP7_75t_L g6286 ( 
.A1(n_6095),
.A2(n_747),
.B1(n_749),
.B2(n_746),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_6133),
.Y(n_6287)
);

AND2x2_ASAP7_75t_L g6288 ( 
.A(n_6082),
.B(n_90),
.Y(n_6288)
);

OR2x6_ASAP7_75t_L g6289 ( 
.A(n_6137),
.B(n_750),
.Y(n_6289)
);

INVx1_ASAP7_75t_L g6290 ( 
.A(n_6085),
.Y(n_6290)
);

AND2x2_ASAP7_75t_L g6291 ( 
.A(n_6069),
.B(n_90),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_6038),
.Y(n_6292)
);

INVx2_ASAP7_75t_L g6293 ( 
.A(n_5995),
.Y(n_6293)
);

AO21x2_ASAP7_75t_L g6294 ( 
.A1(n_6062),
.A2(n_90),
.B(n_91),
.Y(n_6294)
);

AO21x2_ASAP7_75t_L g6295 ( 
.A1(n_6105),
.A2(n_91),
.B(n_92),
.Y(n_6295)
);

AND2x2_ASAP7_75t_L g6296 ( 
.A(n_6078),
.B(n_91),
.Y(n_6296)
);

INVx2_ASAP7_75t_L g6297 ( 
.A(n_5995),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_6087),
.B(n_91),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6076),
.Y(n_6299)
);

OAI221xp5_ASAP7_75t_L g6300 ( 
.A1(n_6000),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.C(n_95),
.Y(n_6300)
);

INVx2_ASAP7_75t_L g6301 ( 
.A(n_6019),
.Y(n_6301)
);

BUFx3_ASAP7_75t_L g6302 ( 
.A(n_6100),
.Y(n_6302)
);

AND2x2_ASAP7_75t_L g6303 ( 
.A(n_6036),
.B(n_6030),
.Y(n_6303)
);

INVx2_ASAP7_75t_L g6304 ( 
.A(n_6052),
.Y(n_6304)
);

AND2x2_ASAP7_75t_L g6305 ( 
.A(n_6031),
.B(n_6002),
.Y(n_6305)
);

INVx2_ASAP7_75t_L g6306 ( 
.A(n_6083),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_6061),
.Y(n_6307)
);

BUFx2_ASAP7_75t_L g6308 ( 
.A(n_6092),
.Y(n_6308)
);

AOI21xp33_ASAP7_75t_L g6309 ( 
.A1(n_6101),
.A2(n_92),
.B(n_93),
.Y(n_6309)
);

HB1xp67_ASAP7_75t_L g6310 ( 
.A(n_6103),
.Y(n_6310)
);

BUFx3_ASAP7_75t_L g6311 ( 
.A(n_6098),
.Y(n_6311)
);

OR2x6_ASAP7_75t_L g6312 ( 
.A(n_6018),
.B(n_750),
.Y(n_6312)
);

BUFx6f_ASAP7_75t_L g6313 ( 
.A(n_6081),
.Y(n_6313)
);

INVx2_ASAP7_75t_L g6314 ( 
.A(n_6050),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6047),
.Y(n_6315)
);

AND2x2_ASAP7_75t_L g6316 ( 
.A(n_6065),
.B(n_93),
.Y(n_6316)
);

INVx1_ASAP7_75t_L g6317 ( 
.A(n_6102),
.Y(n_6317)
);

NAND2xp5_ASAP7_75t_SL g6318 ( 
.A(n_6011),
.B(n_93),
.Y(n_6318)
);

AND2x2_ASAP7_75t_L g6319 ( 
.A(n_6110),
.B(n_94),
.Y(n_6319)
);

BUFx3_ASAP7_75t_L g6320 ( 
.A(n_5991),
.Y(n_6320)
);

OR2x6_ASAP7_75t_L g6321 ( 
.A(n_6138),
.B(n_751),
.Y(n_6321)
);

INVx2_ASAP7_75t_L g6322 ( 
.A(n_6110),
.Y(n_6322)
);

INVx2_ASAP7_75t_SL g6323 ( 
.A(n_6138),
.Y(n_6323)
);

OA21x2_ASAP7_75t_L g6324 ( 
.A1(n_6089),
.A2(n_94),
.B(n_95),
.Y(n_6324)
);

CKINVDCx5p33_ASAP7_75t_R g6325 ( 
.A(n_6126),
.Y(n_6325)
);

OA21x2_ASAP7_75t_L g6326 ( 
.A1(n_6089),
.A2(n_94),
.B(n_95),
.Y(n_6326)
);

AOI21xp5_ASAP7_75t_L g6327 ( 
.A1(n_6106),
.A2(n_95),
.B(n_96),
.Y(n_6327)
);

INVx1_ASAP7_75t_L g6328 ( 
.A(n_6110),
.Y(n_6328)
);

OAI222xp33_ASAP7_75t_L g6329 ( 
.A1(n_5993),
.A2(n_98),
.B1(n_100),
.B2(n_96),
.C1(n_97),
.C2(n_99),
.Y(n_6329)
);

INVx11_ASAP7_75t_L g6330 ( 
.A(n_5991),
.Y(n_6330)
);

AOI22xp5_ASAP7_75t_L g6331 ( 
.A1(n_6209),
.A2(n_6224),
.B1(n_6263),
.B2(n_6301),
.Y(n_6331)
);

INVx2_ASAP7_75t_L g6332 ( 
.A(n_6322),
.Y(n_6332)
);

INVx2_ASAP7_75t_SL g6333 ( 
.A(n_6330),
.Y(n_6333)
);

NAND2xp5_ASAP7_75t_L g6334 ( 
.A(n_6209),
.B(n_96),
.Y(n_6334)
);

AND2x2_ASAP7_75t_L g6335 ( 
.A(n_6323),
.B(n_96),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_6158),
.Y(n_6336)
);

AND2x4_ASAP7_75t_L g6337 ( 
.A(n_6181),
.B(n_751),
.Y(n_6337)
);

INVx1_ASAP7_75t_L g6338 ( 
.A(n_6162),
.Y(n_6338)
);

AND2x4_ASAP7_75t_L g6339 ( 
.A(n_6161),
.B(n_752),
.Y(n_6339)
);

AOI22xp33_ASAP7_75t_L g6340 ( 
.A1(n_6188),
.A2(n_753),
.B1(n_754),
.B2(n_752),
.Y(n_6340)
);

NAND2xp5_ASAP7_75t_L g6341 ( 
.A(n_6310),
.B(n_97),
.Y(n_6341)
);

INVx1_ASAP7_75t_L g6342 ( 
.A(n_6152),
.Y(n_6342)
);

NOR2xp33_ASAP7_75t_L g6343 ( 
.A(n_6177),
.B(n_97),
.Y(n_6343)
);

AND2x2_ASAP7_75t_L g6344 ( 
.A(n_6180),
.B(n_98),
.Y(n_6344)
);

INVx2_ASAP7_75t_L g6345 ( 
.A(n_6153),
.Y(n_6345)
);

BUFx6f_ASAP7_75t_L g6346 ( 
.A(n_6320),
.Y(n_6346)
);

AND2x2_ASAP7_75t_L g6347 ( 
.A(n_6283),
.B(n_98),
.Y(n_6347)
);

INVx2_ASAP7_75t_L g6348 ( 
.A(n_6155),
.Y(n_6348)
);

AND2x2_ASAP7_75t_L g6349 ( 
.A(n_6175),
.B(n_99),
.Y(n_6349)
);

HB1xp67_ASAP7_75t_L g6350 ( 
.A(n_6189),
.Y(n_6350)
);

AND2x2_ASAP7_75t_L g6351 ( 
.A(n_6187),
.B(n_99),
.Y(n_6351)
);

NAND2xp5_ASAP7_75t_L g6352 ( 
.A(n_6191),
.B(n_100),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_6319),
.Y(n_6353)
);

NAND2xp5_ASAP7_75t_L g6354 ( 
.A(n_6315),
.B(n_100),
.Y(n_6354)
);

NAND2xp5_ASAP7_75t_L g6355 ( 
.A(n_6221),
.B(n_100),
.Y(n_6355)
);

AND2x2_ASAP7_75t_L g6356 ( 
.A(n_6260),
.B(n_101),
.Y(n_6356)
);

INVx1_ASAP7_75t_L g6357 ( 
.A(n_6239),
.Y(n_6357)
);

NOR2x1_ASAP7_75t_L g6358 ( 
.A(n_6229),
.B(n_101),
.Y(n_6358)
);

INVx1_ASAP7_75t_L g6359 ( 
.A(n_6151),
.Y(n_6359)
);

AND2x2_ASAP7_75t_L g6360 ( 
.A(n_6229),
.B(n_101),
.Y(n_6360)
);

NAND2xp5_ASAP7_75t_L g6361 ( 
.A(n_6293),
.B(n_101),
.Y(n_6361)
);

INVx1_ASAP7_75t_L g6362 ( 
.A(n_6328),
.Y(n_6362)
);

AND2x2_ASAP7_75t_L g6363 ( 
.A(n_6210),
.B(n_102),
.Y(n_6363)
);

INVx3_ASAP7_75t_L g6364 ( 
.A(n_6325),
.Y(n_6364)
);

AND2x2_ASAP7_75t_L g6365 ( 
.A(n_6216),
.B(n_6183),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_6156),
.Y(n_6366)
);

INVx2_ASAP7_75t_L g6367 ( 
.A(n_6185),
.Y(n_6367)
);

AOI222xp33_ASAP7_75t_L g6368 ( 
.A1(n_6297),
.A2(n_756),
.B1(n_754),
.B2(n_757),
.C1(n_755),
.C2(n_753),
.Y(n_6368)
);

BUFx2_ASAP7_75t_L g6369 ( 
.A(n_6263),
.Y(n_6369)
);

AND2x4_ASAP7_75t_L g6370 ( 
.A(n_6215),
.B(n_754),
.Y(n_6370)
);

NAND2xp5_ASAP7_75t_L g6371 ( 
.A(n_6299),
.B(n_102),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_6219),
.Y(n_6372)
);

AND2x2_ASAP7_75t_L g6373 ( 
.A(n_6223),
.B(n_102),
.Y(n_6373)
);

HB1xp67_ASAP7_75t_L g6374 ( 
.A(n_6169),
.Y(n_6374)
);

INVx1_ASAP7_75t_SL g6375 ( 
.A(n_6217),
.Y(n_6375)
);

BUFx2_ASAP7_75t_L g6376 ( 
.A(n_6282),
.Y(n_6376)
);

AND2x2_ASAP7_75t_L g6377 ( 
.A(n_6258),
.B(n_102),
.Y(n_6377)
);

INVxp67_ASAP7_75t_SL g6378 ( 
.A(n_6220),
.Y(n_6378)
);

INVx2_ASAP7_75t_L g6379 ( 
.A(n_6231),
.Y(n_6379)
);

INVx1_ASAP7_75t_L g6380 ( 
.A(n_6219),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_6233),
.Y(n_6381)
);

AND2x4_ASAP7_75t_L g6382 ( 
.A(n_6179),
.B(n_6206),
.Y(n_6382)
);

HB1xp67_ASAP7_75t_L g6383 ( 
.A(n_6172),
.Y(n_6383)
);

AOI22xp33_ASAP7_75t_L g6384 ( 
.A1(n_6302),
.A2(n_756),
.B1(n_758),
.B2(n_755),
.Y(n_6384)
);

INVx1_ASAP7_75t_L g6385 ( 
.A(n_6233),
.Y(n_6385)
);

HB1xp67_ASAP7_75t_L g6386 ( 
.A(n_6163),
.Y(n_6386)
);

AND2x2_ASAP7_75t_L g6387 ( 
.A(n_6195),
.B(n_103),
.Y(n_6387)
);

AND2x2_ASAP7_75t_L g6388 ( 
.A(n_6304),
.B(n_103),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_6253),
.Y(n_6389)
);

INVx3_ASAP7_75t_L g6390 ( 
.A(n_6171),
.Y(n_6390)
);

OR2x2_ASAP7_75t_L g6391 ( 
.A(n_6306),
.B(n_103),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6253),
.Y(n_6392)
);

NOR2xp33_ASAP7_75t_L g6393 ( 
.A(n_6308),
.B(n_103),
.Y(n_6393)
);

INVx2_ASAP7_75t_L g6394 ( 
.A(n_6231),
.Y(n_6394)
);

AND2x2_ASAP7_75t_L g6395 ( 
.A(n_6314),
.B(n_104),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_6201),
.Y(n_6396)
);

NAND2xp5_ASAP7_75t_L g6397 ( 
.A(n_6317),
.B(n_104),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_6225),
.Y(n_6398)
);

INVx3_ASAP7_75t_L g6399 ( 
.A(n_6171),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_6211),
.Y(n_6400)
);

AND2x2_ASAP7_75t_L g6401 ( 
.A(n_6290),
.B(n_104),
.Y(n_6401)
);

INVx1_ASAP7_75t_L g6402 ( 
.A(n_6255),
.Y(n_6402)
);

OR2x2_ASAP7_75t_L g6403 ( 
.A(n_6284),
.B(n_104),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_6259),
.Y(n_6404)
);

INVx2_ASAP7_75t_L g6405 ( 
.A(n_6174),
.Y(n_6405)
);

OAI221xp5_ASAP7_75t_SL g6406 ( 
.A1(n_6308),
.A2(n_758),
.B1(n_759),
.B2(n_756),
.C(n_755),
.Y(n_6406)
);

AND2x2_ASAP7_75t_L g6407 ( 
.A(n_6227),
.B(n_105),
.Y(n_6407)
);

INVx2_ASAP7_75t_L g6408 ( 
.A(n_6182),
.Y(n_6408)
);

INVx4_ASAP7_75t_L g6409 ( 
.A(n_6157),
.Y(n_6409)
);

BUFx3_ASAP7_75t_L g6410 ( 
.A(n_6190),
.Y(n_6410)
);

BUFx3_ASAP7_75t_L g6411 ( 
.A(n_6157),
.Y(n_6411)
);

NAND3xp33_ASAP7_75t_L g6412 ( 
.A(n_6165),
.B(n_105),
.C(n_106),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_6182),
.Y(n_6413)
);

INVx2_ASAP7_75t_L g6414 ( 
.A(n_6312),
.Y(n_6414)
);

NAND2xp5_ASAP7_75t_L g6415 ( 
.A(n_6307),
.B(n_105),
.Y(n_6415)
);

INVx2_ASAP7_75t_L g6416 ( 
.A(n_6312),
.Y(n_6416)
);

OR2x6_ASAP7_75t_SL g6417 ( 
.A(n_6234),
.B(n_761),
.Y(n_6417)
);

BUFx3_ASAP7_75t_L g6418 ( 
.A(n_6159),
.Y(n_6418)
);

INVxp67_ASAP7_75t_SL g6419 ( 
.A(n_6170),
.Y(n_6419)
);

BUFx3_ASAP7_75t_L g6420 ( 
.A(n_6159),
.Y(n_6420)
);

AND2x2_ASAP7_75t_L g6421 ( 
.A(n_6285),
.B(n_105),
.Y(n_6421)
);

OR2x2_ASAP7_75t_L g6422 ( 
.A(n_6287),
.B(n_6292),
.Y(n_6422)
);

AO21x2_ASAP7_75t_L g6423 ( 
.A1(n_6173),
.A2(n_106),
.B(n_107),
.Y(n_6423)
);

AND2x2_ASAP7_75t_L g6424 ( 
.A(n_6176),
.B(n_106),
.Y(n_6424)
);

HB1xp67_ASAP7_75t_L g6425 ( 
.A(n_6242),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6160),
.Y(n_6426)
);

NAND2xp5_ASAP7_75t_L g6427 ( 
.A(n_6275),
.B(n_106),
.Y(n_6427)
);

AND2x2_ASAP7_75t_L g6428 ( 
.A(n_6214),
.B(n_107),
.Y(n_6428)
);

INVx2_ASAP7_75t_L g6429 ( 
.A(n_6196),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_6166),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6167),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_6242),
.Y(n_6432)
);

AOI222xp33_ASAP7_75t_L g6433 ( 
.A1(n_6311),
.A2(n_762),
.B1(n_760),
.B2(n_763),
.C1(n_761),
.C2(n_759),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_6250),
.Y(n_6434)
);

INVx1_ASAP7_75t_L g6435 ( 
.A(n_6250),
.Y(n_6435)
);

INVx2_ASAP7_75t_L g6436 ( 
.A(n_6205),
.Y(n_6436)
);

INVx1_ASAP7_75t_L g6437 ( 
.A(n_6154),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_6240),
.B(n_107),
.Y(n_6438)
);

INVx1_ASAP7_75t_L g6439 ( 
.A(n_6154),
.Y(n_6439)
);

BUFx2_ASAP7_75t_L g6440 ( 
.A(n_6324),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_6324),
.Y(n_6441)
);

AND2x2_ASAP7_75t_L g6442 ( 
.A(n_6251),
.B(n_107),
.Y(n_6442)
);

NOR2x1_ASAP7_75t_L g6443 ( 
.A(n_6321),
.B(n_6277),
.Y(n_6443)
);

NAND2xp5_ASAP7_75t_SL g6444 ( 
.A(n_6327),
.B(n_108),
.Y(n_6444)
);

OR2x2_ASAP7_75t_L g6445 ( 
.A(n_6203),
.B(n_6252),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6326),
.Y(n_6446)
);

AND2x4_ASAP7_75t_SL g6447 ( 
.A(n_6321),
.B(n_108),
.Y(n_6447)
);

AND2x4_ASAP7_75t_L g6448 ( 
.A(n_6197),
.B(n_109),
.Y(n_6448)
);

INVx1_ASAP7_75t_L g6449 ( 
.A(n_6326),
.Y(n_6449)
);

AND2x4_ASAP7_75t_L g6450 ( 
.A(n_6168),
.B(n_6186),
.Y(n_6450)
);

OR2x2_ASAP7_75t_L g6451 ( 
.A(n_6194),
.B(n_108),
.Y(n_6451)
);

AND2x2_ASAP7_75t_L g6452 ( 
.A(n_6273),
.B(n_108),
.Y(n_6452)
);

NAND2xp5_ASAP7_75t_L g6453 ( 
.A(n_6303),
.B(n_109),
.Y(n_6453)
);

AND2x4_ASAP7_75t_L g6454 ( 
.A(n_6279),
.B(n_759),
.Y(n_6454)
);

NOR2xp33_ASAP7_75t_L g6455 ( 
.A(n_6313),
.B(n_109),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6247),
.Y(n_6456)
);

INVx1_ASAP7_75t_L g6457 ( 
.A(n_6274),
.Y(n_6457)
);

AND2x2_ASAP7_75t_L g6458 ( 
.A(n_6248),
.B(n_109),
.Y(n_6458)
);

BUFx3_ASAP7_75t_L g6459 ( 
.A(n_6212),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6280),
.Y(n_6460)
);

INVx1_ASAP7_75t_L g6461 ( 
.A(n_6264),
.Y(n_6461)
);

BUFx2_ASAP7_75t_L g6462 ( 
.A(n_6212),
.Y(n_6462)
);

NAND2xp5_ASAP7_75t_L g6463 ( 
.A(n_6305),
.B(n_110),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_6241),
.Y(n_6464)
);

AND2x2_ASAP7_75t_L g6465 ( 
.A(n_6298),
.B(n_110),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6238),
.Y(n_6466)
);

AOI22xp33_ASAP7_75t_L g6467 ( 
.A1(n_6313),
.A2(n_761),
.B1(n_762),
.B2(n_760),
.Y(n_6467)
);

AND2x2_ASAP7_75t_L g6468 ( 
.A(n_6256),
.B(n_110),
.Y(n_6468)
);

AND2x2_ASAP7_75t_L g6469 ( 
.A(n_6256),
.B(n_111),
.Y(n_6469)
);

BUFx6f_ASAP7_75t_L g6470 ( 
.A(n_6199),
.Y(n_6470)
);

NOR2xp67_ASAP7_75t_SL g6471 ( 
.A(n_6232),
.B(n_763),
.Y(n_6471)
);

BUFx2_ASAP7_75t_L g6472 ( 
.A(n_6218),
.Y(n_6472)
);

INVx1_ASAP7_75t_L g6473 ( 
.A(n_6238),
.Y(n_6473)
);

INVx2_ASAP7_75t_L g6474 ( 
.A(n_6192),
.Y(n_6474)
);

NOR3xp33_ASAP7_75t_L g6475 ( 
.A(n_6329),
.B(n_111),
.C(n_112),
.Y(n_6475)
);

OR2x2_ASAP7_75t_L g6476 ( 
.A(n_6245),
.B(n_111),
.Y(n_6476)
);

AND2x2_ASAP7_75t_L g6477 ( 
.A(n_6193),
.B(n_111),
.Y(n_6477)
);

INVx1_ASAP7_75t_L g6478 ( 
.A(n_6236),
.Y(n_6478)
);

AND2x2_ASAP7_75t_L g6479 ( 
.A(n_6288),
.B(n_112),
.Y(n_6479)
);

AND2x2_ASAP7_75t_L g6480 ( 
.A(n_6291),
.B(n_112),
.Y(n_6480)
);

AND2x4_ASAP7_75t_L g6481 ( 
.A(n_6254),
.B(n_113),
.Y(n_6481)
);

AND2x2_ASAP7_75t_L g6482 ( 
.A(n_6249),
.B(n_112),
.Y(n_6482)
);

AOI22xp33_ASAP7_75t_L g6483 ( 
.A1(n_6230),
.A2(n_764),
.B1(n_765),
.B2(n_763),
.Y(n_6483)
);

INVxp33_ASAP7_75t_SL g6484 ( 
.A(n_6296),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_6213),
.Y(n_6485)
);

AND2x2_ASAP7_75t_L g6486 ( 
.A(n_6281),
.B(n_113),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6202),
.Y(n_6487)
);

INVx5_ASAP7_75t_SL g6488 ( 
.A(n_6199),
.Y(n_6488)
);

AND2x2_ASAP7_75t_L g6489 ( 
.A(n_6269),
.B(n_114),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_6222),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_6226),
.Y(n_6491)
);

INVx2_ASAP7_75t_L g6492 ( 
.A(n_6289),
.Y(n_6492)
);

NAND2xp5_ASAP7_75t_L g6493 ( 
.A(n_6230),
.B(n_114),
.Y(n_6493)
);

INVx4_ASAP7_75t_L g6494 ( 
.A(n_6294),
.Y(n_6494)
);

NAND2xp5_ASAP7_75t_L g6495 ( 
.A(n_6230),
.B(n_114),
.Y(n_6495)
);

INVx1_ASAP7_75t_L g6496 ( 
.A(n_6235),
.Y(n_6496)
);

INVx2_ASAP7_75t_SL g6497 ( 
.A(n_6237),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_6243),
.Y(n_6498)
);

AND2x2_ASAP7_75t_L g6499 ( 
.A(n_6257),
.B(n_115),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_6244),
.Y(n_6500)
);

AND2x2_ASAP7_75t_L g6501 ( 
.A(n_6270),
.B(n_115),
.Y(n_6501)
);

INVx1_ASAP7_75t_L g6502 ( 
.A(n_6246),
.Y(n_6502)
);

INVx4_ASAP7_75t_L g6503 ( 
.A(n_6289),
.Y(n_6503)
);

AND2x2_ASAP7_75t_L g6504 ( 
.A(n_6184),
.B(n_115),
.Y(n_6504)
);

OAI22xp5_ASAP7_75t_L g6505 ( 
.A1(n_6268),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_6505)
);

INVx2_ASAP7_75t_L g6506 ( 
.A(n_6375),
.Y(n_6506)
);

NAND2xp5_ASAP7_75t_L g6507 ( 
.A(n_6378),
.B(n_6393),
.Y(n_6507)
);

INVx2_ASAP7_75t_SL g6508 ( 
.A(n_6346),
.Y(n_6508)
);

HB1xp67_ASAP7_75t_L g6509 ( 
.A(n_6377),
.Y(n_6509)
);

INVx2_ASAP7_75t_L g6510 ( 
.A(n_6337),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_6373),
.Y(n_6511)
);

AND2x4_ASAP7_75t_L g6512 ( 
.A(n_6364),
.B(n_6170),
.Y(n_6512)
);

INVx5_ASAP7_75t_SL g6513 ( 
.A(n_6346),
.Y(n_6513)
);

AND2x2_ASAP7_75t_L g6514 ( 
.A(n_6333),
.B(n_6309),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_6349),
.Y(n_6515)
);

BUFx2_ASAP7_75t_L g6516 ( 
.A(n_6409),
.Y(n_6516)
);

BUFx2_ASAP7_75t_SL g6517 ( 
.A(n_6470),
.Y(n_6517)
);

INVx2_ASAP7_75t_L g6518 ( 
.A(n_6337),
.Y(n_6518)
);

AND2x2_ASAP7_75t_L g6519 ( 
.A(n_6382),
.B(n_6271),
.Y(n_6519)
);

INVx3_ASAP7_75t_L g6520 ( 
.A(n_6411),
.Y(n_6520)
);

INVx1_ASAP7_75t_L g6521 ( 
.A(n_6351),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_6347),
.Y(n_6522)
);

OR2x2_ASAP7_75t_L g6523 ( 
.A(n_6341),
.B(n_6295),
.Y(n_6523)
);

AND2x2_ASAP7_75t_L g6524 ( 
.A(n_6410),
.B(n_6278),
.Y(n_6524)
);

INVx2_ASAP7_75t_L g6525 ( 
.A(n_6335),
.Y(n_6525)
);

OR2x2_ASAP7_75t_L g6526 ( 
.A(n_6334),
.B(n_6261),
.Y(n_6526)
);

AND2x2_ASAP7_75t_L g6527 ( 
.A(n_6488),
.B(n_6262),
.Y(n_6527)
);

INVx1_ASAP7_75t_L g6528 ( 
.A(n_6356),
.Y(n_6528)
);

INVx1_ASAP7_75t_L g6529 ( 
.A(n_6360),
.Y(n_6529)
);

AND2x2_ASAP7_75t_L g6530 ( 
.A(n_6488),
.B(n_6266),
.Y(n_6530)
);

INVx1_ASAP7_75t_L g6531 ( 
.A(n_6376),
.Y(n_6531)
);

AND2x2_ASAP7_75t_L g6532 ( 
.A(n_6365),
.B(n_6267),
.Y(n_6532)
);

INVx2_ASAP7_75t_L g6533 ( 
.A(n_6339),
.Y(n_6533)
);

INVx1_ASAP7_75t_L g6534 ( 
.A(n_6376),
.Y(n_6534)
);

AOI22xp33_ASAP7_75t_SL g6535 ( 
.A1(n_6369),
.A2(n_6503),
.B1(n_6462),
.B2(n_6440),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_6344),
.Y(n_6536)
);

AND2x2_ASAP7_75t_L g6537 ( 
.A(n_6390),
.B(n_6265),
.Y(n_6537)
);

AND2x2_ASAP7_75t_L g6538 ( 
.A(n_6399),
.B(n_6272),
.Y(n_6538)
);

AND2x2_ASAP7_75t_L g6539 ( 
.A(n_6388),
.B(n_6276),
.Y(n_6539)
);

NAND2xp5_ASAP7_75t_L g6540 ( 
.A(n_6475),
.B(n_6164),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_6372),
.Y(n_6541)
);

INVx2_ASAP7_75t_L g6542 ( 
.A(n_6339),
.Y(n_6542)
);

AND2x2_ASAP7_75t_L g6543 ( 
.A(n_6418),
.B(n_6286),
.Y(n_6543)
);

INVx1_ASAP7_75t_L g6544 ( 
.A(n_6380),
.Y(n_6544)
);

NAND2xp5_ASAP7_75t_L g6545 ( 
.A(n_6481),
.B(n_6208),
.Y(n_6545)
);

INVx1_ASAP7_75t_L g6546 ( 
.A(n_6343),
.Y(n_6546)
);

AND2x2_ASAP7_75t_L g6547 ( 
.A(n_6420),
.B(n_6316),
.Y(n_6547)
);

AND2x2_ASAP7_75t_L g6548 ( 
.A(n_6414),
.B(n_6198),
.Y(n_6548)
);

INVx1_ASAP7_75t_L g6549 ( 
.A(n_6407),
.Y(n_6549)
);

AND2x2_ASAP7_75t_L g6550 ( 
.A(n_6416),
.B(n_6228),
.Y(n_6550)
);

INVx4_ASAP7_75t_L g6551 ( 
.A(n_6470),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_6494),
.B(n_6178),
.Y(n_6552)
);

NAND2xp5_ASAP7_75t_L g6553 ( 
.A(n_6419),
.B(n_6318),
.Y(n_6553)
);

AO21x2_ASAP7_75t_L g6554 ( 
.A1(n_6381),
.A2(n_6204),
.B(n_6300),
.Y(n_6554)
);

OR2x2_ASAP7_75t_SL g6555 ( 
.A(n_6425),
.B(n_6432),
.Y(n_6555)
);

INVx2_ASAP7_75t_L g6556 ( 
.A(n_6332),
.Y(n_6556)
);

INVx1_ASAP7_75t_L g6557 ( 
.A(n_6350),
.Y(n_6557)
);

INVx1_ASAP7_75t_L g6558 ( 
.A(n_6434),
.Y(n_6558)
);

HB1xp67_ASAP7_75t_L g6559 ( 
.A(n_6374),
.Y(n_6559)
);

AND2x2_ASAP7_75t_L g6560 ( 
.A(n_6462),
.B(n_116),
.Y(n_6560)
);

INVx1_ASAP7_75t_L g6561 ( 
.A(n_6435),
.Y(n_6561)
);

NOR2x1_ASAP7_75t_SL g6562 ( 
.A(n_6459),
.B(n_6379),
.Y(n_6562)
);

HB1xp67_ASAP7_75t_L g6563 ( 
.A(n_6345),
.Y(n_6563)
);

AND2x2_ASAP7_75t_L g6564 ( 
.A(n_6405),
.B(n_116),
.Y(n_6564)
);

INVx5_ASAP7_75t_SL g6565 ( 
.A(n_6370),
.Y(n_6565)
);

INVx1_ASAP7_75t_L g6566 ( 
.A(n_6440),
.Y(n_6566)
);

OR2x6_ASAP7_75t_L g6567 ( 
.A(n_6394),
.B(n_6200),
.Y(n_6567)
);

BUFx2_ASAP7_75t_L g6568 ( 
.A(n_6443),
.Y(n_6568)
);

INVx2_ASAP7_75t_L g6569 ( 
.A(n_6370),
.Y(n_6569)
);

INVx2_ASAP7_75t_SL g6570 ( 
.A(n_6447),
.Y(n_6570)
);

INVx2_ASAP7_75t_L g6571 ( 
.A(n_6348),
.Y(n_6571)
);

INVx1_ASAP7_75t_L g6572 ( 
.A(n_6391),
.Y(n_6572)
);

AND2x2_ASAP7_75t_L g6573 ( 
.A(n_6331),
.B(n_116),
.Y(n_6573)
);

AND2x2_ASAP7_75t_L g6574 ( 
.A(n_6492),
.B(n_117),
.Y(n_6574)
);

INVx2_ASAP7_75t_L g6575 ( 
.A(n_6367),
.Y(n_6575)
);

AND2x2_ASAP7_75t_L g6576 ( 
.A(n_6395),
.B(n_117),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6504),
.Y(n_6577)
);

AND2x2_ASAP7_75t_L g6578 ( 
.A(n_6396),
.B(n_117),
.Y(n_6578)
);

INVx2_ASAP7_75t_L g6579 ( 
.A(n_6474),
.Y(n_6579)
);

NAND2xp5_ASAP7_75t_L g6580 ( 
.A(n_6398),
.B(n_6207),
.Y(n_6580)
);

INVx3_ASAP7_75t_L g6581 ( 
.A(n_6408),
.Y(n_6581)
);

INVx2_ASAP7_75t_L g6582 ( 
.A(n_6413),
.Y(n_6582)
);

INVx2_ASAP7_75t_SL g6583 ( 
.A(n_6448),
.Y(n_6583)
);

NAND2xp5_ASAP7_75t_L g6584 ( 
.A(n_6497),
.B(n_118),
.Y(n_6584)
);

AND2x2_ASAP7_75t_L g6585 ( 
.A(n_6358),
.B(n_118),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_6437),
.Y(n_6586)
);

AND2x2_ASAP7_75t_L g6587 ( 
.A(n_6369),
.B(n_118),
.Y(n_6587)
);

INVx1_ASAP7_75t_SL g6588 ( 
.A(n_6451),
.Y(n_6588)
);

AO21x2_ASAP7_75t_L g6589 ( 
.A1(n_6385),
.A2(n_6200),
.B(n_119),
.Y(n_6589)
);

BUFx2_ASAP7_75t_L g6590 ( 
.A(n_6439),
.Y(n_6590)
);

AND2x2_ASAP7_75t_L g6591 ( 
.A(n_6401),
.B(n_6336),
.Y(n_6591)
);

NAND2xp5_ASAP7_75t_L g6592 ( 
.A(n_6484),
.B(n_119),
.Y(n_6592)
);

AND2x4_ASAP7_75t_L g6593 ( 
.A(n_6359),
.B(n_119),
.Y(n_6593)
);

HB1xp67_ASAP7_75t_L g6594 ( 
.A(n_6355),
.Y(n_6594)
);

INVx2_ASAP7_75t_L g6595 ( 
.A(n_6429),
.Y(n_6595)
);

AND2x4_ASAP7_75t_L g6596 ( 
.A(n_6387),
.B(n_120),
.Y(n_6596)
);

INVx1_ASAP7_75t_L g6597 ( 
.A(n_6441),
.Y(n_6597)
);

INVx2_ASAP7_75t_L g6598 ( 
.A(n_6436),
.Y(n_6598)
);

AND2x2_ASAP7_75t_L g6599 ( 
.A(n_6338),
.B(n_120),
.Y(n_6599)
);

INVx1_ASAP7_75t_L g6600 ( 
.A(n_6446),
.Y(n_6600)
);

INVx1_ASAP7_75t_L g6601 ( 
.A(n_6449),
.Y(n_6601)
);

INVx2_ASAP7_75t_L g6602 ( 
.A(n_6366),
.Y(n_6602)
);

NAND2xp5_ASAP7_75t_L g6603 ( 
.A(n_6433),
.B(n_120),
.Y(n_6603)
);

OR2x2_ASAP7_75t_L g6604 ( 
.A(n_6371),
.B(n_121),
.Y(n_6604)
);

HB1xp67_ASAP7_75t_L g6605 ( 
.A(n_6423),
.Y(n_6605)
);

AND2x4_ASAP7_75t_L g6606 ( 
.A(n_6426),
.B(n_6424),
.Y(n_6606)
);

AND2x2_ASAP7_75t_L g6607 ( 
.A(n_6353),
.B(n_121),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6472),
.Y(n_6608)
);

INVxp67_ASAP7_75t_SL g6609 ( 
.A(n_6455),
.Y(n_6609)
);

HB1xp67_ASAP7_75t_L g6610 ( 
.A(n_6389),
.Y(n_6610)
);

OR2x2_ASAP7_75t_L g6611 ( 
.A(n_6463),
.B(n_121),
.Y(n_6611)
);

AND2x2_ASAP7_75t_L g6612 ( 
.A(n_6357),
.B(n_121),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_6472),
.Y(n_6613)
);

HB1xp67_ASAP7_75t_L g6614 ( 
.A(n_6392),
.Y(n_6614)
);

INVx2_ASAP7_75t_L g6615 ( 
.A(n_6445),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_6464),
.B(n_122),
.Y(n_6616)
);

HB1xp67_ASAP7_75t_L g6617 ( 
.A(n_6460),
.Y(n_6617)
);

INVx1_ASAP7_75t_L g6618 ( 
.A(n_6452),
.Y(n_6618)
);

AO21x2_ASAP7_75t_L g6619 ( 
.A1(n_6383),
.A2(n_122),
.B(n_123),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_6493),
.Y(n_6620)
);

NAND4xp25_ASAP7_75t_L g6621 ( 
.A(n_6483),
.B(n_124),
.C(n_122),
.D(n_123),
.Y(n_6621)
);

INVx1_ASAP7_75t_L g6622 ( 
.A(n_6495),
.Y(n_6622)
);

INVx3_ASAP7_75t_L g6623 ( 
.A(n_6450),
.Y(n_6623)
);

NAND2xp5_ASAP7_75t_L g6624 ( 
.A(n_6368),
.B(n_122),
.Y(n_6624)
);

AND2x2_ASAP7_75t_L g6625 ( 
.A(n_6438),
.B(n_123),
.Y(n_6625)
);

INVx1_ASAP7_75t_L g6626 ( 
.A(n_6468),
.Y(n_6626)
);

INVx2_ASAP7_75t_L g6627 ( 
.A(n_6450),
.Y(n_6627)
);

OR2x2_ASAP7_75t_L g6628 ( 
.A(n_6453),
.B(n_123),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_6469),
.Y(n_6629)
);

INVx2_ASAP7_75t_L g6630 ( 
.A(n_6485),
.Y(n_6630)
);

AND2x2_ASAP7_75t_L g6631 ( 
.A(n_6442),
.B(n_124),
.Y(n_6631)
);

INVx1_ASAP7_75t_L g6632 ( 
.A(n_6466),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6473),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_6400),
.Y(n_6634)
);

HB1xp67_ASAP7_75t_L g6635 ( 
.A(n_6362),
.Y(n_6635)
);

INVx2_ASAP7_75t_L g6636 ( 
.A(n_6490),
.Y(n_6636)
);

INVx2_ASAP7_75t_L g6637 ( 
.A(n_6491),
.Y(n_6637)
);

HB1xp67_ASAP7_75t_L g6638 ( 
.A(n_6402),
.Y(n_6638)
);

BUFx6f_ASAP7_75t_L g6639 ( 
.A(n_6427),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_6404),
.Y(n_6640)
);

NAND2xp33_ASAP7_75t_SL g6641 ( 
.A(n_6456),
.B(n_124),
.Y(n_6641)
);

NAND2xp5_ASAP7_75t_L g6642 ( 
.A(n_6457),
.B(n_125),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6386),
.Y(n_6643)
);

INVx2_ASAP7_75t_L g6644 ( 
.A(n_6496),
.Y(n_6644)
);

HB1xp67_ASAP7_75t_L g6645 ( 
.A(n_6342),
.Y(n_6645)
);

HB1xp67_ASAP7_75t_L g6646 ( 
.A(n_6422),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6363),
.Y(n_6647)
);

INVx2_ASAP7_75t_L g6648 ( 
.A(n_6498),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6361),
.Y(n_6649)
);

INVx4_ASAP7_75t_L g6650 ( 
.A(n_6465),
.Y(n_6650)
);

BUFx3_ASAP7_75t_L g6651 ( 
.A(n_6477),
.Y(n_6651)
);

INVx1_ASAP7_75t_L g6652 ( 
.A(n_6421),
.Y(n_6652)
);

AOI221xp5_ASAP7_75t_L g6653 ( 
.A1(n_6430),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_128),
.Y(n_6653)
);

INVxp67_ASAP7_75t_L g6654 ( 
.A(n_6471),
.Y(n_6654)
);

INVx1_ASAP7_75t_L g6655 ( 
.A(n_6428),
.Y(n_6655)
);

AND2x2_ASAP7_75t_L g6656 ( 
.A(n_6487),
.B(n_126),
.Y(n_6656)
);

INVx3_ASAP7_75t_L g6657 ( 
.A(n_6500),
.Y(n_6657)
);

INVx1_ASAP7_75t_L g6658 ( 
.A(n_6412),
.Y(n_6658)
);

NOR2xp33_ASAP7_75t_L g6659 ( 
.A(n_6417),
.B(n_126),
.Y(n_6659)
);

OR2x2_ASAP7_75t_L g6660 ( 
.A(n_6354),
.B(n_6397),
.Y(n_6660)
);

INVx2_ASAP7_75t_L g6661 ( 
.A(n_6502),
.Y(n_6661)
);

INVx1_ASAP7_75t_L g6662 ( 
.A(n_6403),
.Y(n_6662)
);

OR2x2_ASAP7_75t_L g6663 ( 
.A(n_6415),
.B(n_127),
.Y(n_6663)
);

HB1xp67_ASAP7_75t_L g6664 ( 
.A(n_6431),
.Y(n_6664)
);

INVx2_ASAP7_75t_L g6665 ( 
.A(n_6454),
.Y(n_6665)
);

OAI221xp5_ASAP7_75t_SL g6666 ( 
.A1(n_6461),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.C(n_130),
.Y(n_6666)
);

INVx2_ASAP7_75t_L g6667 ( 
.A(n_6454),
.Y(n_6667)
);

INVxp67_ASAP7_75t_SL g6668 ( 
.A(n_6352),
.Y(n_6668)
);

AND2x2_ASAP7_75t_L g6669 ( 
.A(n_6458),
.B(n_128),
.Y(n_6669)
);

INVx2_ASAP7_75t_L g6670 ( 
.A(n_6476),
.Y(n_6670)
);

AND2x4_ASAP7_75t_L g6671 ( 
.A(n_6444),
.B(n_129),
.Y(n_6671)
);

INVx1_ASAP7_75t_L g6672 ( 
.A(n_6482),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6489),
.Y(n_6673)
);

INVx2_ASAP7_75t_L g6674 ( 
.A(n_6478),
.Y(n_6674)
);

INVx5_ASAP7_75t_L g6675 ( 
.A(n_6499),
.Y(n_6675)
);

INVx1_ASAP7_75t_L g6676 ( 
.A(n_6501),
.Y(n_6676)
);

INVx3_ASAP7_75t_L g6677 ( 
.A(n_6480),
.Y(n_6677)
);

NAND2xp5_ASAP7_75t_L g6678 ( 
.A(n_6384),
.B(n_129),
.Y(n_6678)
);

AND2x2_ASAP7_75t_L g6679 ( 
.A(n_6479),
.B(n_129),
.Y(n_6679)
);

BUFx2_ASAP7_75t_L g6680 ( 
.A(n_6486),
.Y(n_6680)
);

AND2x2_ASAP7_75t_L g6681 ( 
.A(n_6505),
.B(n_130),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_6406),
.Y(n_6682)
);

INVx4_ASAP7_75t_L g6683 ( 
.A(n_6467),
.Y(n_6683)
);

AND2x4_ASAP7_75t_L g6684 ( 
.A(n_6340),
.B(n_130),
.Y(n_6684)
);

AND2x2_ASAP7_75t_L g6685 ( 
.A(n_6364),
.B(n_130),
.Y(n_6685)
);

INVx1_ASAP7_75t_SL g6686 ( 
.A(n_6346),
.Y(n_6686)
);

OR2x2_ASAP7_75t_L g6687 ( 
.A(n_6341),
.B(n_131),
.Y(n_6687)
);

AND2x2_ASAP7_75t_L g6688 ( 
.A(n_6364),
.B(n_131),
.Y(n_6688)
);

OR2x2_ASAP7_75t_L g6689 ( 
.A(n_6341),
.B(n_131),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_6377),
.Y(n_6690)
);

BUFx2_ASAP7_75t_L g6691 ( 
.A(n_6409),
.Y(n_6691)
);

AND2x2_ASAP7_75t_L g6692 ( 
.A(n_6364),
.B(n_132),
.Y(n_6692)
);

INVx2_ASAP7_75t_L g6693 ( 
.A(n_6375),
.Y(n_6693)
);

NAND2xp5_ASAP7_75t_L g6694 ( 
.A(n_6375),
.B(n_132),
.Y(n_6694)
);

OR2x2_ASAP7_75t_L g6695 ( 
.A(n_6341),
.B(n_132),
.Y(n_6695)
);

AND2x4_ASAP7_75t_L g6696 ( 
.A(n_6333),
.B(n_132),
.Y(n_6696)
);

HB1xp67_ASAP7_75t_L g6697 ( 
.A(n_6377),
.Y(n_6697)
);

INVx2_ASAP7_75t_L g6698 ( 
.A(n_6375),
.Y(n_6698)
);

AND2x2_ASAP7_75t_L g6699 ( 
.A(n_6364),
.B(n_133),
.Y(n_6699)
);

NAND3xp33_ASAP7_75t_SL g6700 ( 
.A(n_6375),
.B(n_133),
.C(n_134),
.Y(n_6700)
);

AOI22xp33_ASAP7_75t_L g6701 ( 
.A1(n_6376),
.A2(n_765),
.B1(n_766),
.B2(n_764),
.Y(n_6701)
);

INVx2_ASAP7_75t_SL g6702 ( 
.A(n_6346),
.Y(n_6702)
);

BUFx6f_ASAP7_75t_L g6703 ( 
.A(n_6346),
.Y(n_6703)
);

AND2x2_ASAP7_75t_L g6704 ( 
.A(n_6364),
.B(n_133),
.Y(n_6704)
);

BUFx6f_ASAP7_75t_L g6705 ( 
.A(n_6346),
.Y(n_6705)
);

AOI22xp33_ASAP7_75t_SL g6706 ( 
.A1(n_6376),
.A2(n_766),
.B1(n_767),
.B2(n_765),
.Y(n_6706)
);

AND2x4_ASAP7_75t_L g6707 ( 
.A(n_6364),
.B(n_133),
.Y(n_6707)
);

NOR2x1_ASAP7_75t_L g6708 ( 
.A(n_6364),
.B(n_134),
.Y(n_6708)
);

AOI22xp33_ASAP7_75t_L g6709 ( 
.A1(n_6376),
.A2(n_767),
.B1(n_768),
.B2(n_766),
.Y(n_6709)
);

INVxp67_ASAP7_75t_L g6710 ( 
.A(n_6343),
.Y(n_6710)
);

INVx1_ASAP7_75t_L g6711 ( 
.A(n_6377),
.Y(n_6711)
);

NAND2xp5_ASAP7_75t_L g6712 ( 
.A(n_6375),
.B(n_134),
.Y(n_6712)
);

INVx2_ASAP7_75t_L g6713 ( 
.A(n_6375),
.Y(n_6713)
);

INVx2_ASAP7_75t_L g6714 ( 
.A(n_6375),
.Y(n_6714)
);

AOI22xp5_ASAP7_75t_L g6715 ( 
.A1(n_6503),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.Y(n_6715)
);

OR2x2_ASAP7_75t_L g6716 ( 
.A(n_6341),
.B(n_135),
.Y(n_6716)
);

INVx1_ASAP7_75t_L g6717 ( 
.A(n_6377),
.Y(n_6717)
);

INVx2_ASAP7_75t_L g6718 ( 
.A(n_6520),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_6685),
.Y(n_6719)
);

INVx1_ASAP7_75t_L g6720 ( 
.A(n_6688),
.Y(n_6720)
);

OR2x2_ASAP7_75t_L g6721 ( 
.A(n_6506),
.B(n_135),
.Y(n_6721)
);

NAND2xp5_ASAP7_75t_L g6722 ( 
.A(n_6693),
.B(n_136),
.Y(n_6722)
);

AND2x2_ASAP7_75t_L g6723 ( 
.A(n_6513),
.B(n_137),
.Y(n_6723)
);

NAND2xp5_ASAP7_75t_L g6724 ( 
.A(n_6698),
.B(n_137),
.Y(n_6724)
);

INVx2_ASAP7_75t_L g6725 ( 
.A(n_6703),
.Y(n_6725)
);

INVx1_ASAP7_75t_L g6726 ( 
.A(n_6692),
.Y(n_6726)
);

AND2x2_ASAP7_75t_L g6727 ( 
.A(n_6513),
.B(n_137),
.Y(n_6727)
);

HB1xp67_ASAP7_75t_L g6728 ( 
.A(n_6713),
.Y(n_6728)
);

HB1xp67_ASAP7_75t_L g6729 ( 
.A(n_6714),
.Y(n_6729)
);

AND2x2_ASAP7_75t_L g6730 ( 
.A(n_6686),
.B(n_138),
.Y(n_6730)
);

AND2x4_ASAP7_75t_L g6731 ( 
.A(n_6508),
.B(n_138),
.Y(n_6731)
);

AND2x2_ASAP7_75t_L g6732 ( 
.A(n_6703),
.B(n_138),
.Y(n_6732)
);

NOR2xp67_ASAP7_75t_L g6733 ( 
.A(n_6702),
.B(n_139),
.Y(n_6733)
);

AND2x2_ASAP7_75t_L g6734 ( 
.A(n_6705),
.B(n_139),
.Y(n_6734)
);

AND2x2_ASAP7_75t_L g6735 ( 
.A(n_6705),
.B(n_139),
.Y(n_6735)
);

AND2x2_ASAP7_75t_L g6736 ( 
.A(n_6562),
.B(n_139),
.Y(n_6736)
);

AND2x4_ASAP7_75t_L g6737 ( 
.A(n_6551),
.B(n_140),
.Y(n_6737)
);

AND2x2_ASAP7_75t_L g6738 ( 
.A(n_6514),
.B(n_140),
.Y(n_6738)
);

INVx2_ASAP7_75t_SL g6739 ( 
.A(n_6519),
.Y(n_6739)
);

NOR2x1_ASAP7_75t_L g6740 ( 
.A(n_6516),
.B(n_140),
.Y(n_6740)
);

INVx2_ASAP7_75t_L g6741 ( 
.A(n_6516),
.Y(n_6741)
);

AND2x2_ASAP7_75t_L g6742 ( 
.A(n_6547),
.B(n_141),
.Y(n_6742)
);

NAND2xp5_ASAP7_75t_L g6743 ( 
.A(n_6512),
.B(n_141),
.Y(n_6743)
);

NAND2xp5_ASAP7_75t_L g6744 ( 
.A(n_6512),
.B(n_6587),
.Y(n_6744)
);

AND2x4_ASAP7_75t_L g6745 ( 
.A(n_6691),
.B(n_141),
.Y(n_6745)
);

NAND2xp5_ASAP7_75t_L g6746 ( 
.A(n_6535),
.B(n_142),
.Y(n_6746)
);

INVx1_ASAP7_75t_L g6747 ( 
.A(n_6699),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_6704),
.Y(n_6748)
);

INVx1_ASAP7_75t_L g6749 ( 
.A(n_6590),
.Y(n_6749)
);

HB1xp67_ASAP7_75t_L g6750 ( 
.A(n_6541),
.Y(n_6750)
);

AND2x2_ASAP7_75t_L g6751 ( 
.A(n_6691),
.B(n_142),
.Y(n_6751)
);

NAND2x1p5_ASAP7_75t_L g6752 ( 
.A(n_6707),
.B(n_142),
.Y(n_6752)
);

AND2x2_ASAP7_75t_L g6753 ( 
.A(n_6570),
.B(n_142),
.Y(n_6753)
);

INVx1_ASAP7_75t_L g6754 ( 
.A(n_6590),
.Y(n_6754)
);

NAND2xp5_ASAP7_75t_L g6755 ( 
.A(n_6560),
.B(n_143),
.Y(n_6755)
);

OR2x2_ASAP7_75t_L g6756 ( 
.A(n_6658),
.B(n_143),
.Y(n_6756)
);

AND2x2_ASAP7_75t_L g6757 ( 
.A(n_6573),
.B(n_143),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6694),
.Y(n_6758)
);

NAND2xp5_ASAP7_75t_L g6759 ( 
.A(n_6589),
.B(n_143),
.Y(n_6759)
);

AND2x2_ASAP7_75t_L g6760 ( 
.A(n_6567),
.B(n_144),
.Y(n_6760)
);

OR2x2_ASAP7_75t_L g6761 ( 
.A(n_6555),
.B(n_145),
.Y(n_6761)
);

NAND2xp5_ASAP7_75t_L g6762 ( 
.A(n_6682),
.B(n_145),
.Y(n_6762)
);

OR2x2_ASAP7_75t_L g6763 ( 
.A(n_6531),
.B(n_145),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_6712),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6696),
.Y(n_6765)
);

AND2x2_ASAP7_75t_L g6766 ( 
.A(n_6567),
.B(n_145),
.Y(n_6766)
);

AND2x2_ASAP7_75t_L g6767 ( 
.A(n_6565),
.B(n_146),
.Y(n_6767)
);

NAND2xp5_ASAP7_75t_L g6768 ( 
.A(n_6675),
.B(n_146),
.Y(n_6768)
);

AND2x4_ASAP7_75t_L g6769 ( 
.A(n_6627),
.B(n_146),
.Y(n_6769)
);

NOR2x1_ASAP7_75t_L g6770 ( 
.A(n_6568),
.B(n_146),
.Y(n_6770)
);

INVx2_ASAP7_75t_SL g6771 ( 
.A(n_6556),
.Y(n_6771)
);

INVx1_ASAP7_75t_L g6772 ( 
.A(n_6563),
.Y(n_6772)
);

AND2x2_ASAP7_75t_L g6773 ( 
.A(n_6565),
.B(n_147),
.Y(n_6773)
);

NAND2xp5_ASAP7_75t_SL g6774 ( 
.A(n_6675),
.B(n_147),
.Y(n_6774)
);

AND2x2_ASAP7_75t_L g6775 ( 
.A(n_6543),
.B(n_147),
.Y(n_6775)
);

AND2x2_ASAP7_75t_L g6776 ( 
.A(n_6527),
.B(n_147),
.Y(n_6776)
);

AND2x2_ASAP7_75t_L g6777 ( 
.A(n_6530),
.B(n_148),
.Y(n_6777)
);

INVx1_ASAP7_75t_L g6778 ( 
.A(n_6574),
.Y(n_6778)
);

AND2x2_ASAP7_75t_L g6779 ( 
.A(n_6675),
.B(n_148),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_6707),
.Y(n_6780)
);

AND2x2_ASAP7_75t_L g6781 ( 
.A(n_6680),
.B(n_148),
.Y(n_6781)
);

NAND2xp5_ASAP7_75t_SL g6782 ( 
.A(n_6654),
.B(n_148),
.Y(n_6782)
);

INVx2_ASAP7_75t_L g6783 ( 
.A(n_6581),
.Y(n_6783)
);

NAND2xp5_ASAP7_75t_L g6784 ( 
.A(n_6539),
.B(n_6650),
.Y(n_6784)
);

OR2x2_ASAP7_75t_L g6785 ( 
.A(n_6534),
.B(n_149),
.Y(n_6785)
);

AND2x2_ASAP7_75t_L g6786 ( 
.A(n_6680),
.B(n_6524),
.Y(n_6786)
);

BUFx2_ASAP7_75t_L g6787 ( 
.A(n_6544),
.Y(n_6787)
);

NAND2x1p5_ASAP7_75t_L g6788 ( 
.A(n_6671),
.B(n_149),
.Y(n_6788)
);

AND2x2_ASAP7_75t_L g6789 ( 
.A(n_6517),
.B(n_149),
.Y(n_6789)
);

NAND2xp5_ASAP7_75t_SL g6790 ( 
.A(n_6568),
.B(n_150),
.Y(n_6790)
);

OR2x2_ASAP7_75t_L g6791 ( 
.A(n_6540),
.B(n_150),
.Y(n_6791)
);

NAND2xp5_ASAP7_75t_L g6792 ( 
.A(n_6585),
.B(n_150),
.Y(n_6792)
);

AND2x2_ASAP7_75t_L g6793 ( 
.A(n_6578),
.B(n_151),
.Y(n_6793)
);

INVx1_ASAP7_75t_L g6794 ( 
.A(n_6558),
.Y(n_6794)
);

AND2x4_ASAP7_75t_L g6795 ( 
.A(n_6583),
.B(n_151),
.Y(n_6795)
);

INVx1_ASAP7_75t_L g6796 ( 
.A(n_6561),
.Y(n_6796)
);

INVx1_ASAP7_75t_L g6797 ( 
.A(n_6564),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6559),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_6576),
.Y(n_6799)
);

NAND2xp5_ASAP7_75t_L g6800 ( 
.A(n_6659),
.B(n_151),
.Y(n_6800)
);

INVx1_ASAP7_75t_L g6801 ( 
.A(n_6584),
.Y(n_6801)
);

AND2x4_ASAP7_75t_SL g6802 ( 
.A(n_6665),
.B(n_152),
.Y(n_6802)
);

OR2x2_ASAP7_75t_L g6803 ( 
.A(n_6603),
.B(n_152),
.Y(n_6803)
);

INVx1_ASAP7_75t_L g6804 ( 
.A(n_6586),
.Y(n_6804)
);

HB1xp67_ASAP7_75t_L g6805 ( 
.A(n_6597),
.Y(n_6805)
);

AND2x2_ASAP7_75t_L g6806 ( 
.A(n_6532),
.B(n_6550),
.Y(n_6806)
);

INVx1_ASAP7_75t_L g6807 ( 
.A(n_6600),
.Y(n_6807)
);

AND2x2_ASAP7_75t_L g6808 ( 
.A(n_6509),
.B(n_152),
.Y(n_6808)
);

AND2x2_ASAP7_75t_L g6809 ( 
.A(n_6697),
.B(n_152),
.Y(n_6809)
);

NAND2xp5_ASAP7_75t_L g6810 ( 
.A(n_6671),
.B(n_153),
.Y(n_6810)
);

HB1xp67_ASAP7_75t_L g6811 ( 
.A(n_6601),
.Y(n_6811)
);

AND2x4_ASAP7_75t_L g6812 ( 
.A(n_6623),
.B(n_153),
.Y(n_6812)
);

INVx2_ASAP7_75t_L g6813 ( 
.A(n_6571),
.Y(n_6813)
);

NAND2xp5_ASAP7_75t_L g6814 ( 
.A(n_6708),
.B(n_153),
.Y(n_6814)
);

INVx1_ASAP7_75t_L g6815 ( 
.A(n_6593),
.Y(n_6815)
);

OR2x2_ASAP7_75t_L g6816 ( 
.A(n_6624),
.B(n_154),
.Y(n_6816)
);

INVx2_ASAP7_75t_L g6817 ( 
.A(n_6575),
.Y(n_6817)
);

INVxp67_ASAP7_75t_SL g6818 ( 
.A(n_6592),
.Y(n_6818)
);

INVx1_ASAP7_75t_L g6819 ( 
.A(n_6593),
.Y(n_6819)
);

AND2x2_ASAP7_75t_L g6820 ( 
.A(n_6599),
.B(n_154),
.Y(n_6820)
);

INVx1_ASAP7_75t_L g6821 ( 
.A(n_6617),
.Y(n_6821)
);

INVxp67_ASAP7_75t_L g6822 ( 
.A(n_6641),
.Y(n_6822)
);

INVx1_ASAP7_75t_L g6823 ( 
.A(n_6579),
.Y(n_6823)
);

NAND2xp5_ASAP7_75t_L g6824 ( 
.A(n_6684),
.B(n_155),
.Y(n_6824)
);

AND2x2_ASAP7_75t_L g6825 ( 
.A(n_6607),
.B(n_155),
.Y(n_6825)
);

NAND2xp5_ASAP7_75t_SL g6826 ( 
.A(n_6566),
.B(n_155),
.Y(n_6826)
);

AND2x2_ASAP7_75t_L g6827 ( 
.A(n_6651),
.B(n_155),
.Y(n_6827)
);

INVx2_ASAP7_75t_L g6828 ( 
.A(n_6595),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_6598),
.Y(n_6829)
);

INVx1_ASAP7_75t_L g6830 ( 
.A(n_6610),
.Y(n_6830)
);

INVx1_ASAP7_75t_L g6831 ( 
.A(n_6614),
.Y(n_6831)
);

NAND2xp5_ASAP7_75t_L g6832 ( 
.A(n_6684),
.B(n_156),
.Y(n_6832)
);

HB1xp67_ASAP7_75t_L g6833 ( 
.A(n_6582),
.Y(n_6833)
);

NOR2x1p5_ASAP7_75t_L g6834 ( 
.A(n_6609),
.B(n_156),
.Y(n_6834)
);

OR2x2_ASAP7_75t_L g6835 ( 
.A(n_6553),
.B(n_156),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_6569),
.Y(n_6836)
);

INVx1_ASAP7_75t_L g6837 ( 
.A(n_6646),
.Y(n_6837)
);

INVx1_ASAP7_75t_L g6838 ( 
.A(n_6667),
.Y(n_6838)
);

OR2x2_ASAP7_75t_L g6839 ( 
.A(n_6507),
.B(n_156),
.Y(n_6839)
);

INVx1_ASAP7_75t_L g6840 ( 
.A(n_6638),
.Y(n_6840)
);

INVx1_ASAP7_75t_L g6841 ( 
.A(n_6615),
.Y(n_6841)
);

AND2x2_ASAP7_75t_L g6842 ( 
.A(n_6548),
.B(n_157),
.Y(n_6842)
);

NAND2xp5_ASAP7_75t_L g6843 ( 
.A(n_6677),
.B(n_157),
.Y(n_6843)
);

NAND2xp5_ASAP7_75t_L g6844 ( 
.A(n_6510),
.B(n_157),
.Y(n_6844)
);

INVx2_ASAP7_75t_L g6845 ( 
.A(n_6518),
.Y(n_6845)
);

AND2x2_ASAP7_75t_L g6846 ( 
.A(n_6612),
.B(n_157),
.Y(n_6846)
);

OR2x2_ASAP7_75t_L g6847 ( 
.A(n_6690),
.B(n_158),
.Y(n_6847)
);

OR2x2_ASAP7_75t_L g6848 ( 
.A(n_6711),
.B(n_158),
.Y(n_6848)
);

BUFx2_ASAP7_75t_L g6849 ( 
.A(n_6606),
.Y(n_6849)
);

INVx1_ASAP7_75t_L g6850 ( 
.A(n_6525),
.Y(n_6850)
);

INVxp67_ASAP7_75t_L g6851 ( 
.A(n_6625),
.Y(n_6851)
);

BUFx2_ASAP7_75t_L g6852 ( 
.A(n_6533),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6608),
.Y(n_6853)
);

NAND2xp5_ASAP7_75t_L g6854 ( 
.A(n_6554),
.B(n_159),
.Y(n_6854)
);

AND2x4_ASAP7_75t_SL g6855 ( 
.A(n_6683),
.B(n_159),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_6613),
.Y(n_6856)
);

INVx1_ASAP7_75t_L g6857 ( 
.A(n_6549),
.Y(n_6857)
);

NAND2xp5_ASAP7_75t_SL g6858 ( 
.A(n_6552),
.B(n_159),
.Y(n_6858)
);

OR2x2_ASAP7_75t_L g6859 ( 
.A(n_6717),
.B(n_159),
.Y(n_6859)
);

AND2x2_ASAP7_75t_L g6860 ( 
.A(n_6656),
.B(n_160),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6591),
.B(n_160),
.Y(n_6861)
);

AND2x2_ASAP7_75t_L g6862 ( 
.A(n_6647),
.B(n_160),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6632),
.Y(n_6863)
);

INVx1_ASAP7_75t_L g6864 ( 
.A(n_6633),
.Y(n_6864)
);

NAND2xp5_ASAP7_75t_L g6865 ( 
.A(n_6542),
.B(n_160),
.Y(n_6865)
);

INVx2_ASAP7_75t_L g6866 ( 
.A(n_6657),
.Y(n_6866)
);

AND2x4_ASAP7_75t_L g6867 ( 
.A(n_6537),
.B(n_161),
.Y(n_6867)
);

INVxp67_ASAP7_75t_SL g6868 ( 
.A(n_6611),
.Y(n_6868)
);

INVx1_ASAP7_75t_L g6869 ( 
.A(n_6681),
.Y(n_6869)
);

AND2x2_ASAP7_75t_L g6870 ( 
.A(n_6538),
.B(n_161),
.Y(n_6870)
);

INVx2_ASAP7_75t_L g6871 ( 
.A(n_6630),
.Y(n_6871)
);

AND2x2_ASAP7_75t_L g6872 ( 
.A(n_6511),
.B(n_161),
.Y(n_6872)
);

NAND2xp5_ASAP7_75t_L g6873 ( 
.A(n_6706),
.B(n_162),
.Y(n_6873)
);

AND2x4_ASAP7_75t_SL g6874 ( 
.A(n_6596),
.B(n_162),
.Y(n_6874)
);

AND2x2_ASAP7_75t_L g6875 ( 
.A(n_6618),
.B(n_162),
.Y(n_6875)
);

INVx2_ASAP7_75t_L g6876 ( 
.A(n_6636),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_6515),
.B(n_162),
.Y(n_6877)
);

NAND2xp5_ASAP7_75t_L g6878 ( 
.A(n_6521),
.B(n_163),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6557),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_6631),
.Y(n_6880)
);

NAND2xp5_ASAP7_75t_L g6881 ( 
.A(n_6652),
.B(n_163),
.Y(n_6881)
);

OAI221xp5_ASAP7_75t_SL g6882 ( 
.A1(n_6634),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.C(n_166),
.Y(n_6882)
);

OR2x2_ASAP7_75t_L g6883 ( 
.A(n_6580),
.B(n_164),
.Y(n_6883)
);

AND2x4_ASAP7_75t_L g6884 ( 
.A(n_6718),
.B(n_6725),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6806),
.B(n_6536),
.Y(n_6885)
);

INVx1_ASAP7_75t_L g6886 ( 
.A(n_6723),
.Y(n_6886)
);

NOR2xp33_ASAP7_75t_L g6887 ( 
.A(n_6741),
.B(n_6710),
.Y(n_6887)
);

INVx1_ASAP7_75t_L g6888 ( 
.A(n_6727),
.Y(n_6888)
);

NAND2xp5_ASAP7_75t_L g6889 ( 
.A(n_6736),
.B(n_6701),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6767),
.Y(n_6890)
);

INVx2_ASAP7_75t_SL g6891 ( 
.A(n_6737),
.Y(n_6891)
);

INVx1_ASAP7_75t_L g6892 ( 
.A(n_6773),
.Y(n_6892)
);

INVx1_ASAP7_75t_L g6893 ( 
.A(n_6751),
.Y(n_6893)
);

NOR2xp33_ASAP7_75t_L g6894 ( 
.A(n_6822),
.B(n_6626),
.Y(n_6894)
);

AND2x2_ASAP7_75t_L g6895 ( 
.A(n_6786),
.B(n_6629),
.Y(n_6895)
);

INVx1_ASAP7_75t_L g6896 ( 
.A(n_6753),
.Y(n_6896)
);

INVx1_ASAP7_75t_L g6897 ( 
.A(n_6730),
.Y(n_6897)
);

OR2x2_ASAP7_75t_L g6898 ( 
.A(n_6759),
.B(n_6523),
.Y(n_6898)
);

AND2x2_ASAP7_75t_L g6899 ( 
.A(n_6789),
.B(n_6672),
.Y(n_6899)
);

OR2x2_ASAP7_75t_L g6900 ( 
.A(n_6761),
.B(n_6743),
.Y(n_6900)
);

NAND2xp5_ASAP7_75t_L g6901 ( 
.A(n_6795),
.B(n_6709),
.Y(n_6901)
);

AND2x2_ASAP7_75t_L g6902 ( 
.A(n_6742),
.B(n_6776),
.Y(n_6902)
);

NAND2xp5_ASAP7_75t_L g6903 ( 
.A(n_6795),
.B(n_6715),
.Y(n_6903)
);

NAND2xp5_ASAP7_75t_L g6904 ( 
.A(n_6731),
.B(n_6655),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6833),
.Y(n_6905)
);

NAND2xp67_ASAP7_75t_L g6906 ( 
.A(n_6855),
.B(n_6674),
.Y(n_6906)
);

AND2x2_ASAP7_75t_L g6907 ( 
.A(n_6777),
.B(n_6673),
.Y(n_6907)
);

INVx1_ASAP7_75t_L g6908 ( 
.A(n_6728),
.Y(n_6908)
);

INVx1_ASAP7_75t_L g6909 ( 
.A(n_6729),
.Y(n_6909)
);

BUFx3_ASAP7_75t_L g6910 ( 
.A(n_6737),
.Y(n_6910)
);

AND2x2_ASAP7_75t_L g6911 ( 
.A(n_6870),
.B(n_6775),
.Y(n_6911)
);

AND2x2_ASAP7_75t_L g6912 ( 
.A(n_6842),
.B(n_6676),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_6731),
.Y(n_6913)
);

OR2x2_ASAP7_75t_L g6914 ( 
.A(n_6768),
.B(n_6588),
.Y(n_6914)
);

BUFx3_ASAP7_75t_L g6915 ( 
.A(n_6732),
.Y(n_6915)
);

OR2x2_ASAP7_75t_L g6916 ( 
.A(n_6762),
.B(n_6526),
.Y(n_6916)
);

OR2x2_ASAP7_75t_L g6917 ( 
.A(n_6803),
.B(n_6522),
.Y(n_6917)
);

AND2x2_ASAP7_75t_L g6918 ( 
.A(n_6861),
.B(n_6760),
.Y(n_6918)
);

INVx1_ASAP7_75t_L g6919 ( 
.A(n_6766),
.Y(n_6919)
);

INVx2_ASAP7_75t_L g6920 ( 
.A(n_6783),
.Y(n_6920)
);

OR2x2_ASAP7_75t_L g6921 ( 
.A(n_6746),
.B(n_6528),
.Y(n_6921)
);

INVx2_ASAP7_75t_L g6922 ( 
.A(n_6734),
.Y(n_6922)
);

HB1xp67_ASAP7_75t_L g6923 ( 
.A(n_6745),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_6779),
.Y(n_6924)
);

NAND3xp33_ASAP7_75t_L g6925 ( 
.A(n_6854),
.B(n_6643),
.C(n_6653),
.Y(n_6925)
);

AND2x2_ASAP7_75t_L g6926 ( 
.A(n_6827),
.B(n_6529),
.Y(n_6926)
);

AND2x2_ASAP7_75t_L g6927 ( 
.A(n_6849),
.B(n_6577),
.Y(n_6927)
);

NAND2xp5_ASAP7_75t_L g6928 ( 
.A(n_6745),
.B(n_6668),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_L g6929 ( 
.A(n_6769),
.B(n_6670),
.Y(n_6929)
);

AND2x2_ASAP7_75t_L g6930 ( 
.A(n_6739),
.B(n_6572),
.Y(n_6930)
);

OR2x2_ASAP7_75t_L g6931 ( 
.A(n_6816),
.B(n_6771),
.Y(n_6931)
);

INVx2_ASAP7_75t_L g6932 ( 
.A(n_6735),
.Y(n_6932)
);

OR2x2_ASAP7_75t_L g6933 ( 
.A(n_6814),
.B(n_6616),
.Y(n_6933)
);

HB1xp67_ASAP7_75t_L g6934 ( 
.A(n_6812),
.Y(n_6934)
);

NAND2xp5_ASAP7_75t_L g6935 ( 
.A(n_6769),
.B(n_6781),
.Y(n_6935)
);

NOR2xp33_ASAP7_75t_L g6936 ( 
.A(n_6774),
.B(n_6744),
.Y(n_6936)
);

AND2x2_ASAP7_75t_L g6937 ( 
.A(n_6738),
.B(n_6546),
.Y(n_6937)
);

NOR2xp33_ASAP7_75t_L g6938 ( 
.A(n_6765),
.B(n_6545),
.Y(n_6938)
);

INVx1_ASAP7_75t_L g6939 ( 
.A(n_6812),
.Y(n_6939)
);

INVx1_ASAP7_75t_L g6940 ( 
.A(n_6810),
.Y(n_6940)
);

INVx1_ASAP7_75t_SL g6941 ( 
.A(n_6802),
.Y(n_6941)
);

INVx1_ASAP7_75t_L g6942 ( 
.A(n_6788),
.Y(n_6942)
);

INVx2_ASAP7_75t_L g6943 ( 
.A(n_6836),
.Y(n_6943)
);

NOR2x1_ASAP7_75t_L g6944 ( 
.A(n_6740),
.B(n_6619),
.Y(n_6944)
);

NAND2xp5_ASAP7_75t_L g6945 ( 
.A(n_6733),
.B(n_6620),
.Y(n_6945)
);

AND2x2_ASAP7_75t_L g6946 ( 
.A(n_6757),
.B(n_6662),
.Y(n_6946)
);

INVxp67_ASAP7_75t_L g6947 ( 
.A(n_6793),
.Y(n_6947)
);

AND2x2_ASAP7_75t_L g6948 ( 
.A(n_6862),
.B(n_6594),
.Y(n_6948)
);

AND2x2_ASAP7_75t_L g6949 ( 
.A(n_6875),
.B(n_6669),
.Y(n_6949)
);

NOR2xp33_ASAP7_75t_L g6950 ( 
.A(n_6869),
.B(n_6749),
.Y(n_6950)
);

NOR2xp33_ASAP7_75t_L g6951 ( 
.A(n_6754),
.B(n_6639),
.Y(n_6951)
);

AND2x4_ASAP7_75t_L g6952 ( 
.A(n_6845),
.B(n_6640),
.Y(n_6952)
);

INVx2_ASAP7_75t_L g6953 ( 
.A(n_6813),
.Y(n_6953)
);

AND2x2_ASAP7_75t_L g6954 ( 
.A(n_6808),
.B(n_6679),
.Y(n_6954)
);

AND2x2_ASAP7_75t_L g6955 ( 
.A(n_6809),
.B(n_6649),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_6852),
.Y(n_6956)
);

AND2x2_ASAP7_75t_L g6957 ( 
.A(n_6872),
.B(n_6622),
.Y(n_6957)
);

AND2x2_ASAP7_75t_L g6958 ( 
.A(n_6877),
.B(n_6639),
.Y(n_6958)
);

OR2x2_ASAP7_75t_L g6959 ( 
.A(n_6791),
.B(n_6642),
.Y(n_6959)
);

NAND2xp5_ASAP7_75t_L g6960 ( 
.A(n_6867),
.B(n_6605),
.Y(n_6960)
);

HB1xp67_ASAP7_75t_L g6961 ( 
.A(n_6772),
.Y(n_6961)
);

INVx1_ASAP7_75t_L g6962 ( 
.A(n_6722),
.Y(n_6962)
);

NAND2xp5_ASAP7_75t_L g6963 ( 
.A(n_6867),
.B(n_6637),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_6780),
.B(n_6660),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6724),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6752),
.Y(n_6966)
);

NAND4xp25_ASAP7_75t_L g6967 ( 
.A(n_6784),
.B(n_6700),
.C(n_6621),
.D(n_6666),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6820),
.B(n_6644),
.Y(n_6968)
);

AND2x2_ASAP7_75t_L g6969 ( 
.A(n_6825),
.B(n_6648),
.Y(n_6969)
);

AOI22xp33_ASAP7_75t_L g6970 ( 
.A1(n_6866),
.A2(n_6661),
.B1(n_6635),
.B2(n_6602),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_6721),
.Y(n_6971)
);

BUFx2_ASAP7_75t_L g6972 ( 
.A(n_6817),
.Y(n_6972)
);

AND2x2_ASAP7_75t_L g6973 ( 
.A(n_6846),
.B(n_6628),
.Y(n_6973)
);

INVx1_ASAP7_75t_L g6974 ( 
.A(n_6843),
.Y(n_6974)
);

NAND2xp5_ASAP7_75t_L g6975 ( 
.A(n_6860),
.B(n_6645),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_6851),
.B(n_6663),
.Y(n_6976)
);

INVx1_ASAP7_75t_L g6977 ( 
.A(n_6824),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6832),
.Y(n_6978)
);

NOR2xp33_ASAP7_75t_L g6979 ( 
.A(n_6790),
.B(n_6828),
.Y(n_6979)
);

NAND2xp5_ASAP7_75t_L g6980 ( 
.A(n_6770),
.B(n_6664),
.Y(n_6980)
);

AND2x2_ASAP7_75t_L g6981 ( 
.A(n_6868),
.B(n_6687),
.Y(n_6981)
);

INVx3_ASAP7_75t_L g6982 ( 
.A(n_6871),
.Y(n_6982)
);

AND2x2_ASAP7_75t_L g6983 ( 
.A(n_6815),
.B(n_6689),
.Y(n_6983)
);

NAND2xp5_ASAP7_75t_L g6984 ( 
.A(n_6823),
.B(n_6678),
.Y(n_6984)
);

AND2x2_ASAP7_75t_L g6985 ( 
.A(n_6819),
.B(n_6695),
.Y(n_6985)
);

BUFx2_ASAP7_75t_L g6986 ( 
.A(n_6829),
.Y(n_6986)
);

NAND2xp5_ASAP7_75t_L g6987 ( 
.A(n_6838),
.B(n_6716),
.Y(n_6987)
);

NAND2xp5_ASAP7_75t_L g6988 ( 
.A(n_6799),
.B(n_6604),
.Y(n_6988)
);

AND3x2_ASAP7_75t_L g6989 ( 
.A(n_6787),
.B(n_164),
.C(n_165),
.Y(n_6989)
);

AND2x2_ASAP7_75t_L g6990 ( 
.A(n_6880),
.B(n_164),
.Y(n_6990)
);

OR2x2_ASAP7_75t_L g6991 ( 
.A(n_6763),
.B(n_166),
.Y(n_6991)
);

INVx1_ASAP7_75t_L g6992 ( 
.A(n_6750),
.Y(n_6992)
);

INVx2_ASAP7_75t_L g6993 ( 
.A(n_6876),
.Y(n_6993)
);

NAND2xp5_ASAP7_75t_L g6994 ( 
.A(n_6797),
.B(n_166),
.Y(n_6994)
);

INVx1_ASAP7_75t_L g6995 ( 
.A(n_6805),
.Y(n_6995)
);

OR2x2_ASAP7_75t_L g6996 ( 
.A(n_6785),
.B(n_6756),
.Y(n_6996)
);

NAND2x1_ASAP7_75t_L g6997 ( 
.A(n_6841),
.B(n_166),
.Y(n_6997)
);

INVx1_ASAP7_75t_L g6998 ( 
.A(n_6811),
.Y(n_6998)
);

AND2x2_ASAP7_75t_L g6999 ( 
.A(n_6778),
.B(n_167),
.Y(n_6999)
);

NAND2xp5_ASAP7_75t_L g7000 ( 
.A(n_6719),
.B(n_167),
.Y(n_7000)
);

NAND2xp5_ASAP7_75t_L g7001 ( 
.A(n_6720),
.B(n_6726),
.Y(n_7001)
);

HB1xp67_ASAP7_75t_L g7002 ( 
.A(n_6837),
.Y(n_7002)
);

INVx1_ASAP7_75t_L g7003 ( 
.A(n_6844),
.Y(n_7003)
);

AND2x2_ASAP7_75t_L g7004 ( 
.A(n_6834),
.B(n_167),
.Y(n_7004)
);

AOI21xp33_ASAP7_75t_SL g7005 ( 
.A1(n_6858),
.A2(n_167),
.B(n_168),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6747),
.B(n_168),
.Y(n_7006)
);

AND2x2_ASAP7_75t_L g7007 ( 
.A(n_6748),
.B(n_6850),
.Y(n_7007)
);

INVx4_ASAP7_75t_L g7008 ( 
.A(n_6874),
.Y(n_7008)
);

OAI22xp5_ASAP7_75t_L g7009 ( 
.A1(n_6835),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6865),
.Y(n_7010)
);

AND2x2_ASAP7_75t_L g7011 ( 
.A(n_6818),
.B(n_168),
.Y(n_7011)
);

AND2x2_ASAP7_75t_L g7012 ( 
.A(n_6758),
.B(n_169),
.Y(n_7012)
);

INVx3_ASAP7_75t_L g7013 ( 
.A(n_6798),
.Y(n_7013)
);

OR2x2_ASAP7_75t_L g7014 ( 
.A(n_6800),
.B(n_169),
.Y(n_7014)
);

INVx1_ASAP7_75t_L g7015 ( 
.A(n_6792),
.Y(n_7015)
);

INVx2_ASAP7_75t_L g7016 ( 
.A(n_6830),
.Y(n_7016)
);

AND2x2_ASAP7_75t_L g7017 ( 
.A(n_6764),
.B(n_170),
.Y(n_7017)
);

NAND2xp5_ASAP7_75t_L g7018 ( 
.A(n_6831),
.B(n_170),
.Y(n_7018)
);

OR2x2_ASAP7_75t_L g7019 ( 
.A(n_6847),
.B(n_170),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6755),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6848),
.Y(n_7021)
);

OR2x2_ASAP7_75t_L g7022 ( 
.A(n_6859),
.B(n_171),
.Y(n_7022)
);

AND2x2_ASAP7_75t_L g7023 ( 
.A(n_6801),
.B(n_171),
.Y(n_7023)
);

OR2x2_ASAP7_75t_L g7024 ( 
.A(n_6839),
.B(n_171),
.Y(n_7024)
);

INVx1_ASAP7_75t_SL g7025 ( 
.A(n_6821),
.Y(n_7025)
);

INVx2_ASAP7_75t_L g7026 ( 
.A(n_6840),
.Y(n_7026)
);

NAND2xp5_ASAP7_75t_L g7027 ( 
.A(n_6873),
.B(n_171),
.Y(n_7027)
);

AND2x2_ASAP7_75t_L g7028 ( 
.A(n_6857),
.B(n_172),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6782),
.Y(n_7029)
);

BUFx2_ASAP7_75t_L g7030 ( 
.A(n_6853),
.Y(n_7030)
);

OR2x2_ASAP7_75t_L g7031 ( 
.A(n_6883),
.B(n_172),
.Y(n_7031)
);

OR2x2_ASAP7_75t_L g7032 ( 
.A(n_6878),
.B(n_172),
.Y(n_7032)
);

AND2x2_ASAP7_75t_L g7033 ( 
.A(n_6879),
.B(n_172),
.Y(n_7033)
);

INVx2_ASAP7_75t_L g7034 ( 
.A(n_6856),
.Y(n_7034)
);

HB1xp67_ASAP7_75t_L g7035 ( 
.A(n_6794),
.Y(n_7035)
);

NAND2xp5_ASAP7_75t_L g7036 ( 
.A(n_6796),
.B(n_173),
.Y(n_7036)
);

AOI21xp5_ASAP7_75t_L g7037 ( 
.A1(n_6826),
.A2(n_173),
.B(n_174),
.Y(n_7037)
);

AND2x2_ASAP7_75t_L g7038 ( 
.A(n_6881),
.B(n_173),
.Y(n_7038)
);

AOI221x1_ASAP7_75t_SL g7039 ( 
.A1(n_6804),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.C(n_176),
.Y(n_7039)
);

AND2x2_ASAP7_75t_L g7040 ( 
.A(n_6807),
.B(n_174),
.Y(n_7040)
);

NAND2xp5_ASAP7_75t_L g7041 ( 
.A(n_6863),
.B(n_174),
.Y(n_7041)
);

AND2x2_ASAP7_75t_L g7042 ( 
.A(n_6864),
.B(n_175),
.Y(n_7042)
);

NOR2xp33_ASAP7_75t_R g7043 ( 
.A(n_6882),
.B(n_1071),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_6723),
.Y(n_7044)
);

AND2x2_ASAP7_75t_L g7045 ( 
.A(n_6806),
.B(n_175),
.Y(n_7045)
);

NOR2xp33_ASAP7_75t_R g7046 ( 
.A(n_6723),
.B(n_767),
.Y(n_7046)
);

INVx3_ASAP7_75t_L g7047 ( 
.A(n_6731),
.Y(n_7047)
);

NAND2xp5_ASAP7_75t_L g7048 ( 
.A(n_6736),
.B(n_175),
.Y(n_7048)
);

AND2x2_ASAP7_75t_L g7049 ( 
.A(n_6806),
.B(n_176),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6723),
.Y(n_7050)
);

INVx1_ASAP7_75t_L g7051 ( 
.A(n_6723),
.Y(n_7051)
);

AND2x2_ASAP7_75t_L g7052 ( 
.A(n_6806),
.B(n_176),
.Y(n_7052)
);

INVx1_ASAP7_75t_L g7053 ( 
.A(n_6723),
.Y(n_7053)
);

AND2x4_ASAP7_75t_SL g7054 ( 
.A(n_6718),
.B(n_177),
.Y(n_7054)
);

AND2x2_ASAP7_75t_L g7055 ( 
.A(n_6806),
.B(n_177),
.Y(n_7055)
);

INVx2_ASAP7_75t_SL g7056 ( 
.A(n_6718),
.Y(n_7056)
);

AND2x2_ASAP7_75t_L g7057 ( 
.A(n_6806),
.B(n_177),
.Y(n_7057)
);

OR2x2_ASAP7_75t_L g7058 ( 
.A(n_6759),
.B(n_177),
.Y(n_7058)
);

OR2x2_ASAP7_75t_L g7059 ( 
.A(n_6759),
.B(n_178),
.Y(n_7059)
);

INVx1_ASAP7_75t_SL g7060 ( 
.A(n_6941),
.Y(n_7060)
);

HB1xp67_ASAP7_75t_L g7061 ( 
.A(n_6934),
.Y(n_7061)
);

NAND4xp75_ASAP7_75t_SL g7062 ( 
.A(n_6938),
.B(n_180),
.C(n_178),
.D(n_179),
.Y(n_7062)
);

NOR4xp75_ASAP7_75t_L g7063 ( 
.A(n_7056),
.B(n_180),
.C(n_178),
.D(n_179),
.Y(n_7063)
);

OR2x2_ASAP7_75t_L g7064 ( 
.A(n_7048),
.B(n_179),
.Y(n_7064)
);

OA22x2_ASAP7_75t_L g7065 ( 
.A1(n_7008),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_7065)
);

HB1xp67_ASAP7_75t_L g7066 ( 
.A(n_6923),
.Y(n_7066)
);

AND2x2_ASAP7_75t_L g7067 ( 
.A(n_7045),
.B(n_181),
.Y(n_7067)
);

INVx1_ASAP7_75t_L g7068 ( 
.A(n_6997),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_6884),
.Y(n_7069)
);

INVx2_ASAP7_75t_L g7070 ( 
.A(n_6884),
.Y(n_7070)
);

NOR4xp25_ASAP7_75t_L g7071 ( 
.A(n_7025),
.B(n_183),
.C(n_181),
.D(n_182),
.Y(n_7071)
);

NAND2xp5_ASAP7_75t_L g7072 ( 
.A(n_6989),
.B(n_7047),
.Y(n_7072)
);

HB1xp67_ASAP7_75t_L g7073 ( 
.A(n_7047),
.Y(n_7073)
);

INVx2_ASAP7_75t_SL g7074 ( 
.A(n_6943),
.Y(n_7074)
);

NOR4xp25_ASAP7_75t_L g7075 ( 
.A(n_6908),
.B(n_183),
.C(n_181),
.D(n_182),
.Y(n_7075)
);

NAND2x1p5_ASAP7_75t_L g7076 ( 
.A(n_7008),
.B(n_768),
.Y(n_7076)
);

INVx2_ASAP7_75t_L g7077 ( 
.A(n_6910),
.Y(n_7077)
);

NAND2xp5_ASAP7_75t_L g7078 ( 
.A(n_7049),
.B(n_182),
.Y(n_7078)
);

NOR2xp33_ASAP7_75t_SL g7079 ( 
.A(n_6913),
.B(n_182),
.Y(n_7079)
);

INVx1_ASAP7_75t_L g7080 ( 
.A(n_6997),
.Y(n_7080)
);

XOR2x2_ASAP7_75t_L g7081 ( 
.A(n_6889),
.B(n_183),
.Y(n_7081)
);

OR2x2_ASAP7_75t_L g7082 ( 
.A(n_6891),
.B(n_184),
.Y(n_7082)
);

XNOR2x2_ASAP7_75t_L g7083 ( 
.A(n_6967),
.B(n_6951),
.Y(n_7083)
);

INVx2_ASAP7_75t_SL g7084 ( 
.A(n_6953),
.Y(n_7084)
);

INVx2_ASAP7_75t_L g7085 ( 
.A(n_6982),
.Y(n_7085)
);

BUFx3_ASAP7_75t_L g7086 ( 
.A(n_6920),
.Y(n_7086)
);

HB1xp67_ASAP7_75t_L g7087 ( 
.A(n_6956),
.Y(n_7087)
);

INVx1_ASAP7_75t_L g7088 ( 
.A(n_7054),
.Y(n_7088)
);

NOR2xp33_ASAP7_75t_L g7089 ( 
.A(n_6982),
.B(n_184),
.Y(n_7089)
);

AND2x4_ASAP7_75t_L g7090 ( 
.A(n_6915),
.B(n_184),
.Y(n_7090)
);

INVxp67_ASAP7_75t_L g7091 ( 
.A(n_7052),
.Y(n_7091)
);

NAND4xp75_ASAP7_75t_SL g7092 ( 
.A(n_6927),
.B(n_187),
.C(n_185),
.D(n_186),
.Y(n_7092)
);

NOR3xp33_ASAP7_75t_L g7093 ( 
.A(n_7009),
.B(n_185),
.C(n_186),
.Y(n_7093)
);

XOR2xp5_ASAP7_75t_L g7094 ( 
.A(n_6931),
.B(n_185),
.Y(n_7094)
);

NAND4xp75_ASAP7_75t_L g7095 ( 
.A(n_6909),
.B(n_187),
.C(n_185),
.D(n_186),
.Y(n_7095)
);

NAND2xp5_ASAP7_75t_L g7096 ( 
.A(n_7055),
.B(n_187),
.Y(n_7096)
);

INVx2_ASAP7_75t_L g7097 ( 
.A(n_6952),
.Y(n_7097)
);

INVx1_ASAP7_75t_L g7098 ( 
.A(n_6935),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6972),
.Y(n_7099)
);

AND2x2_ASAP7_75t_L g7100 ( 
.A(n_7057),
.B(n_187),
.Y(n_7100)
);

NOR3xp33_ASAP7_75t_L g7101 ( 
.A(n_7018),
.B(n_188),
.C(n_190),
.Y(n_7101)
);

INVx2_ASAP7_75t_SL g7102 ( 
.A(n_6993),
.Y(n_7102)
);

AND2x2_ASAP7_75t_L g7103 ( 
.A(n_6902),
.B(n_188),
.Y(n_7103)
);

NAND4xp75_ASAP7_75t_L g7104 ( 
.A(n_6944),
.B(n_191),
.C(n_188),
.D(n_190),
.Y(n_7104)
);

INVx1_ASAP7_75t_L g7105 ( 
.A(n_6968),
.Y(n_7105)
);

NAND3xp33_ASAP7_75t_L g7106 ( 
.A(n_6887),
.B(n_188),
.C(n_190),
.Y(n_7106)
);

NAND4xp75_ASAP7_75t_L g7107 ( 
.A(n_6905),
.B(n_192),
.C(n_190),
.D(n_191),
.Y(n_7107)
);

NAND4xp75_ASAP7_75t_L g7108 ( 
.A(n_6942),
.B(n_193),
.C(n_191),
.D(n_192),
.Y(n_7108)
);

INVx1_ASAP7_75t_SL g7109 ( 
.A(n_6986),
.Y(n_7109)
);

AND2x4_ASAP7_75t_L g7110 ( 
.A(n_6939),
.B(n_192),
.Y(n_7110)
);

AOI22xp5_ASAP7_75t_L g7111 ( 
.A1(n_6936),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_7111)
);

INVx1_ASAP7_75t_SL g7112 ( 
.A(n_6958),
.Y(n_7112)
);

INVx1_ASAP7_75t_L g7113 ( 
.A(n_6969),
.Y(n_7113)
);

NAND4xp75_ASAP7_75t_L g7114 ( 
.A(n_6966),
.B(n_6995),
.C(n_6998),
.D(n_6992),
.Y(n_7114)
);

NAND2xp5_ASAP7_75t_L g7115 ( 
.A(n_7039),
.B(n_194),
.Y(n_7115)
);

AOI22xp5_ASAP7_75t_L g7116 ( 
.A1(n_6894),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_7116)
);

INVx2_ASAP7_75t_L g7117 ( 
.A(n_6952),
.Y(n_7117)
);

INVx1_ASAP7_75t_L g7118 ( 
.A(n_6929),
.Y(n_7118)
);

BUFx2_ASAP7_75t_L g7119 ( 
.A(n_7046),
.Y(n_7119)
);

NOR4xp25_ASAP7_75t_L g7120 ( 
.A(n_7013),
.B(n_196),
.C(n_194),
.D(n_195),
.Y(n_7120)
);

NAND2xp5_ASAP7_75t_L g7121 ( 
.A(n_7004),
.B(n_195),
.Y(n_7121)
);

NAND3xp33_ASAP7_75t_L g7122 ( 
.A(n_6961),
.B(n_7002),
.C(n_7011),
.Y(n_7122)
);

AND2x2_ASAP7_75t_L g7123 ( 
.A(n_6954),
.B(n_195),
.Y(n_7123)
);

NAND2xp5_ASAP7_75t_L g7124 ( 
.A(n_6885),
.B(n_196),
.Y(n_7124)
);

BUFx3_ASAP7_75t_L g7125 ( 
.A(n_6922),
.Y(n_7125)
);

INVx2_ASAP7_75t_L g7126 ( 
.A(n_6906),
.Y(n_7126)
);

INVx4_ASAP7_75t_L g7127 ( 
.A(n_7013),
.Y(n_7127)
);

NOR3xp33_ASAP7_75t_L g7128 ( 
.A(n_7027),
.B(n_196),
.C(n_197),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6930),
.Y(n_7129)
);

INVx2_ASAP7_75t_SL g7130 ( 
.A(n_6932),
.Y(n_7130)
);

AND2x2_ASAP7_75t_L g7131 ( 
.A(n_6911),
.B(n_197),
.Y(n_7131)
);

INVx1_ASAP7_75t_L g7132 ( 
.A(n_6899),
.Y(n_7132)
);

AND2x2_ASAP7_75t_L g7133 ( 
.A(n_6949),
.B(n_197),
.Y(n_7133)
);

NAND4xp75_ASAP7_75t_SL g7134 ( 
.A(n_6918),
.B(n_200),
.C(n_198),
.D(n_199),
.Y(n_7134)
);

NAND4xp75_ASAP7_75t_SL g7135 ( 
.A(n_6950),
.B(n_200),
.C(n_198),
.D(n_199),
.Y(n_7135)
);

AND2x4_ASAP7_75t_L g7136 ( 
.A(n_7007),
.B(n_198),
.Y(n_7136)
);

INVxp33_ASAP7_75t_L g7137 ( 
.A(n_6979),
.Y(n_7137)
);

INVx2_ASAP7_75t_SL g7138 ( 
.A(n_7016),
.Y(n_7138)
);

INVx1_ASAP7_75t_SL g7139 ( 
.A(n_6963),
.Y(n_7139)
);

INVx1_ASAP7_75t_L g7140 ( 
.A(n_6904),
.Y(n_7140)
);

NOR2xp33_ASAP7_75t_L g7141 ( 
.A(n_6947),
.B(n_199),
.Y(n_7141)
);

XOR2x2_ASAP7_75t_L g7142 ( 
.A(n_6903),
.B(n_200),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_6983),
.Y(n_7143)
);

BUFx3_ASAP7_75t_L g7144 ( 
.A(n_7026),
.Y(n_7144)
);

OR2x2_ASAP7_75t_L g7145 ( 
.A(n_7019),
.B(n_200),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6985),
.Y(n_7146)
);

NAND4xp75_ASAP7_75t_L g7147 ( 
.A(n_6928),
.B(n_203),
.C(n_201),
.D(n_202),
.Y(n_7147)
);

INVx1_ASAP7_75t_L g7148 ( 
.A(n_6987),
.Y(n_7148)
);

INVx1_ASAP7_75t_L g7149 ( 
.A(n_6964),
.Y(n_7149)
);

INVx1_ASAP7_75t_L g7150 ( 
.A(n_6981),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_6926),
.Y(n_7151)
);

AND2x2_ASAP7_75t_L g7152 ( 
.A(n_6895),
.B(n_201),
.Y(n_7152)
);

AND2x4_ASAP7_75t_L g7153 ( 
.A(n_6971),
.B(n_201),
.Y(n_7153)
);

NAND4xp75_ASAP7_75t_SL g7154 ( 
.A(n_6948),
.B(n_204),
.C(n_202),
.D(n_203),
.Y(n_7154)
);

INVx1_ASAP7_75t_L g7155 ( 
.A(n_6886),
.Y(n_7155)
);

NAND2xp5_ASAP7_75t_L g7156 ( 
.A(n_7033),
.B(n_202),
.Y(n_7156)
);

XOR2x2_ASAP7_75t_L g7157 ( 
.A(n_6901),
.B(n_202),
.Y(n_7157)
);

AND2x2_ASAP7_75t_L g7158 ( 
.A(n_6907),
.B(n_203),
.Y(n_7158)
);

INVx2_ASAP7_75t_L g7159 ( 
.A(n_6914),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_6888),
.Y(n_7160)
);

INVx2_ASAP7_75t_L g7161 ( 
.A(n_7034),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_7044),
.Y(n_7162)
);

INVx2_ASAP7_75t_L g7163 ( 
.A(n_6917),
.Y(n_7163)
);

INVx3_ASAP7_75t_L g7164 ( 
.A(n_7014),
.Y(n_7164)
);

NAND3xp33_ASAP7_75t_L g7165 ( 
.A(n_7036),
.B(n_203),
.C(n_204),
.Y(n_7165)
);

NOR3xp33_ASAP7_75t_L g7166 ( 
.A(n_7041),
.B(n_204),
.C(n_205),
.Y(n_7166)
);

NAND3xp33_ASAP7_75t_SL g7167 ( 
.A(n_7043),
.B(n_204),
.C(n_205),
.Y(n_7167)
);

AND2x4_ASAP7_75t_SL g7168 ( 
.A(n_6897),
.B(n_205),
.Y(n_7168)
);

XOR2x2_ASAP7_75t_L g7169 ( 
.A(n_6975),
.B(n_205),
.Y(n_7169)
);

AND2x2_ASAP7_75t_L g7170 ( 
.A(n_6973),
.B(n_206),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_7050),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_7051),
.Y(n_7172)
);

INVx6_ASAP7_75t_L g7173 ( 
.A(n_7058),
.Y(n_7173)
);

INVx3_ASAP7_75t_L g7174 ( 
.A(n_6991),
.Y(n_7174)
);

XNOR2x1_ASAP7_75t_L g7175 ( 
.A(n_7022),
.B(n_206),
.Y(n_7175)
);

NAND4xp75_ASAP7_75t_L g7176 ( 
.A(n_6890),
.B(n_208),
.C(n_206),
.D(n_207),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_7053),
.Y(n_7177)
);

INVx2_ASAP7_75t_SL g7178 ( 
.A(n_7059),
.Y(n_7178)
);

NAND2xp5_ASAP7_75t_SL g7179 ( 
.A(n_6970),
.B(n_207),
.Y(n_7179)
);

OR2x2_ASAP7_75t_L g7180 ( 
.A(n_7031),
.B(n_207),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_6892),
.Y(n_7181)
);

INVx2_ASAP7_75t_L g7182 ( 
.A(n_6896),
.Y(n_7182)
);

AND2x2_ASAP7_75t_L g7183 ( 
.A(n_6912),
.B(n_208),
.Y(n_7183)
);

INVx5_ASAP7_75t_L g7184 ( 
.A(n_7038),
.Y(n_7184)
);

XOR2x2_ASAP7_75t_L g7185 ( 
.A(n_6925),
.B(n_208),
.Y(n_7185)
);

NAND4xp75_ASAP7_75t_L g7186 ( 
.A(n_7029),
.B(n_211),
.C(n_209),
.D(n_210),
.Y(n_7186)
);

NAND2xp5_ASAP7_75t_L g7187 ( 
.A(n_6990),
.B(n_209),
.Y(n_7187)
);

NAND4xp75_ASAP7_75t_L g7188 ( 
.A(n_6919),
.B(n_211),
.C(n_209),
.D(n_210),
.Y(n_7188)
);

AND2x2_ASAP7_75t_L g7189 ( 
.A(n_7006),
.B(n_6946),
.Y(n_7189)
);

HB1xp67_ASAP7_75t_L g7190 ( 
.A(n_6924),
.Y(n_7190)
);

NOR2x1_ASAP7_75t_L g7191 ( 
.A(n_7032),
.B(n_209),
.Y(n_7191)
);

BUFx2_ASAP7_75t_SL g7192 ( 
.A(n_7040),
.Y(n_7192)
);

AND2x4_ASAP7_75t_L g7193 ( 
.A(n_6999),
.B(n_210),
.Y(n_7193)
);

INVx2_ASAP7_75t_L g7194 ( 
.A(n_7024),
.Y(n_7194)
);

AND2x2_ASAP7_75t_L g7195 ( 
.A(n_6937),
.B(n_210),
.Y(n_7195)
);

INVx1_ASAP7_75t_L g7196 ( 
.A(n_7028),
.Y(n_7196)
);

INVx1_ASAP7_75t_L g7197 ( 
.A(n_7042),
.Y(n_7197)
);

AOI22xp5_ASAP7_75t_L g7198 ( 
.A1(n_6893),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_7198)
);

AND2x2_ASAP7_75t_L g7199 ( 
.A(n_6957),
.B(n_211),
.Y(n_7199)
);

INVx1_ASAP7_75t_L g7200 ( 
.A(n_6996),
.Y(n_7200)
);

OR2x2_ASAP7_75t_L g7201 ( 
.A(n_6960),
.B(n_6900),
.Y(n_7201)
);

AND2x2_ASAP7_75t_L g7202 ( 
.A(n_7023),
.B(n_212),
.Y(n_7202)
);

INVx3_ASAP7_75t_L g7203 ( 
.A(n_6916),
.Y(n_7203)
);

INVx2_ASAP7_75t_L g7204 ( 
.A(n_7069),
.Y(n_7204)
);

OR2x6_ASAP7_75t_L g7205 ( 
.A(n_7076),
.B(n_7037),
.Y(n_7205)
);

AND2x2_ASAP7_75t_L g7206 ( 
.A(n_7060),
.B(n_7152),
.Y(n_7206)
);

AND2x2_ASAP7_75t_L g7207 ( 
.A(n_7158),
.B(n_6955),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_7065),
.Y(n_7208)
);

INVx1_ASAP7_75t_L g7209 ( 
.A(n_7066),
.Y(n_7209)
);

AND2x2_ASAP7_75t_L g7210 ( 
.A(n_7183),
.B(n_7012),
.Y(n_7210)
);

NAND2xp5_ASAP7_75t_L g7211 ( 
.A(n_7070),
.B(n_7005),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_7061),
.Y(n_7212)
);

NAND2xp5_ASAP7_75t_L g7213 ( 
.A(n_7071),
.B(n_7112),
.Y(n_7213)
);

INVx1_ASAP7_75t_SL g7214 ( 
.A(n_7086),
.Y(n_7214)
);

INVx1_ASAP7_75t_L g7215 ( 
.A(n_7073),
.Y(n_7215)
);

NAND2xp67_ASAP7_75t_L g7216 ( 
.A(n_7168),
.B(n_7017),
.Y(n_7216)
);

NAND2xp5_ASAP7_75t_L g7217 ( 
.A(n_7077),
.B(n_7075),
.Y(n_7217)
);

INVx1_ASAP7_75t_SL g7218 ( 
.A(n_7109),
.Y(n_7218)
);

AND2x2_ASAP7_75t_L g7219 ( 
.A(n_7195),
.B(n_6976),
.Y(n_7219)
);

NAND2xp5_ASAP7_75t_L g7220 ( 
.A(n_7120),
.B(n_7021),
.Y(n_7220)
);

INVx2_ASAP7_75t_L g7221 ( 
.A(n_7097),
.Y(n_7221)
);

NAND2xp5_ASAP7_75t_L g7222 ( 
.A(n_7074),
.B(n_7030),
.Y(n_7222)
);

INVx1_ASAP7_75t_L g7223 ( 
.A(n_7108),
.Y(n_7223)
);

OR2x6_ASAP7_75t_L g7224 ( 
.A(n_7084),
.B(n_7000),
.Y(n_7224)
);

AND2x2_ASAP7_75t_L g7225 ( 
.A(n_7170),
.B(n_7067),
.Y(n_7225)
);

NAND2x1p5_ASAP7_75t_L g7226 ( 
.A(n_7088),
.B(n_6940),
.Y(n_7226)
);

NAND2xp5_ASAP7_75t_L g7227 ( 
.A(n_7102),
.B(n_7020),
.Y(n_7227)
);

INVx2_ASAP7_75t_L g7228 ( 
.A(n_7117),
.Y(n_7228)
);

AND2x4_ASAP7_75t_L g7229 ( 
.A(n_7085),
.B(n_7003),
.Y(n_7229)
);

INVx1_ASAP7_75t_L g7230 ( 
.A(n_7082),
.Y(n_7230)
);

AND2x2_ASAP7_75t_L g7231 ( 
.A(n_7100),
.B(n_7103),
.Y(n_7231)
);

INVx2_ASAP7_75t_L g7232 ( 
.A(n_7127),
.Y(n_7232)
);

INVx1_ASAP7_75t_L g7233 ( 
.A(n_7083),
.Y(n_7233)
);

INVx2_ASAP7_75t_SL g7234 ( 
.A(n_7144),
.Y(n_7234)
);

NAND2xp5_ASAP7_75t_L g7235 ( 
.A(n_7199),
.B(n_7015),
.Y(n_7235)
);

NAND2xp5_ASAP7_75t_L g7236 ( 
.A(n_7131),
.B(n_6977),
.Y(n_7236)
);

NAND2xp5_ASAP7_75t_L g7237 ( 
.A(n_7123),
.B(n_6978),
.Y(n_7237)
);

INVx1_ASAP7_75t_L g7238 ( 
.A(n_7072),
.Y(n_7238)
);

BUFx3_ASAP7_75t_L g7239 ( 
.A(n_7099),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_7186),
.Y(n_7240)
);

NAND2xp5_ASAP7_75t_L g7241 ( 
.A(n_7202),
.B(n_7010),
.Y(n_7241)
);

OR2x2_ASAP7_75t_L g7242 ( 
.A(n_7150),
.B(n_6945),
.Y(n_7242)
);

INVx1_ASAP7_75t_SL g7243 ( 
.A(n_7110),
.Y(n_7243)
);

INVx1_ASAP7_75t_L g7244 ( 
.A(n_7087),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_7094),
.Y(n_7245)
);

NOR2x1p5_ASAP7_75t_L g7246 ( 
.A(n_7114),
.B(n_6984),
.Y(n_7246)
);

INVx1_ASAP7_75t_L g7247 ( 
.A(n_7095),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_7107),
.Y(n_7248)
);

OR2x2_ASAP7_75t_L g7249 ( 
.A(n_7149),
.B(n_6980),
.Y(n_7249)
);

INVx1_ASAP7_75t_L g7250 ( 
.A(n_7068),
.Y(n_7250)
);

AND2x2_ASAP7_75t_L g7251 ( 
.A(n_7133),
.B(n_6974),
.Y(n_7251)
);

NAND2xp5_ASAP7_75t_L g7252 ( 
.A(n_7189),
.B(n_6962),
.Y(n_7252)
);

AND2x2_ASAP7_75t_L g7253 ( 
.A(n_7129),
.B(n_6965),
.Y(n_7253)
);

NOR2xp33_ASAP7_75t_L g7254 ( 
.A(n_7167),
.B(n_7079),
.Y(n_7254)
);

OR2x2_ASAP7_75t_L g7255 ( 
.A(n_7124),
.B(n_6994),
.Y(n_7255)
);

INVx2_ASAP7_75t_SL g7256 ( 
.A(n_7125),
.Y(n_7256)
);

INVx2_ASAP7_75t_L g7257 ( 
.A(n_7159),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_7080),
.Y(n_7258)
);

AND2x2_ASAP7_75t_L g7259 ( 
.A(n_7193),
.B(n_6898),
.Y(n_7259)
);

NAND2xp5_ASAP7_75t_L g7260 ( 
.A(n_7184),
.B(n_7035),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_7121),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_7192),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_7176),
.Y(n_7263)
);

AOI21xp33_ASAP7_75t_SL g7264 ( 
.A1(n_7115),
.A2(n_7001),
.B(n_6921),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_7136),
.Y(n_7265)
);

NAND2xp5_ASAP7_75t_L g7266 ( 
.A(n_7184),
.B(n_6959),
.Y(n_7266)
);

AND2x2_ASAP7_75t_L g7267 ( 
.A(n_7105),
.B(n_6988),
.Y(n_7267)
);

AND2x2_ASAP7_75t_L g7268 ( 
.A(n_7113),
.B(n_7143),
.Y(n_7268)
);

NAND2xp5_ASAP7_75t_L g7269 ( 
.A(n_7184),
.B(n_6933),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_7147),
.Y(n_7270)
);

NAND2x1_ASAP7_75t_L g7271 ( 
.A(n_7173),
.B(n_213),
.Y(n_7271)
);

INVx2_ASAP7_75t_L g7272 ( 
.A(n_7138),
.Y(n_7272)
);

AND2x2_ASAP7_75t_L g7273 ( 
.A(n_7146),
.B(n_213),
.Y(n_7273)
);

AOI222xp33_ASAP7_75t_L g7274 ( 
.A1(n_7139),
.A2(n_216),
.B1(n_218),
.B2(n_214),
.C1(n_215),
.C2(n_217),
.Y(n_7274)
);

INVx3_ASAP7_75t_L g7275 ( 
.A(n_7090),
.Y(n_7275)
);

OR2x2_ASAP7_75t_L g7276 ( 
.A(n_7187),
.B(n_7145),
.Y(n_7276)
);

AND2x2_ASAP7_75t_L g7277 ( 
.A(n_7163),
.B(n_214),
.Y(n_7277)
);

AND2x2_ASAP7_75t_L g7278 ( 
.A(n_7132),
.B(n_214),
.Y(n_7278)
);

NAND2xp5_ASAP7_75t_SL g7279 ( 
.A(n_7116),
.B(n_214),
.Y(n_7279)
);

HB1xp67_ASAP7_75t_L g7280 ( 
.A(n_7063),
.Y(n_7280)
);

NAND2xp5_ASAP7_75t_L g7281 ( 
.A(n_7089),
.B(n_7141),
.Y(n_7281)
);

INVx2_ASAP7_75t_L g7282 ( 
.A(n_7161),
.Y(n_7282)
);

NAND2xp5_ASAP7_75t_L g7283 ( 
.A(n_7151),
.B(n_215),
.Y(n_7283)
);

INVx2_ASAP7_75t_L g7284 ( 
.A(n_7130),
.Y(n_7284)
);

AND2x4_ASAP7_75t_L g7285 ( 
.A(n_7126),
.B(n_215),
.Y(n_7285)
);

NAND2xp5_ASAP7_75t_L g7286 ( 
.A(n_7188),
.B(n_215),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_7180),
.Y(n_7287)
);

AND2x4_ASAP7_75t_L g7288 ( 
.A(n_7153),
.B(n_7200),
.Y(n_7288)
);

INVxp67_ASAP7_75t_L g7289 ( 
.A(n_7104),
.Y(n_7289)
);

AND2x2_ASAP7_75t_L g7290 ( 
.A(n_7203),
.B(n_216),
.Y(n_7290)
);

OR2x2_ASAP7_75t_L g7291 ( 
.A(n_7156),
.B(n_216),
.Y(n_7291)
);

NAND3xp33_ASAP7_75t_L g7292 ( 
.A(n_7106),
.B(n_216),
.C(n_217),
.Y(n_7292)
);

CKINVDCx16_ASAP7_75t_R g7293 ( 
.A(n_7064),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_7078),
.Y(n_7294)
);

OR2x2_ASAP7_75t_L g7295 ( 
.A(n_7096),
.B(n_217),
.Y(n_7295)
);

OAI32xp33_ASAP7_75t_L g7296 ( 
.A1(n_7137),
.A2(n_219),
.A3(n_217),
.B1(n_218),
.B2(n_220),
.Y(n_7296)
);

NAND2xp5_ASAP7_75t_L g7297 ( 
.A(n_7091),
.B(n_218),
.Y(n_7297)
);

OR2x2_ASAP7_75t_L g7298 ( 
.A(n_7201),
.B(n_7118),
.Y(n_7298)
);

NAND2xp67_ASAP7_75t_SL g7299 ( 
.A(n_7092),
.B(n_218),
.Y(n_7299)
);

INVx1_ASAP7_75t_L g7300 ( 
.A(n_7190),
.Y(n_7300)
);

INVx1_ASAP7_75t_L g7301 ( 
.A(n_7119),
.Y(n_7301)
);

INVx2_ASAP7_75t_L g7302 ( 
.A(n_7173),
.Y(n_7302)
);

INVx2_ASAP7_75t_L g7303 ( 
.A(n_7182),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_7119),
.Y(n_7304)
);

AND2x2_ASAP7_75t_L g7305 ( 
.A(n_7194),
.B(n_7174),
.Y(n_7305)
);

AND2x2_ASAP7_75t_L g7306 ( 
.A(n_7196),
.B(n_219),
.Y(n_7306)
);

AND2x4_ASAP7_75t_SL g7307 ( 
.A(n_7164),
.B(n_219),
.Y(n_7307)
);

OR2x2_ASAP7_75t_L g7308 ( 
.A(n_7179),
.B(n_219),
.Y(n_7308)
);

INVx1_ASAP7_75t_L g7309 ( 
.A(n_7191),
.Y(n_7309)
);

AND2x4_ASAP7_75t_L g7310 ( 
.A(n_7178),
.B(n_220),
.Y(n_7310)
);

AND2x2_ASAP7_75t_L g7311 ( 
.A(n_7197),
.B(n_220),
.Y(n_7311)
);

AND2x2_ASAP7_75t_L g7312 ( 
.A(n_7140),
.B(n_220),
.Y(n_7312)
);

INVx2_ASAP7_75t_L g7313 ( 
.A(n_7098),
.Y(n_7313)
);

OR2x2_ASAP7_75t_L g7314 ( 
.A(n_7122),
.B(n_221),
.Y(n_7314)
);

OR2x2_ASAP7_75t_L g7315 ( 
.A(n_7148),
.B(n_221),
.Y(n_7315)
);

OR2x2_ASAP7_75t_L g7316 ( 
.A(n_7165),
.B(n_221),
.Y(n_7316)
);

AOI22xp33_ASAP7_75t_L g7317 ( 
.A1(n_7093),
.A2(n_224),
.B1(n_221),
.B2(n_223),
.Y(n_7317)
);

INVx1_ASAP7_75t_SL g7318 ( 
.A(n_7134),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_7198),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_7128),
.B(n_223),
.Y(n_7320)
);

AND3x2_ASAP7_75t_L g7321 ( 
.A(n_7166),
.B(n_223),
.C(n_224),
.Y(n_7321)
);

INVx2_ASAP7_75t_L g7322 ( 
.A(n_7155),
.Y(n_7322)
);

OR2x2_ASAP7_75t_L g7323 ( 
.A(n_7160),
.B(n_7162),
.Y(n_7323)
);

AND2x2_ASAP7_75t_L g7324 ( 
.A(n_7175),
.B(n_223),
.Y(n_7324)
);

NAND2xp5_ASAP7_75t_L g7325 ( 
.A(n_7111),
.B(n_225),
.Y(n_7325)
);

INVx1_ASAP7_75t_L g7326 ( 
.A(n_7171),
.Y(n_7326)
);

OR2x2_ASAP7_75t_L g7327 ( 
.A(n_7172),
.B(n_225),
.Y(n_7327)
);

INVx4_ASAP7_75t_L g7328 ( 
.A(n_7142),
.Y(n_7328)
);

AND2x2_ASAP7_75t_SL g7329 ( 
.A(n_7101),
.B(n_225),
.Y(n_7329)
);

HB1xp67_ASAP7_75t_L g7330 ( 
.A(n_7154),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_7177),
.Y(n_7331)
);

NAND2xp5_ASAP7_75t_L g7332 ( 
.A(n_7081),
.B(n_226),
.Y(n_7332)
);

INVx2_ASAP7_75t_L g7333 ( 
.A(n_7181),
.Y(n_7333)
);

INVxp67_ASAP7_75t_L g7334 ( 
.A(n_7157),
.Y(n_7334)
);

AND2x2_ASAP7_75t_L g7335 ( 
.A(n_7169),
.B(n_226),
.Y(n_7335)
);

NOR2x1_ASAP7_75t_L g7336 ( 
.A(n_7135),
.B(n_226),
.Y(n_7336)
);

AND2x2_ASAP7_75t_L g7337 ( 
.A(n_7185),
.B(n_227),
.Y(n_7337)
);

AND2x2_ASAP7_75t_L g7338 ( 
.A(n_7062),
.B(n_227),
.Y(n_7338)
);

INVx2_ASAP7_75t_L g7339 ( 
.A(n_7069),
.Y(n_7339)
);

NOR2xp33_ASAP7_75t_L g7340 ( 
.A(n_7060),
.B(n_227),
.Y(n_7340)
);

AND2x2_ASAP7_75t_L g7341 ( 
.A(n_7060),
.B(n_228),
.Y(n_7341)
);

INVx1_ASAP7_75t_L g7342 ( 
.A(n_7065),
.Y(n_7342)
);

NAND2xp5_ASAP7_75t_L g7343 ( 
.A(n_7060),
.B(n_228),
.Y(n_7343)
);

OR2x2_ASAP7_75t_L g7344 ( 
.A(n_7060),
.B(n_228),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_7060),
.B(n_228),
.Y(n_7345)
);

AND2x4_ASAP7_75t_L g7346 ( 
.A(n_7069),
.B(n_229),
.Y(n_7346)
);

AND2x2_ASAP7_75t_L g7347 ( 
.A(n_7060),
.B(n_229),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_7065),
.Y(n_7348)
);

NAND2xp5_ASAP7_75t_L g7349 ( 
.A(n_7060),
.B(n_229),
.Y(n_7349)
);

AND2x4_ASAP7_75t_L g7350 ( 
.A(n_7204),
.B(n_229),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_L g7351 ( 
.A(n_7233),
.B(n_230),
.Y(n_7351)
);

AND2x2_ASAP7_75t_L g7352 ( 
.A(n_7206),
.B(n_230),
.Y(n_7352)
);

NAND2xp5_ASAP7_75t_L g7353 ( 
.A(n_7214),
.B(n_230),
.Y(n_7353)
);

HB1xp67_ASAP7_75t_L g7354 ( 
.A(n_7339),
.Y(n_7354)
);

NAND2xp5_ASAP7_75t_SL g7355 ( 
.A(n_7257),
.B(n_230),
.Y(n_7355)
);

INVx2_ASAP7_75t_L g7356 ( 
.A(n_7256),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_7341),
.Y(n_7357)
);

OAI22xp33_ASAP7_75t_L g7358 ( 
.A1(n_7318),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_7358)
);

NAND2xp5_ASAP7_75t_L g7359 ( 
.A(n_7234),
.B(n_231),
.Y(n_7359)
);

NAND2xp5_ASAP7_75t_L g7360 ( 
.A(n_7208),
.B(n_231),
.Y(n_7360)
);

BUFx3_ASAP7_75t_L g7361 ( 
.A(n_7232),
.Y(n_7361)
);

NOR2xp33_ASAP7_75t_L g7362 ( 
.A(n_7342),
.B(n_231),
.Y(n_7362)
);

AND2x2_ASAP7_75t_L g7363 ( 
.A(n_7345),
.B(n_233),
.Y(n_7363)
);

INVx2_ASAP7_75t_L g7364 ( 
.A(n_7221),
.Y(n_7364)
);

AND2x2_ASAP7_75t_L g7365 ( 
.A(n_7347),
.B(n_233),
.Y(n_7365)
);

AOI21xp33_ASAP7_75t_R g7366 ( 
.A1(n_7348),
.A2(n_234),
.B(n_235),
.Y(n_7366)
);

BUFx3_ASAP7_75t_L g7367 ( 
.A(n_7302),
.Y(n_7367)
);

NAND2xp5_ASAP7_75t_L g7368 ( 
.A(n_7285),
.B(n_234),
.Y(n_7368)
);

INVx2_ASAP7_75t_SL g7369 ( 
.A(n_7228),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_7338),
.Y(n_7370)
);

AND2x2_ASAP7_75t_L g7371 ( 
.A(n_7207),
.B(n_234),
.Y(n_7371)
);

NAND2xp5_ASAP7_75t_L g7372 ( 
.A(n_7285),
.B(n_235),
.Y(n_7372)
);

OR2x2_ASAP7_75t_L g7373 ( 
.A(n_7298),
.B(n_235),
.Y(n_7373)
);

NAND2xp33_ASAP7_75t_SL g7374 ( 
.A(n_7280),
.B(n_235),
.Y(n_7374)
);

BUFx4f_ASAP7_75t_SL g7375 ( 
.A(n_7218),
.Y(n_7375)
);

INVx1_ASAP7_75t_L g7376 ( 
.A(n_7290),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_7277),
.Y(n_7377)
);

NAND2xp5_ASAP7_75t_L g7378 ( 
.A(n_7346),
.B(n_236),
.Y(n_7378)
);

OR2x2_ASAP7_75t_L g7379 ( 
.A(n_7284),
.B(n_236),
.Y(n_7379)
);

AOI21xp33_ASAP7_75t_SL g7380 ( 
.A1(n_7286),
.A2(n_236),
.B(n_237),
.Y(n_7380)
);

OR2x2_ASAP7_75t_L g7381 ( 
.A(n_7344),
.B(n_237),
.Y(n_7381)
);

INVx1_ASAP7_75t_SL g7382 ( 
.A(n_7243),
.Y(n_7382)
);

NAND2xp5_ASAP7_75t_L g7383 ( 
.A(n_7321),
.B(n_237),
.Y(n_7383)
);

INVx2_ASAP7_75t_SL g7384 ( 
.A(n_7272),
.Y(n_7384)
);

INVx2_ASAP7_75t_L g7385 ( 
.A(n_7282),
.Y(n_7385)
);

INVx1_ASAP7_75t_L g7386 ( 
.A(n_7343),
.Y(n_7386)
);

AND2x2_ASAP7_75t_L g7387 ( 
.A(n_7219),
.B(n_237),
.Y(n_7387)
);

CKINVDCx5p33_ASAP7_75t_R g7388 ( 
.A(n_7239),
.Y(n_7388)
);

O2A1O1Ixp5_ASAP7_75t_L g7389 ( 
.A1(n_7213),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_7389)
);

INVx1_ASAP7_75t_L g7390 ( 
.A(n_7349),
.Y(n_7390)
);

INVx2_ASAP7_75t_L g7391 ( 
.A(n_7226),
.Y(n_7391)
);

INVx1_ASAP7_75t_L g7392 ( 
.A(n_7340),
.Y(n_7392)
);

NAND2xp5_ASAP7_75t_L g7393 ( 
.A(n_7310),
.B(n_238),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7271),
.Y(n_7394)
);

NAND2xp5_ASAP7_75t_L g7395 ( 
.A(n_7262),
.B(n_7273),
.Y(n_7395)
);

NAND2xp5_ASAP7_75t_L g7396 ( 
.A(n_7336),
.B(n_238),
.Y(n_7396)
);

NOR2xp33_ASAP7_75t_SL g7397 ( 
.A(n_7215),
.B(n_7303),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_7307),
.Y(n_7398)
);

INVxp67_ASAP7_75t_L g7399 ( 
.A(n_7330),
.Y(n_7399)
);

AND2x2_ASAP7_75t_L g7400 ( 
.A(n_7231),
.B(n_238),
.Y(n_7400)
);

INVx1_ASAP7_75t_L g7401 ( 
.A(n_7216),
.Y(n_7401)
);

AND2x2_ASAP7_75t_L g7402 ( 
.A(n_7225),
.B(n_239),
.Y(n_7402)
);

NAND2xp5_ASAP7_75t_L g7403 ( 
.A(n_7278),
.B(n_239),
.Y(n_7403)
);

OAI22xp5_ASAP7_75t_L g7404 ( 
.A1(n_7289),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_7316),
.Y(n_7405)
);

NAND2xp5_ASAP7_75t_L g7406 ( 
.A(n_7312),
.B(n_240),
.Y(n_7406)
);

NAND2xp5_ASAP7_75t_L g7407 ( 
.A(n_7335),
.B(n_240),
.Y(n_7407)
);

NAND2xp5_ASAP7_75t_L g7408 ( 
.A(n_7324),
.B(n_241),
.Y(n_7408)
);

NAND2xp5_ASAP7_75t_L g7409 ( 
.A(n_7274),
.B(n_7337),
.Y(n_7409)
);

INVx1_ASAP7_75t_SL g7410 ( 
.A(n_7305),
.Y(n_7410)
);

NAND2xp5_ASAP7_75t_L g7411 ( 
.A(n_7210),
.B(n_241),
.Y(n_7411)
);

NAND2xp5_ASAP7_75t_L g7412 ( 
.A(n_7306),
.B(n_7311),
.Y(n_7412)
);

AND2x2_ASAP7_75t_L g7413 ( 
.A(n_7267),
.B(n_242),
.Y(n_7413)
);

INVx1_ASAP7_75t_L g7414 ( 
.A(n_7217),
.Y(n_7414)
);

OR2x2_ASAP7_75t_L g7415 ( 
.A(n_7209),
.B(n_242),
.Y(n_7415)
);

NAND2xp5_ASAP7_75t_L g7416 ( 
.A(n_7212),
.B(n_242),
.Y(n_7416)
);

NAND2xp5_ASAP7_75t_L g7417 ( 
.A(n_7288),
.B(n_243),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_7222),
.Y(n_7418)
);

NAND2xp5_ASAP7_75t_SL g7419 ( 
.A(n_7313),
.B(n_243),
.Y(n_7419)
);

OR2x2_ASAP7_75t_L g7420 ( 
.A(n_7205),
.B(n_243),
.Y(n_7420)
);

INVxp67_ASAP7_75t_L g7421 ( 
.A(n_7254),
.Y(n_7421)
);

NAND2xp5_ASAP7_75t_L g7422 ( 
.A(n_7223),
.B(n_243),
.Y(n_7422)
);

NAND2x1_ASAP7_75t_SL g7423 ( 
.A(n_7240),
.B(n_244),
.Y(n_7423)
);

INVx2_ASAP7_75t_L g7424 ( 
.A(n_7275),
.Y(n_7424)
);

OR2x2_ASAP7_75t_L g7425 ( 
.A(n_7205),
.B(n_244),
.Y(n_7425)
);

OR2x6_ASAP7_75t_L g7426 ( 
.A(n_7266),
.B(n_768),
.Y(n_7426)
);

NAND2xp5_ASAP7_75t_L g7427 ( 
.A(n_7268),
.B(n_7247),
.Y(n_7427)
);

NAND2xp5_ASAP7_75t_L g7428 ( 
.A(n_7248),
.B(n_244),
.Y(n_7428)
);

NOR2xp33_ASAP7_75t_L g7429 ( 
.A(n_7328),
.B(n_244),
.Y(n_7429)
);

NOR2xp33_ASAP7_75t_L g7430 ( 
.A(n_7270),
.B(n_245),
.Y(n_7430)
);

INVx1_ASAP7_75t_L g7431 ( 
.A(n_7260),
.Y(n_7431)
);

AND2x2_ASAP7_75t_L g7432 ( 
.A(n_7259),
.B(n_245),
.Y(n_7432)
);

INVx2_ASAP7_75t_SL g7433 ( 
.A(n_7229),
.Y(n_7433)
);

NAND2xp5_ASAP7_75t_L g7434 ( 
.A(n_7317),
.B(n_245),
.Y(n_7434)
);

INVx1_ASAP7_75t_SL g7435 ( 
.A(n_7269),
.Y(n_7435)
);

HB1xp67_ASAP7_75t_L g7436 ( 
.A(n_7244),
.Y(n_7436)
);

INVx2_ASAP7_75t_L g7437 ( 
.A(n_7229),
.Y(n_7437)
);

CKINVDCx16_ASAP7_75t_R g7438 ( 
.A(n_7293),
.Y(n_7438)
);

AND2x2_ASAP7_75t_L g7439 ( 
.A(n_7251),
.B(n_246),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_7327),
.Y(n_7440)
);

INVx2_ASAP7_75t_L g7441 ( 
.A(n_7361),
.Y(n_7441)
);

NOR2xp33_ASAP7_75t_L g7442 ( 
.A(n_7375),
.B(n_7263),
.Y(n_7442)
);

INVxp67_ASAP7_75t_SL g7443 ( 
.A(n_7354),
.Y(n_7443)
);

INVx2_ASAP7_75t_L g7444 ( 
.A(n_7367),
.Y(n_7444)
);

OAI211xp5_ASAP7_75t_L g7445 ( 
.A1(n_7380),
.A2(n_7264),
.B(n_7332),
.C(n_7334),
.Y(n_7445)
);

INVx2_ASAP7_75t_L g7446 ( 
.A(n_7356),
.Y(n_7446)
);

INVx1_ASAP7_75t_L g7447 ( 
.A(n_7368),
.Y(n_7447)
);

OR2x2_ASAP7_75t_L g7448 ( 
.A(n_7438),
.B(n_7211),
.Y(n_7448)
);

NAND2x1p5_ASAP7_75t_L g7449 ( 
.A(n_7384),
.B(n_7301),
.Y(n_7449)
);

NAND2xp5_ASAP7_75t_L g7450 ( 
.A(n_7433),
.B(n_7300),
.Y(n_7450)
);

OR2x2_ASAP7_75t_L g7451 ( 
.A(n_7410),
.B(n_7242),
.Y(n_7451)
);

NOR2xp67_ASAP7_75t_L g7452 ( 
.A(n_7369),
.B(n_7304),
.Y(n_7452)
);

BUFx2_ASAP7_75t_L g7453 ( 
.A(n_7350),
.Y(n_7453)
);

NAND2xp5_ASAP7_75t_L g7454 ( 
.A(n_7382),
.B(n_7245),
.Y(n_7454)
);

NOR2xp33_ASAP7_75t_L g7455 ( 
.A(n_7435),
.B(n_7315),
.Y(n_7455)
);

INVxp67_ASAP7_75t_L g7456 ( 
.A(n_7397),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_7372),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_7350),
.Y(n_7458)
);

NAND2xp5_ASAP7_75t_L g7459 ( 
.A(n_7364),
.B(n_7250),
.Y(n_7459)
);

AND2x2_ASAP7_75t_L g7460 ( 
.A(n_7387),
.B(n_7253),
.Y(n_7460)
);

OAI21xp33_ASAP7_75t_L g7461 ( 
.A1(n_7427),
.A2(n_7238),
.B(n_7227),
.Y(n_7461)
);

NOR2xp33_ASAP7_75t_L g7462 ( 
.A(n_7370),
.B(n_7314),
.Y(n_7462)
);

OR2x2_ASAP7_75t_L g7463 ( 
.A(n_7437),
.B(n_7308),
.Y(n_7463)
);

OAI22xp5_ASAP7_75t_L g7464 ( 
.A1(n_7391),
.A2(n_7249),
.B1(n_7319),
.B2(n_7283),
.Y(n_7464)
);

OR2x2_ASAP7_75t_L g7465 ( 
.A(n_7385),
.B(n_7258),
.Y(n_7465)
);

NOR2xp33_ASAP7_75t_SL g7466 ( 
.A(n_7388),
.B(n_7265),
.Y(n_7466)
);

NAND2xp5_ASAP7_75t_L g7467 ( 
.A(n_7366),
.B(n_7329),
.Y(n_7467)
);

NOR2x1p5_ASAP7_75t_L g7468 ( 
.A(n_7395),
.B(n_7230),
.Y(n_7468)
);

AND2x2_ASAP7_75t_L g7469 ( 
.A(n_7352),
.B(n_7224),
.Y(n_7469)
);

NOR2xp33_ASAP7_75t_SL g7470 ( 
.A(n_7431),
.B(n_7287),
.Y(n_7470)
);

INVx2_ASAP7_75t_SL g7471 ( 
.A(n_7424),
.Y(n_7471)
);

OAI22xp5_ASAP7_75t_L g7472 ( 
.A1(n_7399),
.A2(n_7297),
.B1(n_7246),
.B2(n_7220),
.Y(n_7472)
);

INVx3_ASAP7_75t_L g7473 ( 
.A(n_7398),
.Y(n_7473)
);

OR2x6_ASAP7_75t_L g7474 ( 
.A(n_7426),
.B(n_7322),
.Y(n_7474)
);

INVx1_ASAP7_75t_L g7475 ( 
.A(n_7378),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_7393),
.Y(n_7476)
);

AND2x4_ASAP7_75t_L g7477 ( 
.A(n_7418),
.B(n_7333),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_7420),
.Y(n_7478)
);

OR2x2_ASAP7_75t_L g7479 ( 
.A(n_7426),
.B(n_7323),
.Y(n_7479)
);

AND2x2_ASAP7_75t_L g7480 ( 
.A(n_7432),
.B(n_7224),
.Y(n_7480)
);

BUFx2_ASAP7_75t_L g7481 ( 
.A(n_7423),
.Y(n_7481)
);

NAND2x1p5_ASAP7_75t_L g7482 ( 
.A(n_7425),
.B(n_7401),
.Y(n_7482)
);

AND2x2_ASAP7_75t_L g7483 ( 
.A(n_7371),
.B(n_7294),
.Y(n_7483)
);

NAND2xp5_ASAP7_75t_L g7484 ( 
.A(n_7413),
.B(n_7326),
.Y(n_7484)
);

NAND2xp5_ASAP7_75t_L g7485 ( 
.A(n_7439),
.B(n_7331),
.Y(n_7485)
);

INVx1_ASAP7_75t_L g7486 ( 
.A(n_7353),
.Y(n_7486)
);

AND2x4_ASAP7_75t_L g7487 ( 
.A(n_7421),
.B(n_7261),
.Y(n_7487)
);

NAND2x1_ASAP7_75t_L g7488 ( 
.A(n_7394),
.B(n_7309),
.Y(n_7488)
);

AND2x2_ASAP7_75t_L g7489 ( 
.A(n_7400),
.B(n_7291),
.Y(n_7489)
);

INVx1_ASAP7_75t_L g7490 ( 
.A(n_7417),
.Y(n_7490)
);

AOI222xp33_ASAP7_75t_L g7491 ( 
.A1(n_7374),
.A2(n_7292),
.B1(n_7252),
.B2(n_7279),
.C1(n_7236),
.C2(n_7237),
.Y(n_7491)
);

NOR2xp33_ASAP7_75t_L g7492 ( 
.A(n_7383),
.B(n_7295),
.Y(n_7492)
);

NAND2xp5_ASAP7_75t_L g7493 ( 
.A(n_7402),
.B(n_7320),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_7373),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_7415),
.Y(n_7495)
);

INVx1_ASAP7_75t_L g7496 ( 
.A(n_7359),
.Y(n_7496)
);

NAND2xp5_ASAP7_75t_L g7497 ( 
.A(n_7363),
.B(n_7325),
.Y(n_7497)
);

OAI22xp33_ASAP7_75t_L g7498 ( 
.A1(n_7396),
.A2(n_7276),
.B1(n_7235),
.B2(n_7281),
.Y(n_7498)
);

OAI22xp5_ASAP7_75t_L g7499 ( 
.A1(n_7351),
.A2(n_7241),
.B1(n_7255),
.B2(n_7299),
.Y(n_7499)
);

AND2x2_ASAP7_75t_L g7500 ( 
.A(n_7365),
.B(n_7296),
.Y(n_7500)
);

INVx1_ASAP7_75t_L g7501 ( 
.A(n_7379),
.Y(n_7501)
);

INVx1_ASAP7_75t_L g7502 ( 
.A(n_7381),
.Y(n_7502)
);

AND2x2_ASAP7_75t_L g7503 ( 
.A(n_7436),
.B(n_246),
.Y(n_7503)
);

NAND2xp5_ASAP7_75t_SL g7504 ( 
.A(n_7358),
.B(n_246),
.Y(n_7504)
);

NAND2xp5_ASAP7_75t_L g7505 ( 
.A(n_7362),
.B(n_246),
.Y(n_7505)
);

AND2x4_ASAP7_75t_L g7506 ( 
.A(n_7405),
.B(n_247),
.Y(n_7506)
);

AOI21xp33_ASAP7_75t_SL g7507 ( 
.A1(n_7360),
.A2(n_247),
.B(n_248),
.Y(n_7507)
);

AND2x2_ASAP7_75t_L g7508 ( 
.A(n_7357),
.B(n_247),
.Y(n_7508)
);

INVx1_ASAP7_75t_L g7509 ( 
.A(n_7422),
.Y(n_7509)
);

NOR2xp67_ASAP7_75t_L g7510 ( 
.A(n_7377),
.B(n_247),
.Y(n_7510)
);

NOR2xp33_ASAP7_75t_L g7511 ( 
.A(n_7403),
.B(n_248),
.Y(n_7511)
);

OAI22xp33_ASAP7_75t_L g7512 ( 
.A1(n_7406),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_7512)
);

NAND2xp5_ASAP7_75t_L g7513 ( 
.A(n_7430),
.B(n_248),
.Y(n_7513)
);

INVx1_ASAP7_75t_SL g7514 ( 
.A(n_7355),
.Y(n_7514)
);

NOR3xp33_ASAP7_75t_L g7515 ( 
.A(n_7389),
.B(n_249),
.C(n_250),
.Y(n_7515)
);

INVx2_ASAP7_75t_L g7516 ( 
.A(n_7376),
.Y(n_7516)
);

HB1xp67_ASAP7_75t_L g7517 ( 
.A(n_7404),
.Y(n_7517)
);

NAND3xp33_ASAP7_75t_L g7518 ( 
.A(n_7429),
.B(n_250),
.C(n_251),
.Y(n_7518)
);

INVx1_ASAP7_75t_SL g7519 ( 
.A(n_7419),
.Y(n_7519)
);

AND2x4_ASAP7_75t_L g7520 ( 
.A(n_7440),
.B(n_250),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7428),
.Y(n_7521)
);

AO21x1_ASAP7_75t_L g7522 ( 
.A1(n_7407),
.A2(n_251),
.B(n_252),
.Y(n_7522)
);

NAND2x1_ASAP7_75t_L g7523 ( 
.A(n_7414),
.B(n_251),
.Y(n_7523)
);

NAND2xp5_ASAP7_75t_L g7524 ( 
.A(n_7408),
.B(n_7411),
.Y(n_7524)
);

INVxp67_ASAP7_75t_L g7525 ( 
.A(n_7416),
.Y(n_7525)
);

NOR2xp33_ASAP7_75t_L g7526 ( 
.A(n_7434),
.B(n_251),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_7412),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_7409),
.Y(n_7528)
);

AND2x2_ASAP7_75t_L g7529 ( 
.A(n_7392),
.B(n_252),
.Y(n_7529)
);

NAND2xp5_ASAP7_75t_L g7530 ( 
.A(n_7386),
.B(n_252),
.Y(n_7530)
);

HB1xp67_ASAP7_75t_L g7531 ( 
.A(n_7390),
.Y(n_7531)
);

NOR2xp33_ASAP7_75t_L g7532 ( 
.A(n_7375),
.B(n_253),
.Y(n_7532)
);

AND2x2_ASAP7_75t_L g7533 ( 
.A(n_7410),
.B(n_253),
.Y(n_7533)
);

AOI22xp5_ASAP7_75t_L g7534 ( 
.A1(n_7375),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_7534)
);

INVxp67_ASAP7_75t_L g7535 ( 
.A(n_7354),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7354),
.Y(n_7536)
);

AOI31xp33_ASAP7_75t_L g7537 ( 
.A1(n_7396),
.A2(n_256),
.A3(n_254),
.B(n_255),
.Y(n_7537)
);

AOI22x1_ASAP7_75t_L g7538 ( 
.A1(n_7364),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_7538)
);

AND2x2_ASAP7_75t_L g7539 ( 
.A(n_7410),
.B(n_254),
.Y(n_7539)
);

OAI22xp33_ASAP7_75t_L g7540 ( 
.A1(n_7375),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_7540)
);

NAND2xp5_ASAP7_75t_L g7541 ( 
.A(n_7438),
.B(n_256),
.Y(n_7541)
);

NAND2xp5_ASAP7_75t_L g7542 ( 
.A(n_7438),
.B(n_257),
.Y(n_7542)
);

CKINVDCx20_ASAP7_75t_R g7543 ( 
.A(n_7451),
.Y(n_7543)
);

INVx1_ASAP7_75t_L g7544 ( 
.A(n_7441),
.Y(n_7544)
);

OR2x2_ASAP7_75t_L g7545 ( 
.A(n_7444),
.B(n_257),
.Y(n_7545)
);

INVx1_ASAP7_75t_L g7546 ( 
.A(n_7443),
.Y(n_7546)
);

INVx2_ASAP7_75t_L g7547 ( 
.A(n_7446),
.Y(n_7547)
);

AND2x2_ASAP7_75t_L g7548 ( 
.A(n_7460),
.B(n_257),
.Y(n_7548)
);

AOI32xp33_ASAP7_75t_L g7549 ( 
.A1(n_7515),
.A2(n_260),
.A3(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7533),
.Y(n_7550)
);

NOR2xp33_ASAP7_75t_L g7551 ( 
.A(n_7473),
.B(n_258),
.Y(n_7551)
);

AND2x2_ASAP7_75t_L g7552 ( 
.A(n_7503),
.B(n_7539),
.Y(n_7552)
);

OAI21xp5_ASAP7_75t_L g7553 ( 
.A1(n_7535),
.A2(n_258),
.B(n_259),
.Y(n_7553)
);

OR2x2_ASAP7_75t_L g7554 ( 
.A(n_7471),
.B(n_7448),
.Y(n_7554)
);

OR2x2_ASAP7_75t_L g7555 ( 
.A(n_7449),
.B(n_258),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7454),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_7538),
.Y(n_7557)
);

OAI21xp5_ASAP7_75t_L g7558 ( 
.A1(n_7456),
.A2(n_259),
.B(n_260),
.Y(n_7558)
);

AOI22xp5_ASAP7_75t_L g7559 ( 
.A1(n_7442),
.A2(n_7470),
.B1(n_7466),
.B2(n_7528),
.Y(n_7559)
);

OAI22xp5_ASAP7_75t_L g7560 ( 
.A1(n_7536),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_7465),
.Y(n_7561)
);

OAI21xp33_ASAP7_75t_L g7562 ( 
.A1(n_7461),
.A2(n_261),
.B(n_262),
.Y(n_7562)
);

AND2x2_ASAP7_75t_L g7563 ( 
.A(n_7469),
.B(n_261),
.Y(n_7563)
);

INVxp67_ASAP7_75t_L g7564 ( 
.A(n_7532),
.Y(n_7564)
);

AOI21xp33_ASAP7_75t_L g7565 ( 
.A1(n_7459),
.A2(n_262),
.B(n_263),
.Y(n_7565)
);

NOR2xp33_ASAP7_75t_L g7566 ( 
.A(n_7504),
.B(n_7458),
.Y(n_7566)
);

INVx1_ASAP7_75t_L g7567 ( 
.A(n_7450),
.Y(n_7567)
);

AOI221xp5_ASAP7_75t_L g7568 ( 
.A1(n_7540),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_769),
.Y(n_7568)
);

NAND2xp5_ASAP7_75t_L g7569 ( 
.A(n_7520),
.B(n_263),
.Y(n_7569)
);

AND2x2_ASAP7_75t_L g7570 ( 
.A(n_7480),
.B(n_264),
.Y(n_7570)
);

AND2x2_ASAP7_75t_L g7571 ( 
.A(n_7508),
.B(n_264),
.Y(n_7571)
);

OR2x2_ASAP7_75t_L g7572 ( 
.A(n_7541),
.B(n_769),
.Y(n_7572)
);

INVx2_ASAP7_75t_L g7573 ( 
.A(n_7477),
.Y(n_7573)
);

NAND2xp5_ASAP7_75t_L g7574 ( 
.A(n_7520),
.B(n_769),
.Y(n_7574)
);

NAND2xp5_ASAP7_75t_L g7575 ( 
.A(n_7452),
.B(n_770),
.Y(n_7575)
);

NOR2xp33_ASAP7_75t_L g7576 ( 
.A(n_7537),
.B(n_770),
.Y(n_7576)
);

INVx5_ASAP7_75t_L g7577 ( 
.A(n_7477),
.Y(n_7577)
);

INVx2_ASAP7_75t_L g7578 ( 
.A(n_7482),
.Y(n_7578)
);

INVx2_ASAP7_75t_L g7579 ( 
.A(n_7453),
.Y(n_7579)
);

OAI21xp5_ASAP7_75t_L g7580 ( 
.A1(n_7518),
.A2(n_770),
.B(n_771),
.Y(n_7580)
);

NOR2xp33_ASAP7_75t_L g7581 ( 
.A(n_7542),
.B(n_771),
.Y(n_7581)
);

CKINVDCx20_ASAP7_75t_R g7582 ( 
.A(n_7464),
.Y(n_7582)
);

OAI32xp33_ASAP7_75t_L g7583 ( 
.A1(n_7505),
.A2(n_1070),
.A3(n_774),
.B1(n_772),
.B2(n_773),
.Y(n_7583)
);

OR2x2_ASAP7_75t_L g7584 ( 
.A(n_7479),
.B(n_1070),
.Y(n_7584)
);

OAI31xp33_ASAP7_75t_L g7585 ( 
.A1(n_7445),
.A2(n_774),
.A3(n_772),
.B(n_773),
.Y(n_7585)
);

NAND2x1p5_ASAP7_75t_L g7586 ( 
.A(n_7488),
.B(n_772),
.Y(n_7586)
);

AOI22xp5_ASAP7_75t_L g7587 ( 
.A1(n_7526),
.A2(n_1059),
.B1(n_777),
.B2(n_775),
.Y(n_7587)
);

OAI22xp33_ASAP7_75t_L g7588 ( 
.A1(n_7467),
.A2(n_7513),
.B1(n_7530),
.B2(n_7474),
.Y(n_7588)
);

OAI21xp5_ASAP7_75t_SL g7589 ( 
.A1(n_7491),
.A2(n_775),
.B(n_776),
.Y(n_7589)
);

INVx2_ASAP7_75t_SL g7590 ( 
.A(n_7463),
.Y(n_7590)
);

INVx1_ASAP7_75t_L g7591 ( 
.A(n_7529),
.Y(n_7591)
);

INVx1_ASAP7_75t_L g7592 ( 
.A(n_7523),
.Y(n_7592)
);

OAI221xp5_ASAP7_75t_L g7593 ( 
.A1(n_7534),
.A2(n_778),
.B1(n_775),
.B2(n_777),
.C(n_779),
.Y(n_7593)
);

AOI22xp5_ASAP7_75t_L g7594 ( 
.A1(n_7511),
.A2(n_780),
.B1(n_778),
.B2(n_779),
.Y(n_7594)
);

NAND2xp5_ASAP7_75t_SL g7595 ( 
.A(n_7512),
.B(n_778),
.Y(n_7595)
);

AND2x2_ASAP7_75t_L g7596 ( 
.A(n_7489),
.B(n_781),
.Y(n_7596)
);

INVx1_ASAP7_75t_SL g7597 ( 
.A(n_7554),
.Y(n_7597)
);

AOI22xp5_ASAP7_75t_L g7598 ( 
.A1(n_7543),
.A2(n_7455),
.B1(n_7462),
.B2(n_7506),
.Y(n_7598)
);

AND2x2_ASAP7_75t_L g7599 ( 
.A(n_7573),
.B(n_7547),
.Y(n_7599)
);

INVx2_ASAP7_75t_SL g7600 ( 
.A(n_7577),
.Y(n_7600)
);

AOI211xp5_ASAP7_75t_L g7601 ( 
.A1(n_7565),
.A2(n_7507),
.B(n_7472),
.C(n_7498),
.Y(n_7601)
);

INVx2_ASAP7_75t_L g7602 ( 
.A(n_7577),
.Y(n_7602)
);

NAND2xp5_ASAP7_75t_SL g7603 ( 
.A(n_7544),
.B(n_7510),
.Y(n_7603)
);

INVx1_ASAP7_75t_L g7604 ( 
.A(n_7563),
.Y(n_7604)
);

INVx2_ASAP7_75t_L g7605 ( 
.A(n_7577),
.Y(n_7605)
);

INVxp67_ASAP7_75t_L g7606 ( 
.A(n_7570),
.Y(n_7606)
);

INVx1_ASAP7_75t_L g7607 ( 
.A(n_7569),
.Y(n_7607)
);

INVx1_ASAP7_75t_L g7608 ( 
.A(n_7546),
.Y(n_7608)
);

NAND2xp5_ASAP7_75t_L g7609 ( 
.A(n_7548),
.B(n_7500),
.Y(n_7609)
);

OAI21xp5_ASAP7_75t_SL g7610 ( 
.A1(n_7559),
.A2(n_7589),
.B(n_7549),
.Y(n_7610)
);

OR2x2_ASAP7_75t_L g7611 ( 
.A(n_7590),
.B(n_7474),
.Y(n_7611)
);

INVx2_ASAP7_75t_L g7612 ( 
.A(n_7578),
.Y(n_7612)
);

INVxp67_ASAP7_75t_L g7613 ( 
.A(n_7551),
.Y(n_7613)
);

INVx1_ASAP7_75t_L g7614 ( 
.A(n_7596),
.Y(n_7614)
);

INVx1_ASAP7_75t_L g7615 ( 
.A(n_7574),
.Y(n_7615)
);

INVxp67_ASAP7_75t_L g7616 ( 
.A(n_7575),
.Y(n_7616)
);

NAND2xp5_ASAP7_75t_L g7617 ( 
.A(n_7571),
.B(n_7483),
.Y(n_7617)
);

NAND2xp5_ASAP7_75t_L g7618 ( 
.A(n_7561),
.B(n_7478),
.Y(n_7618)
);

O2A1O1Ixp33_ASAP7_75t_L g7619 ( 
.A1(n_7583),
.A2(n_7517),
.B(n_7499),
.C(n_7531),
.Y(n_7619)
);

INVx1_ASAP7_75t_L g7620 ( 
.A(n_7555),
.Y(n_7620)
);

AOI21xp33_ASAP7_75t_L g7621 ( 
.A1(n_7560),
.A2(n_7527),
.B(n_7485),
.Y(n_7621)
);

INVx2_ASAP7_75t_L g7622 ( 
.A(n_7545),
.Y(n_7622)
);

OR2x2_ASAP7_75t_L g7623 ( 
.A(n_7556),
.B(n_7494),
.Y(n_7623)
);

AOI21xp5_ASAP7_75t_L g7624 ( 
.A1(n_7595),
.A2(n_7484),
.B(n_7493),
.Y(n_7624)
);

O2A1O1Ixp33_ASAP7_75t_L g7625 ( 
.A1(n_7562),
.A2(n_7516),
.B(n_7501),
.C(n_7502),
.Y(n_7625)
);

INVx1_ASAP7_75t_L g7626 ( 
.A(n_7586),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_7584),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7552),
.Y(n_7628)
);

OAI21xp33_ASAP7_75t_L g7629 ( 
.A1(n_7567),
.A2(n_7492),
.B(n_7497),
.Y(n_7629)
);

AND2x2_ASAP7_75t_L g7630 ( 
.A(n_7579),
.B(n_7468),
.Y(n_7630)
);

NAND2xp5_ASAP7_75t_SL g7631 ( 
.A(n_7585),
.B(n_7487),
.Y(n_7631)
);

NOR2xp33_ASAP7_75t_L g7632 ( 
.A(n_7582),
.B(n_7522),
.Y(n_7632)
);

NAND2xp5_ASAP7_75t_L g7633 ( 
.A(n_7576),
.B(n_7495),
.Y(n_7633)
);

INVx2_ASAP7_75t_SL g7634 ( 
.A(n_7592),
.Y(n_7634)
);

AOI322xp5_ASAP7_75t_L g7635 ( 
.A1(n_7581),
.A2(n_7514),
.A3(n_7519),
.B1(n_7486),
.B2(n_7490),
.C1(n_7457),
.C2(n_7447),
.Y(n_7635)
);

INVxp67_ASAP7_75t_SL g7636 ( 
.A(n_7566),
.Y(n_7636)
);

INVx1_ASAP7_75t_L g7637 ( 
.A(n_7572),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_7557),
.Y(n_7638)
);

A2O1A1Ixp33_ASAP7_75t_L g7639 ( 
.A1(n_7568),
.A2(n_7553),
.B(n_7558),
.C(n_7594),
.Y(n_7639)
);

AOI22xp33_ASAP7_75t_SL g7640 ( 
.A1(n_7550),
.A2(n_7481),
.B1(n_7521),
.B2(n_7509),
.Y(n_7640)
);

OAI21xp5_ASAP7_75t_L g7641 ( 
.A1(n_7580),
.A2(n_7524),
.B(n_7525),
.Y(n_7641)
);

INVx1_ASAP7_75t_L g7642 ( 
.A(n_7591),
.Y(n_7642)
);

INVx1_ASAP7_75t_L g7643 ( 
.A(n_7587),
.Y(n_7643)
);

INVx1_ASAP7_75t_L g7644 ( 
.A(n_7593),
.Y(n_7644)
);

NOR2xp33_ASAP7_75t_L g7645 ( 
.A(n_7588),
.B(n_7476),
.Y(n_7645)
);

OAI21xp5_ASAP7_75t_SL g7646 ( 
.A1(n_7564),
.A2(n_7496),
.B(n_7475),
.Y(n_7646)
);

INVx1_ASAP7_75t_SL g7647 ( 
.A(n_7554),
.Y(n_7647)
);

OAI221xp5_ASAP7_75t_L g7648 ( 
.A1(n_7585),
.A2(n_783),
.B1(n_781),
.B2(n_782),
.C(n_784),
.Y(n_7648)
);

O2A1O1Ixp33_ASAP7_75t_L g7649 ( 
.A1(n_7583),
.A2(n_783),
.B(n_781),
.C(n_782),
.Y(n_7649)
);

NAND2xp5_ASAP7_75t_L g7650 ( 
.A(n_7577),
.B(n_782),
.Y(n_7650)
);

INVx1_ASAP7_75t_L g7651 ( 
.A(n_7554),
.Y(n_7651)
);

OAI21xp33_ASAP7_75t_L g7652 ( 
.A1(n_7544),
.A2(n_783),
.B(n_784),
.Y(n_7652)
);

AOI21xp33_ASAP7_75t_L g7653 ( 
.A1(n_7554),
.A2(n_784),
.B(n_785),
.Y(n_7653)
);

INVxp67_ASAP7_75t_L g7654 ( 
.A(n_7554),
.Y(n_7654)
);

INVx1_ASAP7_75t_L g7655 ( 
.A(n_7599),
.Y(n_7655)
);

NOR3xp33_ASAP7_75t_L g7656 ( 
.A(n_7654),
.B(n_1059),
.C(n_785),
.Y(n_7656)
);

AOI21xp33_ASAP7_75t_L g7657 ( 
.A1(n_7597),
.A2(n_786),
.B(n_787),
.Y(n_7657)
);

OAI21xp33_ASAP7_75t_L g7658 ( 
.A1(n_7647),
.A2(n_786),
.B(n_787),
.Y(n_7658)
);

OAI22xp5_ASAP7_75t_L g7659 ( 
.A1(n_7612),
.A2(n_788),
.B1(n_786),
.B2(n_787),
.Y(n_7659)
);

OAI321xp33_ASAP7_75t_L g7660 ( 
.A1(n_7651),
.A2(n_790),
.A3(n_792),
.B1(n_788),
.B2(n_789),
.C(n_791),
.Y(n_7660)
);

INVx1_ASAP7_75t_L g7661 ( 
.A(n_7650),
.Y(n_7661)
);

NOR2x1_ASAP7_75t_L g7662 ( 
.A(n_7611),
.B(n_789),
.Y(n_7662)
);

AOI22xp5_ASAP7_75t_L g7663 ( 
.A1(n_7634),
.A2(n_1055),
.B1(n_792),
.B2(n_790),
.Y(n_7663)
);

A2O1A1Ixp33_ASAP7_75t_L g7664 ( 
.A1(n_7619),
.A2(n_793),
.B(n_791),
.C(n_792),
.Y(n_7664)
);

INVx1_ASAP7_75t_L g7665 ( 
.A(n_7609),
.Y(n_7665)
);

AOI21xp33_ASAP7_75t_L g7666 ( 
.A1(n_7649),
.A2(n_794),
.B(n_795),
.Y(n_7666)
);

O2A1O1Ixp5_ASAP7_75t_L g7667 ( 
.A1(n_7631),
.A2(n_796),
.B(n_794),
.C(n_795),
.Y(n_7667)
);

OAI22xp5_ASAP7_75t_L g7668 ( 
.A1(n_7598),
.A2(n_798),
.B1(n_796),
.B2(n_797),
.Y(n_7668)
);

AOI22xp33_ASAP7_75t_SL g7669 ( 
.A1(n_7636),
.A2(n_7608),
.B1(n_7638),
.B2(n_7630),
.Y(n_7669)
);

NAND2xp5_ASAP7_75t_L g7670 ( 
.A(n_7600),
.B(n_797),
.Y(n_7670)
);

OAI211xp5_ASAP7_75t_L g7671 ( 
.A1(n_7653),
.A2(n_800),
.B(n_798),
.C(n_799),
.Y(n_7671)
);

INVxp33_ASAP7_75t_L g7672 ( 
.A(n_7645),
.Y(n_7672)
);

O2A1O1Ixp33_ASAP7_75t_L g7673 ( 
.A1(n_7618),
.A2(n_800),
.B(n_798),
.C(n_799),
.Y(n_7673)
);

AOI222xp33_ASAP7_75t_L g7674 ( 
.A1(n_7652),
.A2(n_801),
.B1(n_803),
.B2(n_799),
.C1(n_800),
.C2(n_802),
.Y(n_7674)
);

INVx1_ASAP7_75t_L g7675 ( 
.A(n_7617),
.Y(n_7675)
);

AOI31xp33_ASAP7_75t_L g7676 ( 
.A1(n_7601),
.A2(n_803),
.A3(n_801),
.B(n_802),
.Y(n_7676)
);

A2O1A1Ixp33_ASAP7_75t_L g7677 ( 
.A1(n_7625),
.A2(n_803),
.B(n_801),
.C(n_802),
.Y(n_7677)
);

AOI211xp5_ASAP7_75t_L g7678 ( 
.A1(n_7648),
.A2(n_806),
.B(n_804),
.C(n_805),
.Y(n_7678)
);

AOI21xp5_ASAP7_75t_L g7679 ( 
.A1(n_7603),
.A2(n_804),
.B(n_805),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_7623),
.Y(n_7680)
);

O2A1O1Ixp33_ASAP7_75t_L g7681 ( 
.A1(n_7621),
.A2(n_807),
.B(n_805),
.C(n_806),
.Y(n_7681)
);

OAI21xp33_ASAP7_75t_L g7682 ( 
.A1(n_7629),
.A2(n_806),
.B(n_807),
.Y(n_7682)
);

AOI211x1_ASAP7_75t_L g7683 ( 
.A1(n_7624),
.A2(n_809),
.B(n_807),
.C(n_808),
.Y(n_7683)
);

AOI322xp5_ASAP7_75t_L g7684 ( 
.A1(n_7632),
.A2(n_808),
.A3(n_809),
.B1(n_810),
.B2(n_811),
.C1(n_812),
.C2(n_813),
.Y(n_7684)
);

AOI21xp33_ASAP7_75t_L g7685 ( 
.A1(n_7602),
.A2(n_808),
.B(n_810),
.Y(n_7685)
);

AOI32xp33_ASAP7_75t_L g7686 ( 
.A1(n_7644),
.A2(n_812),
.A3(n_810),
.B1(n_811),
.B2(n_813),
.Y(n_7686)
);

AOI221xp5_ASAP7_75t_L g7687 ( 
.A1(n_7610),
.A2(n_814),
.B1(n_811),
.B2(n_813),
.C(n_815),
.Y(n_7687)
);

OR2x2_ASAP7_75t_L g7688 ( 
.A(n_7605),
.B(n_814),
.Y(n_7688)
);

AOI221xp5_ASAP7_75t_L g7689 ( 
.A1(n_7628),
.A2(n_816),
.B1(n_814),
.B2(n_815),
.C(n_817),
.Y(n_7689)
);

NOR2xp33_ASAP7_75t_L g7690 ( 
.A(n_7606),
.B(n_815),
.Y(n_7690)
);

INVx1_ASAP7_75t_SL g7691 ( 
.A(n_7620),
.Y(n_7691)
);

INVx1_ASAP7_75t_L g7692 ( 
.A(n_7604),
.Y(n_7692)
);

AOI221x1_ASAP7_75t_L g7693 ( 
.A1(n_7627),
.A2(n_818),
.B1(n_816),
.B2(n_817),
.C(n_819),
.Y(n_7693)
);

INVx1_ASAP7_75t_L g7694 ( 
.A(n_7598),
.Y(n_7694)
);

AOI211xp5_ASAP7_75t_SL g7695 ( 
.A1(n_7613),
.A2(n_820),
.B(n_818),
.C(n_819),
.Y(n_7695)
);

NAND2xp33_ASAP7_75t_R g7696 ( 
.A(n_7626),
.B(n_818),
.Y(n_7696)
);

INVx1_ASAP7_75t_L g7697 ( 
.A(n_7614),
.Y(n_7697)
);

NAND2xp5_ASAP7_75t_L g7698 ( 
.A(n_7655),
.B(n_7622),
.Y(n_7698)
);

OAI21xp5_ASAP7_75t_L g7699 ( 
.A1(n_7664),
.A2(n_7639),
.B(n_7635),
.Y(n_7699)
);

NAND2xp5_ASAP7_75t_L g7700 ( 
.A(n_7684),
.B(n_7642),
.Y(n_7700)
);

OAI21xp33_ASAP7_75t_SL g7701 ( 
.A1(n_7665),
.A2(n_7633),
.B(n_7643),
.Y(n_7701)
);

AOI322xp5_ASAP7_75t_L g7702 ( 
.A1(n_7691),
.A2(n_7637),
.A3(n_7607),
.B1(n_7615),
.B2(n_7640),
.C1(n_7616),
.C2(n_7646),
.Y(n_7702)
);

AOI221xp5_ASAP7_75t_L g7703 ( 
.A1(n_7685),
.A2(n_7641),
.B1(n_821),
.B2(n_819),
.C(n_820),
.Y(n_7703)
);

OAI31xp33_ASAP7_75t_L g7704 ( 
.A1(n_7671),
.A2(n_822),
.A3(n_820),
.B(n_821),
.Y(n_7704)
);

AOI322xp5_ASAP7_75t_L g7705 ( 
.A1(n_7690),
.A2(n_822),
.A3(n_823),
.B1(n_824),
.B2(n_825),
.C1(n_826),
.C2(n_827),
.Y(n_7705)
);

AOI21xp5_ASAP7_75t_L g7706 ( 
.A1(n_7670),
.A2(n_823),
.B(n_824),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_7688),
.Y(n_7707)
);

AOI22xp5_ASAP7_75t_L g7708 ( 
.A1(n_7675),
.A2(n_7694),
.B1(n_7680),
.B2(n_7692),
.Y(n_7708)
);

OR2x2_ASAP7_75t_L g7709 ( 
.A(n_7668),
.B(n_825),
.Y(n_7709)
);

OA22x2_ASAP7_75t_L g7710 ( 
.A1(n_7697),
.A2(n_827),
.B1(n_825),
.B2(n_826),
.Y(n_7710)
);

AOI322xp5_ASAP7_75t_L g7711 ( 
.A1(n_7669),
.A2(n_827),
.A3(n_828),
.B1(n_829),
.B2(n_830),
.C1(n_831),
.C2(n_832),
.Y(n_7711)
);

NAND2xp5_ASAP7_75t_L g7712 ( 
.A(n_7687),
.B(n_7689),
.Y(n_7712)
);

AOI221xp5_ASAP7_75t_L g7713 ( 
.A1(n_7676),
.A2(n_830),
.B1(n_828),
.B2(n_829),
.C(n_831),
.Y(n_7713)
);

OAI221xp5_ASAP7_75t_L g7714 ( 
.A1(n_7686),
.A2(n_831),
.B1(n_828),
.B2(n_830),
.C(n_832),
.Y(n_7714)
);

OAI221xp5_ASAP7_75t_L g7715 ( 
.A1(n_7658),
.A2(n_834),
.B1(n_832),
.B2(n_833),
.C(n_835),
.Y(n_7715)
);

NOR4xp25_ASAP7_75t_SL g7716 ( 
.A(n_7696),
.B(n_835),
.C(n_833),
.D(n_834),
.Y(n_7716)
);

AOI22xp5_ASAP7_75t_L g7717 ( 
.A1(n_7672),
.A2(n_835),
.B1(n_833),
.B2(n_834),
.Y(n_7717)
);

AOI221xp5_ASAP7_75t_L g7718 ( 
.A1(n_7657),
.A2(n_838),
.B1(n_836),
.B2(n_837),
.C(n_839),
.Y(n_7718)
);

AOI211xp5_ASAP7_75t_L g7719 ( 
.A1(n_7666),
.A2(n_838),
.B(n_836),
.C(n_837),
.Y(n_7719)
);

NOR2x1_ASAP7_75t_L g7720 ( 
.A(n_7662),
.B(n_836),
.Y(n_7720)
);

AND4x1_ASAP7_75t_L g7721 ( 
.A(n_7695),
.B(n_841),
.C(n_838),
.D(n_839),
.Y(n_7721)
);

AOI222xp33_ASAP7_75t_L g7722 ( 
.A1(n_7682),
.A2(n_843),
.B1(n_845),
.B2(n_841),
.C1(n_842),
.C2(n_844),
.Y(n_7722)
);

NOR3xp33_ASAP7_75t_L g7723 ( 
.A(n_7660),
.B(n_841),
.C(n_842),
.Y(n_7723)
);

AOI211xp5_ASAP7_75t_L g7724 ( 
.A1(n_7659),
.A2(n_844),
.B(n_842),
.C(n_843),
.Y(n_7724)
);

NAND2xp5_ASAP7_75t_SL g7725 ( 
.A(n_7678),
.B(n_843),
.Y(n_7725)
);

INVxp67_ASAP7_75t_SL g7726 ( 
.A(n_7681),
.Y(n_7726)
);

INVx1_ASAP7_75t_L g7727 ( 
.A(n_7663),
.Y(n_7727)
);

AOI21xp5_ASAP7_75t_L g7728 ( 
.A1(n_7677),
.A2(n_844),
.B(n_845),
.Y(n_7728)
);

AOI31xp33_ASAP7_75t_L g7729 ( 
.A1(n_7674),
.A2(n_847),
.A3(n_845),
.B(n_846),
.Y(n_7729)
);

AOI322xp5_ASAP7_75t_L g7730 ( 
.A1(n_7656),
.A2(n_846),
.A3(n_847),
.B1(n_848),
.B2(n_849),
.C1(n_850),
.C2(n_851),
.Y(n_7730)
);

NAND2xp5_ASAP7_75t_SL g7731 ( 
.A(n_7667),
.B(n_846),
.Y(n_7731)
);

OAI22xp5_ASAP7_75t_L g7732 ( 
.A1(n_7661),
.A2(n_850),
.B1(n_848),
.B2(n_849),
.Y(n_7732)
);

OAI22xp5_ASAP7_75t_L g7733 ( 
.A1(n_7683),
.A2(n_850),
.B1(n_848),
.B2(n_849),
.Y(n_7733)
);

NAND3xp33_ASAP7_75t_L g7734 ( 
.A(n_7673),
.B(n_7679),
.C(n_7693),
.Y(n_7734)
);

OAI322xp33_ASAP7_75t_SL g7735 ( 
.A1(n_7655),
.A2(n_851),
.A3(n_852),
.B1(n_853),
.B2(n_854),
.C1(n_855),
.C2(n_856),
.Y(n_7735)
);

NAND2xp5_ASAP7_75t_L g7736 ( 
.A(n_7655),
.B(n_852),
.Y(n_7736)
);

NAND2xp5_ASAP7_75t_L g7737 ( 
.A(n_7655),
.B(n_852),
.Y(n_7737)
);

XNOR2x1_ASAP7_75t_L g7738 ( 
.A(n_7662),
.B(n_853),
.Y(n_7738)
);

INVx2_ASAP7_75t_L g7739 ( 
.A(n_7655),
.Y(n_7739)
);

NOR2xp67_ASAP7_75t_L g7740 ( 
.A(n_7655),
.B(n_854),
.Y(n_7740)
);

INVx1_ASAP7_75t_L g7741 ( 
.A(n_7655),
.Y(n_7741)
);

AOI22xp33_ASAP7_75t_SL g7742 ( 
.A1(n_7655),
.A2(n_857),
.B1(n_855),
.B2(n_856),
.Y(n_7742)
);

AOI221xp5_ASAP7_75t_L g7743 ( 
.A1(n_7685),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.C(n_860),
.Y(n_7743)
);

NAND4xp25_ASAP7_75t_L g7744 ( 
.A(n_7655),
.B(n_859),
.C(n_857),
.D(n_858),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_7655),
.Y(n_7745)
);

INVx1_ASAP7_75t_L g7746 ( 
.A(n_7710),
.Y(n_7746)
);

NAND2xp5_ASAP7_75t_L g7747 ( 
.A(n_7711),
.B(n_858),
.Y(n_7747)
);

AND2x2_ASAP7_75t_L g7748 ( 
.A(n_7739),
.B(n_859),
.Y(n_7748)
);

NAND2xp5_ASAP7_75t_L g7749 ( 
.A(n_7705),
.B(n_860),
.Y(n_7749)
);

OAI32xp33_ASAP7_75t_L g7750 ( 
.A1(n_7701),
.A2(n_862),
.A3(n_860),
.B1(n_861),
.B2(n_863),
.Y(n_7750)
);

INVx1_ASAP7_75t_L g7751 ( 
.A(n_7736),
.Y(n_7751)
);

INVx1_ASAP7_75t_L g7752 ( 
.A(n_7737),
.Y(n_7752)
);

INVx1_ASAP7_75t_L g7753 ( 
.A(n_7698),
.Y(n_7753)
);

AND2x2_ASAP7_75t_L g7754 ( 
.A(n_7741),
.B(n_861),
.Y(n_7754)
);

NAND2xp5_ASAP7_75t_L g7755 ( 
.A(n_7742),
.B(n_7745),
.Y(n_7755)
);

AND2x2_ASAP7_75t_L g7756 ( 
.A(n_7708),
.B(n_862),
.Y(n_7756)
);

NAND2xp5_ASAP7_75t_L g7757 ( 
.A(n_7740),
.B(n_7730),
.Y(n_7757)
);

NOR2x1_ASAP7_75t_L g7758 ( 
.A(n_7734),
.B(n_862),
.Y(n_7758)
);

INVx1_ASAP7_75t_SL g7759 ( 
.A(n_7709),
.Y(n_7759)
);

OR2x2_ASAP7_75t_L g7760 ( 
.A(n_7744),
.B(n_863),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_7717),
.Y(n_7761)
);

INVxp67_ASAP7_75t_L g7762 ( 
.A(n_7715),
.Y(n_7762)
);

NAND2xp5_ASAP7_75t_L g7763 ( 
.A(n_7722),
.B(n_863),
.Y(n_7763)
);

NAND2xp5_ASAP7_75t_SL g7764 ( 
.A(n_7703),
.B(n_864),
.Y(n_7764)
);

NAND2xp5_ASAP7_75t_SL g7765 ( 
.A(n_7704),
.B(n_864),
.Y(n_7765)
);

AND2x2_ASAP7_75t_L g7766 ( 
.A(n_7707),
.B(n_864),
.Y(n_7766)
);

NAND2xp5_ASAP7_75t_L g7767 ( 
.A(n_7743),
.B(n_865),
.Y(n_7767)
);

HB1xp67_ASAP7_75t_L g7768 ( 
.A(n_7699),
.Y(n_7768)
);

INVxp67_ASAP7_75t_SL g7769 ( 
.A(n_7700),
.Y(n_7769)
);

OAI22xp33_ASAP7_75t_L g7770 ( 
.A1(n_7729),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_7732),
.Y(n_7771)
);

INVx2_ASAP7_75t_L g7772 ( 
.A(n_7738),
.Y(n_7772)
);

INVx1_ASAP7_75t_L g7773 ( 
.A(n_7726),
.Y(n_7773)
);

INVx1_ASAP7_75t_L g7774 ( 
.A(n_7720),
.Y(n_7774)
);

INVx1_ASAP7_75t_L g7775 ( 
.A(n_7721),
.Y(n_7775)
);

NAND2xp5_ASAP7_75t_L g7776 ( 
.A(n_7718),
.B(n_865),
.Y(n_7776)
);

INVx1_ASAP7_75t_L g7777 ( 
.A(n_7731),
.Y(n_7777)
);

INVx1_ASAP7_75t_L g7778 ( 
.A(n_7733),
.Y(n_7778)
);

NOR2xp33_ASAP7_75t_L g7779 ( 
.A(n_7714),
.B(n_866),
.Y(n_7779)
);

NAND2xp5_ASAP7_75t_L g7780 ( 
.A(n_7713),
.B(n_867),
.Y(n_7780)
);

OR2x2_ASAP7_75t_L g7781 ( 
.A(n_7712),
.B(n_867),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_7719),
.Y(n_7782)
);

OAI221xp5_ASAP7_75t_L g7783 ( 
.A1(n_7724),
.A2(n_870),
.B1(n_868),
.B2(n_869),
.C(n_871),
.Y(n_7783)
);

INVx1_ASAP7_75t_L g7784 ( 
.A(n_7727),
.Y(n_7784)
);

INVx1_ASAP7_75t_L g7785 ( 
.A(n_7723),
.Y(n_7785)
);

NOR2xp33_ASAP7_75t_L g7786 ( 
.A(n_7725),
.B(n_869),
.Y(n_7786)
);

INVx1_ASAP7_75t_L g7787 ( 
.A(n_7706),
.Y(n_7787)
);

NOR2xp33_ASAP7_75t_L g7788 ( 
.A(n_7728),
.B(n_870),
.Y(n_7788)
);

INVx2_ASAP7_75t_L g7789 ( 
.A(n_7702),
.Y(n_7789)
);

INVx1_ASAP7_75t_SL g7790 ( 
.A(n_7753),
.Y(n_7790)
);

A2O1A1Ixp33_ASAP7_75t_L g7791 ( 
.A1(n_7779),
.A2(n_7735),
.B(n_7716),
.C(n_873),
.Y(n_7791)
);

OAI21xp33_ASAP7_75t_SL g7792 ( 
.A1(n_7769),
.A2(n_871),
.B(n_872),
.Y(n_7792)
);

AOI221xp5_ASAP7_75t_SL g7793 ( 
.A1(n_7783),
.A2(n_874),
.B1(n_871),
.B2(n_872),
.C(n_875),
.Y(n_7793)
);

AOI222xp33_ASAP7_75t_L g7794 ( 
.A1(n_7773),
.A2(n_872),
.B1(n_874),
.B2(n_875),
.C1(n_876),
.C2(n_877),
.Y(n_7794)
);

O2A1O1Ixp33_ASAP7_75t_L g7795 ( 
.A1(n_7768),
.A2(n_877),
.B(n_875),
.C(n_876),
.Y(n_7795)
);

AND2x2_ASAP7_75t_L g7796 ( 
.A(n_7754),
.B(n_877),
.Y(n_7796)
);

INVx1_ASAP7_75t_L g7797 ( 
.A(n_7789),
.Y(n_7797)
);

INVxp33_ASAP7_75t_L g7798 ( 
.A(n_7766),
.Y(n_7798)
);

AOI21xp5_ASAP7_75t_L g7799 ( 
.A1(n_7747),
.A2(n_7749),
.B(n_7763),
.Y(n_7799)
);

O2A1O1Ixp33_ASAP7_75t_L g7800 ( 
.A1(n_7784),
.A2(n_880),
.B(n_878),
.C(n_879),
.Y(n_7800)
);

NAND3xp33_ASAP7_75t_L g7801 ( 
.A(n_7788),
.B(n_878),
.C(n_879),
.Y(n_7801)
);

NAND4xp25_ASAP7_75t_L g7802 ( 
.A(n_7762),
.B(n_880),
.C(n_878),
.D(n_879),
.Y(n_7802)
);

AOI22x1_ASAP7_75t_SL g7803 ( 
.A1(n_7771),
.A2(n_882),
.B1(n_880),
.B2(n_881),
.Y(n_7803)
);

AOI221xp5_ASAP7_75t_L g7804 ( 
.A1(n_7770),
.A2(n_1055),
.B1(n_883),
.B2(n_881),
.C(n_882),
.Y(n_7804)
);

AOI221xp5_ASAP7_75t_L g7805 ( 
.A1(n_7750),
.A2(n_1054),
.B1(n_884),
.B2(n_881),
.C(n_883),
.Y(n_7805)
);

NAND2xp5_ASAP7_75t_L g7806 ( 
.A(n_7748),
.B(n_883),
.Y(n_7806)
);

AOI221xp5_ASAP7_75t_L g7807 ( 
.A1(n_7786),
.A2(n_1054),
.B1(n_886),
.B2(n_884),
.C(n_885),
.Y(n_7807)
);

NOR3xp33_ASAP7_75t_L g7808 ( 
.A(n_7755),
.B(n_884),
.C(n_885),
.Y(n_7808)
);

AOI221xp5_ASAP7_75t_L g7809 ( 
.A1(n_7778),
.A2(n_1054),
.B1(n_888),
.B2(n_886),
.C(n_887),
.Y(n_7809)
);

AOI22xp33_ASAP7_75t_L g7810 ( 
.A1(n_7756),
.A2(n_888),
.B1(n_886),
.B2(n_887),
.Y(n_7810)
);

NAND2xp5_ASAP7_75t_L g7811 ( 
.A(n_7758),
.B(n_887),
.Y(n_7811)
);

INVx1_ASAP7_75t_L g7812 ( 
.A(n_7760),
.Y(n_7812)
);

AOI211xp5_ASAP7_75t_L g7813 ( 
.A1(n_7780),
.A2(n_891),
.B(n_889),
.C(n_890),
.Y(n_7813)
);

O2A1O1Ixp33_ASAP7_75t_L g7814 ( 
.A1(n_7776),
.A2(n_891),
.B(n_889),
.C(n_890),
.Y(n_7814)
);

AOI322xp5_ASAP7_75t_L g7815 ( 
.A1(n_7759),
.A2(n_892),
.A3(n_893),
.B1(n_894),
.B2(n_895),
.C1(n_896),
.C2(n_897),
.Y(n_7815)
);

NAND4xp25_ASAP7_75t_SL g7816 ( 
.A(n_7759),
.B(n_7767),
.C(n_7785),
.D(n_7781),
.Y(n_7816)
);

NOR2xp33_ASAP7_75t_L g7817 ( 
.A(n_7746),
.B(n_892),
.Y(n_7817)
);

A2O1A1Ixp33_ASAP7_75t_L g7818 ( 
.A1(n_7787),
.A2(n_897),
.B(n_893),
.C(n_895),
.Y(n_7818)
);

AND4x1_ASAP7_75t_L g7819 ( 
.A(n_7761),
.B(n_897),
.C(n_893),
.D(n_895),
.Y(n_7819)
);

OAI211xp5_ASAP7_75t_L g7820 ( 
.A1(n_7765),
.A2(n_900),
.B(n_898),
.C(n_899),
.Y(n_7820)
);

AOI221xp5_ASAP7_75t_L g7821 ( 
.A1(n_7764),
.A2(n_1053),
.B1(n_901),
.B2(n_898),
.C(n_899),
.Y(n_7821)
);

NAND3xp33_ASAP7_75t_L g7822 ( 
.A(n_7797),
.B(n_7775),
.C(n_7777),
.Y(n_7822)
);

NAND2xp5_ASAP7_75t_SL g7823 ( 
.A(n_7813),
.B(n_7782),
.Y(n_7823)
);

AND3x4_ASAP7_75t_L g7824 ( 
.A(n_7819),
.B(n_7772),
.C(n_7752),
.Y(n_7824)
);

OAI21xp5_ASAP7_75t_L g7825 ( 
.A1(n_7790),
.A2(n_7757),
.B(n_7751),
.Y(n_7825)
);

INVx2_ASAP7_75t_L g7826 ( 
.A(n_7812),
.Y(n_7826)
);

AND2x4_ASAP7_75t_L g7827 ( 
.A(n_7796),
.B(n_7774),
.Y(n_7827)
);

OAI22xp5_ASAP7_75t_L g7828 ( 
.A1(n_7806),
.A2(n_902),
.B1(n_898),
.B2(n_901),
.Y(n_7828)
);

NAND2xp5_ASAP7_75t_L g7829 ( 
.A(n_7809),
.B(n_901),
.Y(n_7829)
);

NAND2xp5_ASAP7_75t_L g7830 ( 
.A(n_7794),
.B(n_902),
.Y(n_7830)
);

AOI22xp5_ASAP7_75t_L g7831 ( 
.A1(n_7816),
.A2(n_905),
.B1(n_903),
.B2(n_904),
.Y(n_7831)
);

INVx1_ASAP7_75t_L g7832 ( 
.A(n_7803),
.Y(n_7832)
);

AOI21xp5_ASAP7_75t_L g7833 ( 
.A1(n_7795),
.A2(n_903),
.B(n_904),
.Y(n_7833)
);

INVxp67_ASAP7_75t_L g7834 ( 
.A(n_7817),
.Y(n_7834)
);

AOI221xp5_ASAP7_75t_L g7835 ( 
.A1(n_7802),
.A2(n_906),
.B1(n_903),
.B2(n_905),
.C(n_907),
.Y(n_7835)
);

AOI22xp5_ASAP7_75t_L g7836 ( 
.A1(n_7808),
.A2(n_908),
.B1(n_906),
.B2(n_907),
.Y(n_7836)
);

OR2x2_ASAP7_75t_L g7837 ( 
.A(n_7791),
.B(n_906),
.Y(n_7837)
);

AOI22xp5_ASAP7_75t_L g7838 ( 
.A1(n_7801),
.A2(n_910),
.B1(n_907),
.B2(n_909),
.Y(n_7838)
);

NOR2xp33_ASAP7_75t_L g7839 ( 
.A(n_7798),
.B(n_909),
.Y(n_7839)
);

OAI21xp33_ASAP7_75t_SL g7840 ( 
.A1(n_7811),
.A2(n_909),
.B(n_911),
.Y(n_7840)
);

NAND2xp5_ASAP7_75t_SL g7841 ( 
.A(n_7814),
.B(n_911),
.Y(n_7841)
);

NOR2xp33_ASAP7_75t_L g7842 ( 
.A(n_7792),
.B(n_7820),
.Y(n_7842)
);

INVx1_ASAP7_75t_L g7843 ( 
.A(n_7800),
.Y(n_7843)
);

NOR2x1_ASAP7_75t_L g7844 ( 
.A(n_7799),
.B(n_912),
.Y(n_7844)
);

NOR3x1_ASAP7_75t_L g7845 ( 
.A(n_7793),
.B(n_912),
.C(n_913),
.Y(n_7845)
);

AOI21xp5_ASAP7_75t_L g7846 ( 
.A1(n_7821),
.A2(n_912),
.B(n_913),
.Y(n_7846)
);

AOI22xp33_ASAP7_75t_L g7847 ( 
.A1(n_7807),
.A2(n_915),
.B1(n_913),
.B2(n_914),
.Y(n_7847)
);

INVxp67_ASAP7_75t_SL g7848 ( 
.A(n_7810),
.Y(n_7848)
);

AOI21xp33_ASAP7_75t_L g7849 ( 
.A1(n_7804),
.A2(n_914),
.B(n_915),
.Y(n_7849)
);

NOR4xp25_ASAP7_75t_L g7850 ( 
.A(n_7822),
.B(n_7805),
.C(n_7818),
.D(n_7815),
.Y(n_7850)
);

AND2x4_ASAP7_75t_L g7851 ( 
.A(n_7826),
.B(n_915),
.Y(n_7851)
);

OR2x2_ASAP7_75t_L g7852 ( 
.A(n_7825),
.B(n_916),
.Y(n_7852)
);

NOR2x1_ASAP7_75t_L g7853 ( 
.A(n_7830),
.B(n_916),
.Y(n_7853)
);

AOI21xp5_ASAP7_75t_L g7854 ( 
.A1(n_7839),
.A2(n_916),
.B(n_917),
.Y(n_7854)
);

AOI221x1_ASAP7_75t_L g7855 ( 
.A1(n_7843),
.A2(n_919),
.B1(n_917),
.B2(n_918),
.C(n_920),
.Y(n_7855)
);

NOR3xp33_ASAP7_75t_L g7856 ( 
.A(n_7823),
.B(n_917),
.C(n_918),
.Y(n_7856)
);

NOR2x1_ASAP7_75t_L g7857 ( 
.A(n_7829),
.B(n_919),
.Y(n_7857)
);

NAND2xp5_ASAP7_75t_L g7858 ( 
.A(n_7827),
.B(n_920),
.Y(n_7858)
);

AND2x4_ASAP7_75t_L g7859 ( 
.A(n_7827),
.B(n_920),
.Y(n_7859)
);

NOR3xp33_ASAP7_75t_L g7860 ( 
.A(n_7848),
.B(n_921),
.C(n_922),
.Y(n_7860)
);

NAND2xp5_ASAP7_75t_L g7861 ( 
.A(n_7832),
.B(n_1053),
.Y(n_7861)
);

OAI211xp5_ASAP7_75t_SL g7862 ( 
.A1(n_7834),
.A2(n_923),
.B(n_921),
.C(n_922),
.Y(n_7862)
);

NOR3xp33_ASAP7_75t_L g7863 ( 
.A(n_7837),
.B(n_7842),
.C(n_7841),
.Y(n_7863)
);

NOR5xp2_ASAP7_75t_L g7864 ( 
.A(n_7849),
.B(n_921),
.C(n_923),
.D(n_924),
.E(n_925),
.Y(n_7864)
);

NOR2x1_ASAP7_75t_L g7865 ( 
.A(n_7824),
.B(n_923),
.Y(n_7865)
);

AOI22xp5_ASAP7_75t_L g7866 ( 
.A1(n_7863),
.A2(n_7844),
.B1(n_7840),
.B2(n_7828),
.Y(n_7866)
);

NOR2x1_ASAP7_75t_L g7867 ( 
.A(n_7853),
.B(n_7833),
.Y(n_7867)
);

INVx2_ASAP7_75t_L g7868 ( 
.A(n_7859),
.Y(n_7868)
);

INVx1_ASAP7_75t_L g7869 ( 
.A(n_7861),
.Y(n_7869)
);

INVx1_ASAP7_75t_L g7870 ( 
.A(n_7858),
.Y(n_7870)
);

INVx1_ASAP7_75t_L g7871 ( 
.A(n_7865),
.Y(n_7871)
);

NAND5xp2_ASAP7_75t_L g7872 ( 
.A(n_7866),
.B(n_7850),
.C(n_7857),
.D(n_7845),
.E(n_7854),
.Y(n_7872)
);

OR4x2_ASAP7_75t_L g7873 ( 
.A(n_7868),
.B(n_7862),
.C(n_7860),
.D(n_7864),
.Y(n_7873)
);

INVx1_ASAP7_75t_L g7874 ( 
.A(n_7871),
.Y(n_7874)
);

CKINVDCx5p33_ASAP7_75t_R g7875 ( 
.A(n_7874),
.Y(n_7875)
);

INVx3_ASAP7_75t_SL g7876 ( 
.A(n_7872),
.Y(n_7876)
);

NAND4xp25_ASAP7_75t_L g7877 ( 
.A(n_7876),
.B(n_7869),
.C(n_7870),
.D(n_7867),
.Y(n_7877)
);

AOI221xp5_ASAP7_75t_L g7878 ( 
.A1(n_7877),
.A2(n_7875),
.B1(n_7873),
.B2(n_7852),
.C(n_7851),
.Y(n_7878)
);

INVx2_ASAP7_75t_SL g7879 ( 
.A(n_7878),
.Y(n_7879)
);

INVx3_ASAP7_75t_L g7880 ( 
.A(n_7878),
.Y(n_7880)
);

AND2x4_ASAP7_75t_L g7881 ( 
.A(n_7880),
.B(n_7846),
.Y(n_7881)
);

NOR2x1_ASAP7_75t_L g7882 ( 
.A(n_7879),
.B(n_7847),
.Y(n_7882)
);

AOI22x1_ASAP7_75t_L g7883 ( 
.A1(n_7881),
.A2(n_7856),
.B1(n_7836),
.B2(n_7835),
.Y(n_7883)
);

HB1xp67_ASAP7_75t_L g7884 ( 
.A(n_7883),
.Y(n_7884)
);

AOI222xp33_ASAP7_75t_L g7885 ( 
.A1(n_7884),
.A2(n_7882),
.B1(n_7838),
.B2(n_7855),
.C1(n_7831),
.C2(n_928),
.Y(n_7885)
);

AOI321xp33_ASAP7_75t_L g7886 ( 
.A1(n_7885),
.A2(n_924),
.A3(n_925),
.B1(n_926),
.B2(n_927),
.C(n_928),
.Y(n_7886)
);

NAND3xp33_ASAP7_75t_L g7887 ( 
.A(n_7886),
.B(n_924),
.C(n_925),
.Y(n_7887)
);

AOI22xp33_ASAP7_75t_R g7888 ( 
.A1(n_7887),
.A2(n_1048),
.B1(n_928),
.B2(n_926),
.Y(n_7888)
);

AO221x1_ASAP7_75t_L g7889 ( 
.A1(n_7888),
.A2(n_926),
.B1(n_927),
.B2(n_929),
.C(n_930),
.Y(n_7889)
);

OAI221xp5_ASAP7_75t_R g7890 ( 
.A1(n_7889),
.A2(n_1048),
.B1(n_929),
.B2(n_930),
.C(n_931),
.Y(n_7890)
);

AOI22xp33_ASAP7_75t_L g7891 ( 
.A1(n_7890),
.A2(n_931),
.B1(n_927),
.B2(n_930),
.Y(n_7891)
);

AOI211xp5_ASAP7_75t_L g7892 ( 
.A1(n_7891),
.A2(n_933),
.B(n_931),
.C(n_932),
.Y(n_7892)
);


endmodule