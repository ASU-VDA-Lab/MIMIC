module fake_jpeg_5675_n_89 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_89);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_89;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_14),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_55),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_51),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_47),
.B1(n_37),
.B2(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_64),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_56),
.B(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_48),
.B1(n_35),
.B2(n_50),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_72),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_49),
.B1(n_41),
.B2(n_39),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_75),
.B1(n_74),
.B2(n_46),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_60),
.Y(n_72)
);

A2O1A1O1Ixp25_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_20),
.B(n_2),
.C(n_4),
.D(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_45),
.C(n_65),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_76),
.A2(n_77),
.B(n_1),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_78),
.B(n_79),
.C(n_9),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_6),
.C(n_8),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_11),
.B(n_12),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_15),
.C(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_18),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_19),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_21),
.C(n_22),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_24),
.Y(n_89)
);


endmodule