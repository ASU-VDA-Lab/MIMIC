module fake_jpeg_32005_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_28),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_55),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_79),
.Y(n_91)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_54),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_66),
.B(n_72),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_60),
.A3(n_49),
.B1(n_64),
.B2(n_68),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_72),
.B(n_55),
.C(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_54),
.B1(n_53),
.B2(n_51),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_67),
.B1(n_61),
.B2(n_59),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_111),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_114),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_57),
.C(n_50),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_48),
.B1(n_24),
.B2(n_31),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

BUFx2_ASAP7_75t_SL g120 ( 
.A(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_1),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_23),
.B1(n_44),
.B2(n_43),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_129),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_4),
.B(n_5),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_133),
.B(n_13),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_7),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_34),
.B(n_41),
.C(n_9),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_36),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_7),
.B(n_8),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_12),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_20),
.C(n_33),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_47),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_136),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_137),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_136),
.B(n_129),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_150),
.C(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_141),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_138),
.B(n_132),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_151),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_158),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_165),
.A2(n_156),
.B(n_160),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_154),
.B(n_134),
.Y(n_167)
);


endmodule