module fake_jpeg_17029_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_29),
.A2(n_21),
.B1(n_15),
.B2(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_21),
.B1(n_17),
.B2(n_18),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_37),
.B1(n_43),
.B2(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_21),
.B1(n_18),
.B2(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_26),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_15),
.B1(n_30),
.B2(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_51),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_29),
.A3(n_31),
.B1(n_27),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_55),
.B1(n_33),
.B2(n_43),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_52),
.B1(n_36),
.B2(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_23),
.B1(n_25),
.B2(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_23),
.B1(n_22),
.B2(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx9p33_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_62),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_54),
.B1(n_45),
.B2(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_53),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_69),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_50),
.B1(n_48),
.B2(n_54),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_6),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_51),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_16),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_46),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_41),
.C(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_78),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_80),
.B1(n_86),
.B2(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_82),
.B1(n_85),
.B2(n_65),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_54),
.B1(n_45),
.B2(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_49),
.B1(n_42),
.B2(n_32),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_41),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_65),
.B1(n_68),
.B2(n_62),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_91),
.B1(n_94),
.B2(n_81),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_85),
.B(n_80),
.C(n_82),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_99),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_76),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_113),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_79),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_114),
.C(n_41),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_112),
.B1(n_105),
.B2(n_103),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_9),
.B1(n_7),
.B2(n_11),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_66),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_70),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_110),
.A2(n_96),
.B1(n_98),
.B2(n_94),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_109),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_90),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_120),
.C(n_121),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_34),
.C(n_38),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_34),
.C(n_38),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_19),
.C(n_14),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_126),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_128),
.B1(n_109),
.B2(n_16),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_41),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_139),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_133),
.B(n_143),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_106),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_19),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_112),
.B(n_109),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_13),
.B(n_32),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_22),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_122),
.C(n_121),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_13),
.B1(n_128),
.B2(n_11),
.Y(n_148)
);

OAI322xp33_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_13),
.A3(n_16),
.B1(n_41),
.B2(n_20),
.C1(n_19),
.C2(n_14),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_133),
.B(n_141),
.C(n_140),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_152),
.B(n_20),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_139),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_149),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_136),
.B1(n_134),
.B2(n_119),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_153),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_20),
.CI(n_14),
.CON(n_151),
.SN(n_151)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_20),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_19),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_145),
.A2(n_11),
.B(n_10),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_156),
.B(n_159),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_144),
.A2(n_150),
.B(n_146),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_162),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_10),
.B(n_9),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_8),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_158),
.A2(n_148),
.B1(n_153),
.B2(n_151),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_164),
.A2(n_5),
.B(n_1),
.Y(n_175)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_161),
.B(n_159),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_0),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_147),
.B1(n_8),
.B2(n_5),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_12),
.C(n_34),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_8),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_171),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_38),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_5),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_176),
.A3(n_165),
.B1(n_32),
.B2(n_3),
.C1(n_4),
.C2(n_1),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_177),
.C(n_12),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_180),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_25),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_168),
.A3(n_38),
.B1(n_25),
.B2(n_12),
.C1(n_4),
.C2(n_3),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_12),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.C(n_178),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_SL g185 ( 
.A1(n_184),
.A2(n_2),
.B(n_4),
.C(n_25),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_2),
.Y(n_186)
);


endmodule