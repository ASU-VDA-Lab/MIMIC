module real_aes_2240_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_0), .B(n_140), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_1), .A2(n_148), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_2), .B(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_3), .B(n_140), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_4), .B(n_167), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_5), .B(n_167), .Y(n_465) );
INVx1_ASAP7_75t_L g136 ( .A(n_6), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_7), .B(n_167), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g749 ( .A(n_8), .Y(n_749) );
NAND2xp33_ASAP7_75t_L g535 ( .A(n_9), .B(n_165), .Y(n_535) );
AND2x2_ASAP7_75t_L g170 ( .A(n_10), .B(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g181 ( .A(n_11), .B(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g127 ( .A(n_12), .Y(n_127) );
AOI221x1_ASAP7_75t_L g440 ( .A1(n_13), .A2(n_24), .B1(n_140), .B2(n_148), .C(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_14), .B(n_167), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_15), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_16), .B(n_140), .Y(n_531) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_17), .A2(n_182), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_18), .B(n_125), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_19), .B(n_167), .Y(n_518) );
AO21x1_ASAP7_75t_L g460 ( .A1(n_20), .A2(n_140), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_21), .B(n_140), .Y(n_221) );
INVx1_ASAP7_75t_L g112 ( .A(n_22), .Y(n_112) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_23), .A2(n_88), .B1(n_131), .B2(n_140), .Y(n_130) );
NAND2x1_ASAP7_75t_L g452 ( .A(n_25), .B(n_167), .Y(n_452) );
NAND2x1_ASAP7_75t_L g493 ( .A(n_26), .B(n_165), .Y(n_493) );
OR2x2_ASAP7_75t_L g128 ( .A(n_27), .B(n_85), .Y(n_128) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_27), .A2(n_85), .B(n_127), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_28), .B(n_165), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_29), .B(n_167), .Y(n_534) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_30), .A2(n_171), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_31), .B(n_165), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_32), .A2(n_148), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_33), .B(n_167), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_34), .A2(n_148), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g138 ( .A(n_35), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g146 ( .A(n_35), .B(n_136), .Y(n_146) );
INVx1_ASAP7_75t_L g152 ( .A(n_35), .Y(n_152) );
OR2x6_ASAP7_75t_L g110 ( .A(n_36), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_37), .B(n_140), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_38), .B(n_140), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_39), .B(n_167), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_40), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_41), .B(n_165), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_42), .B(n_140), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_43), .A2(n_148), .B(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_44), .A2(n_148), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_45), .B(n_165), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_46), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_47), .B(n_165), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_48), .B(n_140), .Y(n_233) );
INVx1_ASAP7_75t_L g134 ( .A(n_49), .Y(n_134) );
INVx1_ASAP7_75t_L g143 ( .A(n_49), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_50), .B(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g201 ( .A(n_51), .B(n_125), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_52), .B(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_53), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_54), .B(n_167), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_55), .B(n_165), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_56), .A2(n_148), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_57), .B(n_140), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_58), .A2(n_114), .B1(n_721), .B2(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_58), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_59), .B(n_140), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_60), .A2(n_148), .B(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g227 ( .A(n_61), .B(n_126), .Y(n_227) );
AO21x1_ASAP7_75t_L g462 ( .A1(n_62), .A2(n_148), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_63), .B(n_140), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_64), .B(n_165), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_65), .B(n_140), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_66), .B(n_165), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_67), .A2(n_92), .B1(n_148), .B2(n_150), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_68), .B(n_167), .Y(n_224) );
AND2x2_ASAP7_75t_L g476 ( .A(n_69), .B(n_126), .Y(n_476) );
INVx1_ASAP7_75t_L g139 ( .A(n_70), .Y(n_139) );
INVx1_ASAP7_75t_L g145 ( .A(n_70), .Y(n_145) );
AND2x2_ASAP7_75t_L g496 ( .A(n_71), .B(n_171), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_72), .B(n_165), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_73), .A2(n_148), .B(n_205), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_74), .A2(n_148), .B(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_75), .A2(n_148), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g218 ( .A(n_76), .B(n_126), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_77), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g113 ( .A(n_78), .Y(n_113) );
AND2x2_ASAP7_75t_L g481 ( .A(n_79), .B(n_171), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_80), .B(n_140), .Y(n_520) );
AND2x2_ASAP7_75t_L g194 ( .A(n_81), .B(n_182), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_82), .A2(n_102), .B1(n_719), .B2(n_724), .Y(n_718) );
AND2x2_ASAP7_75t_L g461 ( .A(n_83), .B(n_208), .Y(n_461) );
INVx1_ASAP7_75t_L g102 ( .A(n_84), .Y(n_102) );
AND2x2_ASAP7_75t_L g455 ( .A(n_86), .B(n_171), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_87), .B(n_165), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_89), .B(n_167), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_90), .B(n_165), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_91), .A2(n_148), .B(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_93), .A2(n_148), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_94), .B(n_167), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_95), .B(n_167), .Y(n_486) );
BUFx2_ASAP7_75t_L g226 ( .A(n_96), .Y(n_226) );
BUFx2_ASAP7_75t_L g730 ( .A(n_97), .Y(n_730) );
BUFx2_ASAP7_75t_SL g739 ( .A(n_97), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_98), .A2(n_148), .B(n_533), .Y(n_532) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_743), .B(n_750), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_726), .B(n_737), .Y(n_100) );
OAI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_103), .B(n_718), .Y(n_101) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_114), .B1(n_433), .B2(n_713), .Y(n_104) );
CKINVDCx6p67_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx11_ASAP7_75t_R g720 ( .A(n_106), .Y(n_720) );
INVx3_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x6_ASAP7_75t_SL g108 ( .A(n_109), .B(n_110), .Y(n_108) );
OR2x6_ASAP7_75t_SL g716 ( .A(n_109), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g725 ( .A(n_109), .B(n_110), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_109), .B(n_717), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g717 ( .A(n_110), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx4_ASAP7_75t_L g721 ( .A(n_114), .Y(n_721) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_370), .Y(n_114) );
NAND3xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_286), .C(n_323), .Y(n_115) );
NOR3xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_254), .C(n_269), .Y(n_116) );
OAI221xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_198), .B1(n_228), .B2(n_240), .C(n_241), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_120), .B(n_183), .Y(n_119) );
OAI22xp33_ASAP7_75t_SL g314 ( .A1(n_120), .A2(n_278), .B1(n_315), .B2(n_318), .Y(n_314) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_155), .Y(n_120) );
OAI21xp33_ASAP7_75t_SL g324 ( .A1(n_121), .A2(n_325), .B(n_331), .Y(n_324) );
OR2x2_ASAP7_75t_L g353 ( .A(n_121), .B(n_185), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_121), .B(n_273), .Y(n_354) );
INVx2_ASAP7_75t_L g385 ( .A(n_121), .Y(n_385) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_122), .B(n_245), .Y(n_366) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g240 ( .A(n_123), .B(n_158), .Y(n_240) );
BUFx3_ASAP7_75t_L g266 ( .A(n_123), .Y(n_266) );
AND2x2_ASAP7_75t_L g402 ( .A(n_123), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g425 ( .A(n_123), .B(n_186), .Y(n_425) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
AND2x4_ASAP7_75t_L g197 ( .A(n_124), .B(n_129), .Y(n_197) );
AO21x2_ASAP7_75t_L g129 ( .A1(n_125), .A2(n_130), .B(n_147), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_125), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_125), .A2(n_189), .B(n_190), .Y(n_188) );
OA21x2_ASAP7_75t_L g439 ( .A1(n_125), .A2(n_440), .B(n_444), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_125), .A2(n_483), .B(n_484), .Y(n_482) );
OA21x2_ASAP7_75t_L g583 ( .A1(n_125), .A2(n_440), .B(n_444), .Y(n_583) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x4_ASAP7_75t_L g208 ( .A(n_127), .B(n_128), .Y(n_208) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g149 ( .A(n_134), .B(n_136), .Y(n_149) );
AND2x4_ASAP7_75t_L g167 ( .A(n_134), .B(n_144), .Y(n_167) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x6_ASAP7_75t_L g148 ( .A(n_138), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
AND2x6_ASAP7_75t_L g165 ( .A(n_139), .B(n_142), .Y(n_165) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
AND2x4_ASAP7_75t_L g150 ( .A(n_149), .B(n_151), .Y(n_150) );
NOR2x1p5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_156), .B(n_186), .Y(n_345) );
INVx1_ASAP7_75t_L g382 ( .A(n_156), .Y(n_382) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_172), .Y(n_156) );
AND2x2_ASAP7_75t_L g196 ( .A(n_157), .B(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g403 ( .A(n_157), .Y(n_403) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g246 ( .A(n_158), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_158), .B(n_172), .Y(n_247) );
AND2x2_ASAP7_75t_L g268 ( .A(n_158), .B(n_187), .Y(n_268) );
AND2x2_ASAP7_75t_L g350 ( .A(n_158), .B(n_173), .Y(n_350) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_170), .Y(n_158) );
INVx4_ASAP7_75t_L g171 ( .A(n_159), .Y(n_171) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx4f_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_169), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_166), .B(n_168), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_165), .B(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_168), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_168), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_168), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_168), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_168), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_168), .A2(n_236), .B(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_168), .A2(n_442), .B(n_443), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_168), .A2(n_452), .B(n_453), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_168), .A2(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_168), .A2(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_168), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_168), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_168), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_168), .A2(n_534), .B(n_535), .Y(n_533) );
INVx3_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
AND2x4_ASAP7_75t_SL g243 ( .A(n_172), .B(n_187), .Y(n_243) );
INVx1_ASAP7_75t_L g274 ( .A(n_172), .Y(n_274) );
INVx2_ASAP7_75t_L g282 ( .A(n_172), .Y(n_282) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_172), .Y(n_306) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_173), .Y(n_195) );
AOI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_181), .Y(n_173) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_174), .A2(n_490), .B(n_496), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_180), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_182), .A2(n_221), .B(n_222), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_196), .Y(n_183) );
AND2x2_ASAP7_75t_L g421 ( .A(n_184), .B(n_284), .Y(n_421) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_195), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g280 ( .A(n_186), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g332 ( .A(n_186), .B(n_247), .Y(n_332) );
AND2x2_ASAP7_75t_L g349 ( .A(n_186), .B(n_350), .Y(n_349) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x4_ASAP7_75t_L g273 ( .A(n_187), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g289 ( .A(n_187), .Y(n_289) );
AND2x2_ASAP7_75t_L g333 ( .A(n_187), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g340 ( .A(n_187), .B(n_341), .Y(n_340) );
NOR2x1_ASAP7_75t_L g355 ( .A(n_187), .B(n_246), .Y(n_355) );
BUFx2_ASAP7_75t_L g365 ( .A(n_187), .Y(n_365) );
AND2x2_ASAP7_75t_L g390 ( .A(n_187), .B(n_350), .Y(n_390) );
AND2x2_ASAP7_75t_L g411 ( .A(n_187), .B(n_412), .Y(n_411) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_194), .Y(n_187) );
INVx1_ASAP7_75t_L g342 ( .A(n_195), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_196), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g372 ( .A(n_196), .B(n_243), .Y(n_372) );
INVx3_ASAP7_75t_L g279 ( .A(n_197), .Y(n_279) );
AND2x2_ASAP7_75t_L g412 ( .A(n_197), .B(n_334), .Y(n_412) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_199), .A2(n_242), .B1(n_247), .B2(n_248), .Y(n_241) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
INVx4_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
INVx2_ASAP7_75t_L g276 ( .A(n_200), .Y(n_276) );
NAND2x1_ASAP7_75t_L g302 ( .A(n_200), .B(n_219), .Y(n_302) );
OR2x2_ASAP7_75t_L g317 ( .A(n_200), .B(n_252), .Y(n_317) );
OR2x2_ASAP7_75t_SL g344 ( .A(n_200), .B(n_316), .Y(n_344) );
AND2x2_ASAP7_75t_L g357 ( .A(n_200), .B(n_231), .Y(n_357) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_200), .Y(n_378) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_208), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_208), .A2(n_233), .B(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_208), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_SL g514 ( .A(n_208), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_208), .A2(n_531), .B(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g257 ( .A(n_209), .Y(n_257) );
AND2x2_ASAP7_75t_L g389 ( .A(n_209), .B(n_363), .Y(n_389) );
NOR2x1_ASAP7_75t_SL g209 ( .A(n_210), .B(n_219), .Y(n_209) );
AND2x2_ASAP7_75t_L g230 ( .A(n_210), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g406 ( .A(n_210), .B(n_329), .Y(n_406) );
AO21x1_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_210) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_253) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_211), .A2(n_449), .B(n_455), .Y(n_448) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_211), .A2(n_470), .B(n_476), .Y(n_469) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_211), .A2(n_470), .B(n_476), .Y(n_503) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_211), .A2(n_449), .B(n_455), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_217), .Y(n_212) );
OR2x2_ASAP7_75t_L g238 ( .A(n_219), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g249 ( .A(n_219), .B(n_239), .Y(n_249) );
AND2x2_ASAP7_75t_L g295 ( .A(n_219), .B(n_252), .Y(n_295) );
OR2x2_ASAP7_75t_L g316 ( .A(n_219), .B(n_231), .Y(n_316) );
INVx2_ASAP7_75t_SL g322 ( .A(n_219), .Y(n_322) );
AND2x2_ASAP7_75t_L g328 ( .A(n_219), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g338 ( .A(n_219), .B(n_321), .Y(n_338) );
BUFx2_ASAP7_75t_L g360 ( .A(n_219), .Y(n_360) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_227), .Y(n_219) );
INVx2_ASAP7_75t_L g407 ( .A(n_228), .Y(n_407) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_238), .Y(n_228) );
OR2x2_ASAP7_75t_L g432 ( .A(n_229), .B(n_276), .Y(n_432) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_230), .B(n_239), .Y(n_298) );
AND2x2_ASAP7_75t_L g369 ( .A(n_230), .B(n_249), .Y(n_369) );
INVx1_ASAP7_75t_L g251 ( .A(n_231), .Y(n_251) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_231), .Y(n_260) );
INVx1_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
INVx2_ASAP7_75t_L g329 ( .A(n_231), .Y(n_329) );
NOR2xp67_ASAP7_75t_L g259 ( .A(n_239), .B(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_L g319 ( .A(n_239), .Y(n_319) );
INVx2_ASAP7_75t_SL g395 ( .A(n_240), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_242), .A2(n_297), .B1(n_299), .B2(n_303), .Y(n_296) );
AND2x2_ASAP7_75t_SL g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g423 ( .A(n_243), .B(n_279), .Y(n_423) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_245), .B(n_289), .Y(n_368) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g334 ( .A(n_246), .B(n_282), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_247), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g277 ( .A(n_248), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_248), .A2(n_392), .B1(n_396), .B2(n_398), .C(n_400), .Y(n_391) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
AND2x2_ASAP7_75t_L g261 ( .A(n_249), .B(n_262), .Y(n_261) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_249), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_249), .B(n_292), .Y(n_347) );
INVx1_ASAP7_75t_SL g343 ( .A(n_250), .Y(n_343) );
AOI221xp5_ASAP7_75t_SL g371 ( .A1(n_250), .A2(n_261), .B1(n_372), .B2(n_373), .C(n_376), .Y(n_371) );
AOI322xp5_ASAP7_75t_L g404 ( .A1(n_250), .A2(n_322), .A3(n_349), .B1(n_405), .B2(n_407), .C1(n_408), .C2(n_411), .Y(n_404) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
BUFx2_ASAP7_75t_L g271 ( .A(n_251), .Y(n_271) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_252), .Y(n_263) );
INVx2_ASAP7_75t_L g321 ( .A(n_252), .Y(n_321) );
AND2x2_ASAP7_75t_L g362 ( .A(n_252), .B(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OA21x2_ASAP7_75t_SL g254 ( .A1(n_255), .A2(n_261), .B(n_264), .Y(n_254) );
AOI211xp5_ASAP7_75t_L g424 ( .A1(n_255), .A2(n_425), .B(n_426), .C(n_430), .Y(n_424) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OR2x2_ASAP7_75t_L g313 ( .A(n_257), .B(n_275), .Y(n_313) );
OR2x2_ASAP7_75t_L g397 ( .A(n_257), .B(n_292), .Y(n_397) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g337 ( .A(n_259), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g415 ( .A(n_262), .Y(n_415) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
OR2x2_ASAP7_75t_L g270 ( .A(n_266), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g305 ( .A(n_268), .B(n_306), .Y(n_305) );
OAI322xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_272), .A3(n_275), .B1(n_277), .B2(n_278), .C1(n_283), .C2(n_285), .Y(n_269) );
INVx1_ASAP7_75t_L g311 ( .A(n_270), .Y(n_311) );
OR2x2_ASAP7_75t_L g283 ( .A(n_272), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_272), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g294 ( .A(n_276), .B(n_295), .Y(n_294) );
OAI32xp33_ASAP7_75t_L g339 ( .A1(n_276), .A2(n_340), .A3(n_343), .B1(n_344), .B2(n_345), .Y(n_339) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g284 ( .A(n_279), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_279), .B(n_342), .Y(n_341) );
NOR2x1_ASAP7_75t_L g381 ( .A(n_279), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g405 ( .A(n_279), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g326 ( .A(n_280), .Y(n_326) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_284), .B(n_350), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_307), .Y(n_286) );
OAI21xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B(n_296), .Y(n_287) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_SL g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g356 ( .A(n_295), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_298), .A2(n_318), .B1(n_420), .B2(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_347), .B(n_348), .C(n_351), .Y(n_346) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx3_ASAP7_75t_L g428 ( .A(n_302), .Y(n_428) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g309 ( .A(n_306), .Y(n_309) );
AO21x1_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_310), .B(n_314), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g374 ( .A(n_309), .Y(n_374) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_315), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g330 ( .A(n_317), .Y(n_330) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g387 ( .A(n_320), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NOR3xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_346), .C(n_358), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OAI21xp5_ASAP7_75t_SL g388 ( .A1(n_327), .A2(n_389), .B(n_390), .Y(n_388) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g363 ( .A(n_329), .Y(n_363) );
O2A1O1Ixp5_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_333), .B(n_335), .C(n_339), .Y(n_331) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_341), .Y(n_431) );
INVx2_ASAP7_75t_L g416 ( .A(n_344), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_345), .A2(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g410 ( .A(n_350), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .A3(n_355), .B(n_356), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g429 ( .A(n_357), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_364), .B(n_367), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
BUFx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g379 ( .A(n_362), .Y(n_379) );
AOI21xp33_ASAP7_75t_SL g426 ( .A1(n_364), .A2(n_427), .B(n_429), .Y(n_426) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g394 ( .A(n_365), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_365), .B(n_385), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_365), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g375 ( .A(n_366), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
NAND5xp2_ASAP7_75t_L g370 ( .A(n_371), .B(n_391), .C(n_404), .D(n_413), .E(n_424), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B1(n_383), .B2(n_386), .C(n_388), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B(n_419), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g723 ( .A(n_433), .Y(n_723) );
NAND4xp75_ASAP7_75t_L g433 ( .A(n_434), .B(n_623), .C(n_663), .D(n_692), .Y(n_433) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_585), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_542), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_477), .B(n_497), .Y(n_436) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_438), .B(n_445), .Y(n_437) );
AND2x4_ASAP7_75t_L g541 ( .A(n_438), .B(n_502), .Y(n_541) );
INVx1_ASAP7_75t_SL g594 ( .A(n_438), .Y(n_594) );
AOI21xp33_ASAP7_75t_L g629 ( .A1(n_438), .A2(n_630), .B(n_633), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_SL g633 ( .A1(n_438), .A2(n_634), .B(n_635), .C(n_636), .Y(n_633) );
NAND2x1_ASAP7_75t_L g674 ( .A(n_438), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_438), .B(n_635), .Y(n_696) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g500 ( .A(n_439), .Y(n_500) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_439), .Y(n_573) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_456), .Y(n_445) );
AND2x2_ASAP7_75t_L g565 ( .A(n_446), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g646 ( .A(n_446), .B(n_502), .Y(n_646) );
INVx1_ASAP7_75t_L g706 ( .A(n_446), .Y(n_706) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g550 ( .A(n_447), .B(n_468), .Y(n_550) );
AND2x2_ASAP7_75t_L g675 ( .A(n_447), .B(n_469), .Y(n_675) );
AND2x2_ASAP7_75t_L g680 ( .A(n_447), .B(n_640), .Y(n_680) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g556 ( .A(n_448), .Y(n_556) );
BUFx3_ASAP7_75t_L g589 ( .A(n_448), .Y(n_589) );
AND2x2_ASAP7_75t_L g635 ( .A(n_448), .B(n_469), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_454), .Y(n_449) );
AND2x2_ASAP7_75t_L g620 ( .A(n_456), .B(n_499), .Y(n_620) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_468), .Y(n_456) );
AND2x4_ASAP7_75t_L g502 ( .A(n_457), .B(n_503), .Y(n_502) );
OR2x2_ASAP7_75t_L g612 ( .A(n_457), .B(n_596), .Y(n_612) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_457), .B(n_583), .Y(n_655) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g591 ( .A(n_458), .Y(n_591) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g552 ( .A(n_459), .Y(n_552) );
OAI21x1_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_462), .B(n_466), .Y(n_459) );
INVx1_ASAP7_75t_L g467 ( .A(n_461), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_468), .B(n_552), .Y(n_555) );
AND2x2_ASAP7_75t_L g640 ( .A(n_468), .B(n_583), .Y(n_640) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g637 ( .A(n_469), .B(n_500), .Y(n_637) );
AND2x2_ASAP7_75t_L g657 ( .A(n_469), .B(n_583), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_471), .B(n_475), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_477), .B(n_546), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_477), .A2(n_669), .B1(n_670), .B2(n_671), .C(n_673), .Y(n_668) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI332xp33_ASAP7_75t_L g702 ( .A1(n_478), .A2(n_562), .A3(n_569), .B1(n_628), .B2(n_703), .B3(n_704), .C1(n_705), .C2(n_707), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .Y(n_478) );
AND2x2_ASAP7_75t_L g508 ( .A(n_479), .B(n_489), .Y(n_508) );
AND2x2_ASAP7_75t_L g525 ( .A(n_479), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g537 ( .A(n_479), .Y(n_537) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_479), .B(n_538), .Y(n_597) );
INVx5_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR2x1_ASAP7_75t_SL g559 ( .A(n_480), .B(n_526), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_480), .B(n_488), .Y(n_563) );
AND2x2_ASAP7_75t_L g570 ( .A(n_480), .B(n_489), .Y(n_570) );
BUFx2_ASAP7_75t_L g605 ( .A(n_480), .Y(n_605) );
AND2x2_ASAP7_75t_L g660 ( .A(n_480), .B(n_529), .Y(n_660) );
OR2x6_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
OR2x2_ASAP7_75t_L g528 ( .A(n_488), .B(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g538 ( .A(n_488), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g578 ( .A(n_488), .Y(n_578) );
AND2x2_ASAP7_75t_L g648 ( .A(n_488), .B(n_547), .Y(n_648) );
AND2x2_ASAP7_75t_L g661 ( .A(n_488), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_488), .B(n_662), .Y(n_679) );
INVx4_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_489), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .Y(n_490) );
OAI32xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_504), .A3(n_509), .B1(n_523), .B2(n_540), .Y(n_497) );
INVx2_ASAP7_75t_L g606 ( .A(n_498), .Y(n_606) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g617 ( .A(n_499), .Y(n_617) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g551 ( .A(n_500), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g684 ( .A(n_500), .B(n_589), .Y(n_684) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g596 ( .A(n_503), .Y(n_596) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVx2_ASAP7_75t_L g584 ( .A(n_506), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_506), .B(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_SL g595 ( .A(n_507), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g672 ( .A(n_507), .Y(n_672) );
AND2x2_ASAP7_75t_L g690 ( .A(n_507), .B(n_552), .Y(n_690) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp67_ASAP7_75t_SL g634 ( .A(n_510), .B(n_563), .Y(n_634) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_511), .B(n_545), .Y(n_632) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g708 ( .A(n_512), .B(n_578), .Y(n_708) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g539 ( .A(n_513), .Y(n_539) );
INVx2_ASAP7_75t_L g580 ( .A(n_513), .Y(n_580) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_521), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_514), .B(n_522), .Y(n_521) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_514), .A2(n_515), .B(n_521), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_520), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_536), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_524), .B(n_582), .Y(n_667) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
AND3x2_ASAP7_75t_L g622 ( .A(n_525), .B(n_569), .C(n_578), .Y(n_622) );
AND2x2_ASAP7_75t_L g546 ( .A(n_526), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_526), .B(n_529), .Y(n_603) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g557 ( .A(n_528), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g547 ( .A(n_529), .Y(n_547) );
INVx1_ASAP7_75t_L g562 ( .A(n_529), .Y(n_562) );
BUFx3_ASAP7_75t_L g569 ( .A(n_529), .Y(n_569) );
AND2x2_ASAP7_75t_L g579 ( .A(n_529), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x4_ASAP7_75t_L g588 ( .A(n_537), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_537), .B(n_547), .Y(n_631) );
AND2x2_ASAP7_75t_L g587 ( .A(n_538), .B(n_562), .Y(n_587) );
INVx2_ASAP7_75t_L g614 ( .A(n_538), .Y(n_614) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AOI211xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_548), .B(n_553), .C(n_574), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_543), .A2(n_670), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_546), .B(n_605), .Y(n_604) );
AOI211xp5_ASAP7_75t_SL g624 ( .A1(n_546), .A2(n_625), .B(n_629), .C(n_638), .Y(n_624) );
AND2x2_ASAP7_75t_L g610 ( .A(n_547), .B(n_570), .Y(n_610) );
OR2x2_ASAP7_75t_L g613 ( .A(n_547), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_550), .B(n_655), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_551), .B(n_596), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_551), .A2(n_577), .B1(n_657), .B2(n_660), .C(n_666), .Y(n_665) );
AND2x4_ASAP7_75t_L g582 ( .A(n_552), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g628 ( .A(n_552), .B(n_583), .Y(n_628) );
OAI221xp5_ASAP7_75t_SL g553 ( .A1(n_554), .A2(n_557), .B1(n_560), .B2(n_564), .C(n_567), .Y(n_553) );
AND2x2_ASAP7_75t_L g699 ( .A(n_554), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
INVx1_ASAP7_75t_L g652 ( .A(n_556), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_557), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g571 ( .A(n_559), .B(n_562), .Y(n_571) );
AND2x2_ASAP7_75t_L g647 ( .A(n_559), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g572 ( .A(n_566), .B(n_573), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_571), .B(n_572), .Y(n_567) );
INVx1_ASAP7_75t_L g691 ( .A(n_568), .Y(n_691) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g670 ( .A(n_569), .B(n_597), .Y(n_670) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_570), .B(n_579), .Y(n_643) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_581), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_575), .A2(n_609), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g681 ( .A(n_575), .Y(n_681) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g601 ( .A(n_578), .Y(n_601) );
INVx1_ASAP7_75t_L g662 ( .A(n_580), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_582), .B(n_652), .Y(n_703) );
AND2x2_ASAP7_75t_L g671 ( .A(n_583), .B(n_672), .Y(n_671) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_584), .A2(n_665), .B(n_668), .C(n_676), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_607), .Y(n_585) );
AOI322xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .A3(n_590), .B1(n_592), .B2(n_597), .C1(n_598), .C2(n_606), .Y(n_586) );
CKINVDCx16_ASAP7_75t_R g704 ( .A(n_588), .Y(n_704) );
AND2x2_ASAP7_75t_L g654 ( .A(n_589), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g688 ( .A(n_589), .Y(n_688) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_SL g639 ( .A(n_591), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_SL g645 ( .A(n_591), .B(n_637), .Y(n_645) );
AND2x2_ASAP7_75t_L g669 ( .A(n_591), .B(n_635), .Y(n_669) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_L g641 ( .A(n_595), .Y(n_641) );
NAND2xp33_ASAP7_75t_SL g598 ( .A(n_599), .B(n_604), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_SL g644 ( .A1(n_600), .A2(n_645), .B1(n_646), .B2(n_647), .C(n_649), .Y(n_644) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g711 ( .A(n_603), .Y(n_711) );
AOI211xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B(n_611), .C(n_615), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g686 ( .A(n_610), .Y(n_686) );
INVx1_ASAP7_75t_L g618 ( .A(n_612), .Y(n_618) );
OR2x2_ASAP7_75t_L g705 ( .A(n_612), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_SL g701 ( .A(n_613), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_619), .B(n_621), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_617), .B(n_635), .Y(n_712) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_644), .Y(n_623) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_627), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
OR2x2_ASAP7_75t_L g678 ( .A(n_631), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_641), .B(n_642), .Y(n_638) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AOI31xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .A3(n_656), .B(n_658), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_655), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B1(n_681), .B2(n_682), .C(n_685), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_689), .B2(n_691), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g689 ( .A(n_690), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_702), .C(n_709), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx4f_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g722 ( .A(n_715), .Y(n_722) );
CKINVDCx11_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_724), .B(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_731), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_732), .A2(n_733), .B(n_741), .Y(n_740) );
NOR2xp33_ASAP7_75t_SL g732 ( .A(n_733), .B(n_736), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx3_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g752 ( .A(n_746), .Y(n_752) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
endmodule