module fake_ariane_2189_n_3863 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_541, n_499, n_789, n_788, n_12, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_790, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_738, n_758, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_158, n_69, n_259, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_256, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_780, n_175, n_711, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_804, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_83, n_389, n_800, n_657, n_513, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_785, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_793, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_792, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_799, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_3863);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_790;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_256;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_780;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_804;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_785;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_793;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_3863;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_3619;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_3181;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_2407;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_3765;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_3719;
wire n_2731;
wire n_3703;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_2278;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_829;
wire n_1062;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_3856;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2663;
wire n_2233;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3830;
wire n_821;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_3315;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_3606;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_1074;
wire n_3230;
wire n_859;
wire n_3793;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_2650;
wire n_863;
wire n_1254;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_3828;
wire n_3073;
wire n_2060;
wire n_1295;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_1013;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3728;
wire n_1840;
wire n_1230;
wire n_2739;
wire n_3739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_3271;
wire n_844;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_1267;
wire n_3164;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_1790;
wire n_1354;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_3458;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3850;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_3777;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_851;
wire n_1590;
wire n_3280;
wire n_1351;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_3862;
wire n_930;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_1179;
wire n_3284;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_1468;
wire n_1661;
wire n_1253;
wire n_2791;
wire n_2683;
wire n_3212;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_2970;
wire n_3159;
wire n_966;
wire n_992;
wire n_955;
wire n_3549;
wire n_3624;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_3538;
wire n_1376;
wire n_3839;
wire n_1972;
wire n_1178;
wire n_2015;
wire n_1292;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3666;
wire n_3629;
wire n_3372;
wire n_990;
wire n_1623;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_867;
wire n_2147;
wire n_3479;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3724;
wire n_1920;
wire n_2083;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_3046;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_3741;
wire n_2388;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_2567;
wire n_3496;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_976;
wire n_3567;
wire n_909;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_965;
wire n_1914;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1234;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_2632;
wire n_1255;
wire n_1646;
wire n_3031;
wire n_2262;
wire n_3179;
wire n_2565;
wire n_1237;
wire n_3262;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3615;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_2640;
wire n_1163;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_3642;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3513;
wire n_3498;
wire n_3682;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_3508;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_1304;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3599;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_3477;
wire n_3286;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3788;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_3569;
wire n_3542;
wire n_2523;
wire n_1945;
wire n_3835;
wire n_3837;
wire n_1015;
wire n_2496;
wire n_1377;
wire n_1614;
wire n_2418;
wire n_1162;
wire n_2031;
wire n_1258;
wire n_3260;
wire n_3349;
wire n_3761;
wire n_3819;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3653;
wire n_3035;
wire n_3823;
wire n_887;
wire n_3403;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_1202;
wire n_2254;
wire n_3290;
wire n_3130;
wire n_1498;
wire n_1188;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_3602;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3492;
wire n_3501;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3737;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2949;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_1711;
wire n_1219;
wire n_1919;
wire n_2994;
wire n_2508;
wire n_1791;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_3826;
wire n_2266;
wire n_3417;
wire n_2449;
wire n_890;
wire n_842;
wire n_3626;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_1373;
wire n_1975;
wire n_1081;
wire n_1388;
wire n_2119;
wire n_1540;
wire n_1719;
wire n_1266;
wire n_2742;
wire n_3671;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_915;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_3367;
wire n_3669;
wire n_837;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_3795;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1714;
wire n_1044;
wire n_2696;
wire n_3340;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_873;
wire n_2157;
wire n_1966;
wire n_2468;
wire n_2171;
wire n_1243;
wire n_1400;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_3836;
wire n_3302;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_3097;
wire n_3507;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_1318;
wire n_854;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_3789;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_1873;
wire n_1137;
wire n_1733;
wire n_1856;
wire n_1476;
wire n_1524;
wire n_2723;
wire n_2016;
wire n_2725;
wire n_2667;
wire n_2928;
wire n_943;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_3746;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_3787;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_3753;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2720;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_3843;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3640;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_2936;
wire n_1154;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_3718;
wire n_2022;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2911;
wire n_2890;
wire n_3381;
wire n_3455;
wire n_3736;
wire n_891;
wire n_3313;
wire n_885;
wire n_1659;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_3317;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_1151;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_3605;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_3809;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_3573;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_3654;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_2665;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_3842;
wire n_2044;
wire n_928;
wire n_1153;
wire n_3769;
wire n_825;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_914;
wire n_1116;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_3462;
wire n_1197;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3731;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_3444;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_3851;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_2234;
wire n_1341;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3322;
wire n_1440;
wire n_3175;
wire n_2666;
wire n_3289;
wire n_1370;
wire n_1603;
wire n_2935;
wire n_2401;
wire n_889;
wire n_3822;
wire n_3255;
wire n_3818;
wire n_1549;
wire n_1066;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_911;
wire n_2658;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1534;
wire n_1065;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_3376;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_3770;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_3790;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_3405;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_2007;
wire n_1056;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1803;
wire n_1444;
wire n_1749;
wire n_820;
wire n_1653;
wire n_872;
wire n_3409;
wire n_3522;
wire n_3583;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3241;
wire n_3802;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_3481;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_3442;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_2638;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_2828;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_3553;
wire n_2305;
wire n_3645;
wire n_880;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_1175;
wire n_2299;
wire n_3751;
wire n_3402;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_2951;
wire n_3807;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_932;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_3470;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3844;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3677;
wire n_1564;
wire n_2010;
wire n_3676;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3576;
wire n_3558;
wire n_3782;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3658;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_2639;
wire n_3521;
wire n_3855;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_1663;
wire n_919;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_3360;
wire n_1930;
wire n_3687;
wire n_1809;
wire n_2787;
wire n_3585;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_3575;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_3633;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3379;
wire n_3111;
wire n_2212;
wire n_3838;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_2569;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_3316;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_3351;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_3776;
wire n_2775;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_2351;
wire n_1619;
wire n_3303;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_3445;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3285;
wire n_3824;
wire n_3825;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_1150;
wire n_977;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_3845;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_3371;
wire n_1781;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_881;
wire n_1477;
wire n_1777;
wire n_1019;
wire n_2188;
wire n_2097;
wire n_1982;
wire n_3366;
wire n_3461;
wire n_2430;
wire n_2504;
wire n_910;
wire n_1410;
wire n_939;
wire n_2297;
wire n_3094;
wire n_3441;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_2513;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_2957;
wire n_1199;
wire n_865;
wire n_1983;
wire n_1273;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3820;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_3763;
wire n_1946;
wire n_2148;
wire n_933;
wire n_3244;
wire n_3499;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1821;
wire n_1168;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3762;
wire n_3794;
wire n_3593;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_3293;
wire n_3361;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_3707;
wire n_2052;
wire n_1091;
wire n_2485;
wire n_3779;
wire n_3149;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_1581;
wire n_3849;
wire n_1928;
wire n_946;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_2792;
wire n_1818;
wire n_1146;
wire n_3398;
wire n_3709;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3592;
wire n_3557;
wire n_3725;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_3505;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_3547;
wire n_3771;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_3041;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1981;
wire n_1069;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g817 ( 
.A(n_285),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_460),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_155),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_145),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_471),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_767),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_786),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_489),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_156),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_51),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_130),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_674),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_680),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_438),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_176),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_110),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_155),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_290),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_730),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_593),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_136),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_18),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_791),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_253),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_83),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_636),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_296),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_546),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_115),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_737),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_586),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_659),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_537),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_742),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_554),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_23),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_157),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_59),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_777),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_425),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_219),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_338),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_657),
.Y(n_859)
);

CKINVDCx14_ASAP7_75t_R g860 ( 
.A(n_336),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_183),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_215),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_489),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_256),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_65),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_196),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_286),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_240),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_161),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_769),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_799),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_515),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_233),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_688),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_116),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_136),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_280),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_425),
.Y(n_878)
);

CKINVDCx16_ASAP7_75t_R g879 ( 
.A(n_734),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_153),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_404),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_459),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_812),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_686),
.Y(n_884)
);

INVxp67_ASAP7_75t_L g885 ( 
.A(n_701),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_521),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_521),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_599),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_94),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_128),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_446),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_217),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_46),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_575),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_287),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_60),
.Y(n_896)
);

CKINVDCx16_ASAP7_75t_R g897 ( 
.A(n_661),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_450),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_172),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_330),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_32),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_653),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_494),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_577),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_471),
.Y(n_905)
);

INVx1_ASAP7_75t_SL g906 ( 
.A(n_101),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_545),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_219),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_524),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_583),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_623),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_523),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_269),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_739),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_670),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_760),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_539),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_152),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_169),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_753),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_604),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_781),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_330),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_630),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_794),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_774),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_573),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_774),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_407),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_77),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_169),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_543),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_810),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_434),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_589),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_395),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_93),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_280),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_295),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_314),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_409),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_252),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_349),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_528),
.Y(n_944)
);

BUFx10_ASAP7_75t_L g945 ( 
.A(n_268),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_673),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_700),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_529),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_274),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_122),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_290),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_35),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_103),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_138),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_65),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_616),
.Y(n_956)
);

BUFx10_ASAP7_75t_L g957 ( 
.A(n_381),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_145),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_680),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_560),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_684),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_790),
.Y(n_962)
);

INVx1_ASAP7_75t_SL g963 ( 
.A(n_767),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_607),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_742),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_129),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_14),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_743),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_651),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_620),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_127),
.Y(n_971)
);

CKINVDCx16_ASAP7_75t_R g972 ( 
.A(n_519),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_620),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_801),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_47),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_559),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_286),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_662),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_498),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_241),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_749),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_79),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_367),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_596),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_727),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_95),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_633),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_209),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_191),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_659),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_66),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_776),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_594),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_151),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_212),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_607),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_583),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_105),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_781),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_8),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_738),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_367),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_548),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_207),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_376),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_593),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_152),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_333),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_733),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_274),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_665),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_289),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_382),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_657),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_575),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_22),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_783),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_762),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_728),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_770),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_635),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_472),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_308),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_101),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_282),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_493),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_256),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_690),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_660),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_773),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_664),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_771),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_754),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_480),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_672),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_361),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_168),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_729),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_409),
.Y(n_1039)
);

INVxp33_ASAP7_75t_SL g1040 ( 
.A(n_709),
.Y(n_1040)
);

BUFx8_ASAP7_75t_SL g1041 ( 
.A(n_160),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_462),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_100),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_757),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_612),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_337),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_261),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_402),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_63),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_366),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_2),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_666),
.Y(n_1052)
);

CKINVDCx16_ASAP7_75t_R g1053 ( 
.A(n_764),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_461),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_375),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_770),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_23),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_756),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_335),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_582),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_667),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_525),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_636),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_5),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_321),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_376),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_114),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_270),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_591),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_556),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_384),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_814),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_567),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_301),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_237),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_260),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_741),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_739),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_351),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_87),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_681),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_360),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_476),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_204),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_755),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_628),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_325),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_347),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_806),
.Y(n_1089)
);

BUFx10_ASAP7_75t_L g1090 ( 
.A(n_793),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_651),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_335),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_713),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_360),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_221),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_44),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_676),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_340),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_458),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_488),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_796),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_195),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_772),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_175),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_538),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_217),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_738),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_642),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_551),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_211),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_285),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_592),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_604),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_103),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_163),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_36),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_748),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_334),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_544),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_293),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_31),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_112),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_110),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_785),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_353),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_690),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_252),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_337),
.Y(n_1128)
);

CKINVDCx16_ASAP7_75t_R g1129 ( 
.A(n_746),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_282),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_251),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_747),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_295),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_294),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_325),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_306),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_757),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_27),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_457),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_755),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_52),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_624),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_718),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_509),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_780),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_782),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_715),
.Y(n_1147)
);

CKINVDCx14_ASAP7_75t_R g1148 ( 
.A(n_448),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_35),
.Y(n_1149)
);

CKINVDCx16_ASAP7_75t_R g1150 ( 
.A(n_712),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_185),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_692),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_514),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_323),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_764),
.Y(n_1155)
);

CKINVDCx16_ASAP7_75t_R g1156 ( 
.A(n_73),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_556),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_391),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_192),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_109),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_180),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_212),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_88),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_9),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_125),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_773),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_401),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_445),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_137),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_263),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_4),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_292),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_759),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_313),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_765),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_566),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_744),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_260),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_202),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_160),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_740),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_7),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_424),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_815),
.Y(n_1184)
);

CKINVDCx14_ASAP7_75t_R g1185 ( 
.A(n_508),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_13),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_31),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_745),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_167),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_52),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_721),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_371),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_595),
.Y(n_1193)
);

BUFx10_ASAP7_75t_L g1194 ( 
.A(n_373),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_381),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_2),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_419),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_236),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_291),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_769),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_46),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_535),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_248),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_97),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_312),
.Y(n_1205)
);

CKINVDCx12_ASAP7_75t_R g1206 ( 
.A(n_608),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_36),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_728),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_351),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_741),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_661),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_686),
.Y(n_1212)
);

CKINVDCx16_ASAP7_75t_R g1213 ( 
.A(n_382),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_405),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_269),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_740),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_258),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_736),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_407),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_362),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_363),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_525),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_606),
.Y(n_1223)
);

INVxp67_ASAP7_75t_SL g1224 ( 
.A(n_162),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_518),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_32),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_178),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_255),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_618),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_170),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_276),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_74),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_365),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_658),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_247),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_761),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_232),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_69),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_598),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_112),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_539),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_574),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_782),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_289),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_402),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_752),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_123),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_345),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_669),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_406),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_19),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_768),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_406),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_763),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_297),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_270),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_587),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_186),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_704),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_369),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_244),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_811),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_24),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_283),
.Y(n_1264)
);

CKINVDCx16_ASAP7_75t_R g1265 ( 
.A(n_64),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_735),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_336),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_268),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_779),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_731),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_350),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_805),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_319),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_677),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_595),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_70),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_797),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_20),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_557),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_548),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_98),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_117),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_296),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_497),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_429),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_404),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_248),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_241),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_710),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_694),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_574),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_732),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_813),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_761),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_463),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_751),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_222),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_694),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_73),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_787),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_243),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_766),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_38),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_640),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_750),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_120),
.Y(n_1306)
);

CKINVDCx16_ASAP7_75t_R g1307 ( 
.A(n_768),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_408),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_721),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_526),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_493),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_795),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_447),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_265),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_666),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_529),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_730),
.Y(n_1317)
);

BUFx10_ASAP7_75t_L g1318 ( 
.A(n_63),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_124),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_490),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_128),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_28),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_637),
.Y(n_1323)
);

CKINVDCx16_ASAP7_75t_R g1324 ( 
.A(n_242),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_807),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_318),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_313),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_167),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_586),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_732),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_717),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_705),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_432),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_438),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_726),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_746),
.Y(n_1336)
);

CKINVDCx16_ASAP7_75t_R g1337 ( 
.A(n_532),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_153),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_458),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_316),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_87),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_775),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_0),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_236),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_650),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_195),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_743),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_400),
.Y(n_1348)
);

BUFx2_ASAP7_75t_SL g1349 ( 
.A(n_21),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_149),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_224),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_778),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_816),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_420),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_533),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_92),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_225),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_783),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_669),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_490),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_758),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1115),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1041),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1115),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_868),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1115),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_860),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_870),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1186),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_1186),
.Y(n_1370)
);

INVxp67_ASAP7_75t_L g1371 ( 
.A(n_982),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_879),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_1186),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1148),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_843),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_843),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_849),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_849),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_861),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1293),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_861),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_952),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_990),
.B(n_0),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_952),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1046),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1046),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1185),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1071),
.Y(n_1388)
);

INVxp33_ASAP7_75t_SL g1389 ( 
.A(n_1321),
.Y(n_1389)
);

CKINVDCx16_ASAP7_75t_R g1390 ( 
.A(n_897),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_839),
.Y(n_1391)
);

INVxp33_ASAP7_75t_L g1392 ( 
.A(n_1070),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1071),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_972),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1085),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1085),
.Y(n_1396)
);

CKINVDCx20_ASAP7_75t_R g1397 ( 
.A(n_925),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1112),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1112),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1217),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1217),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1222),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1222),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_827),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_817),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_819),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1053),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_822),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_828),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1132),
.Y(n_1410)
);

INVxp33_ASAP7_75t_L g1411 ( 
.A(n_1153),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_827),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1129),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_829),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_833),
.Y(n_1415)
);

INVxp67_ASAP7_75t_L g1416 ( 
.A(n_1250),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1150),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_844),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_974),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1262),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_847),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1156),
.Y(n_1422)
);

INVx1_ASAP7_75t_SL g1423 ( 
.A(n_859),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1291),
.B(n_1),
.Y(n_1424)
);

INVxp67_ASAP7_75t_SL g1425 ( 
.A(n_857),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_862),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1299),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_851),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_857),
.Y(n_1429)
);

INVxp33_ASAP7_75t_L g1430 ( 
.A(n_852),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_855),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_867),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_869),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_874),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1164),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1213),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_878),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1090),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_882),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_893),
.Y(n_1440)
);

INVxp33_ASAP7_75t_L g1441 ( 
.A(n_896),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1265),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_903),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_910),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1307),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_911),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_912),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_915),
.Y(n_1448)
);

CKINVDCx14_ASAP7_75t_R g1449 ( 
.A(n_1090),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1132),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_924),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_928),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_931),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1324),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_934),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_935),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_937),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_940),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1337),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_944),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_889),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_914),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_900),
.Y(n_1463)
);

BUFx5_ASAP7_75t_L g1464 ( 
.A(n_871),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_948),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_949),
.Y(n_1466)
);

INVxp33_ASAP7_75t_SL g1467 ( 
.A(n_820),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_916),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_950),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_954),
.Y(n_1470)
);

INVxp67_ASAP7_75t_SL g1471 ( 
.A(n_888),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_958),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_965),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_966),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_968),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_917),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_973),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_976),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_978),
.Y(n_1479)
);

INVxp33_ASAP7_75t_SL g1480 ( 
.A(n_820),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_979),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_980),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_888),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_913),
.Y(n_1484)
);

INVxp67_ASAP7_75t_SL g1485 ( 
.A(n_901),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1040),
.B(n_3),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_918),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1132),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_933),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1206),
.Y(n_1490)
);

INVxp67_ASAP7_75t_SL g1491 ( 
.A(n_901),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_989),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1090),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1132),
.Y(n_1494)
);

CKINVDCx14_ASAP7_75t_R g1495 ( 
.A(n_945),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_946),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_991),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1132),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_955),
.Y(n_1499)
);

INVxp33_ASAP7_75t_SL g1500 ( 
.A(n_821),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_992),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_995),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1410),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1450),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1488),
.Y(n_1505)
);

AND2x6_ASAP7_75t_L g1506 ( 
.A(n_1438),
.B(n_933),
.Y(n_1506)
);

BUFx8_ASAP7_75t_SL g1507 ( 
.A(n_1426),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1494),
.Y(n_1508)
);

INVx5_ASAP7_75t_L g1509 ( 
.A(n_1489),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1362),
.A2(n_1072),
.B(n_962),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1498),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1364),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1366),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1391),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1489),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1369),
.A2(n_1101),
.B(n_823),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1489),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1489),
.Y(n_1518)
);

NOR2x1_ASAP7_75t_L g1519 ( 
.A(n_1493),
.B(n_1380),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1382),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1397),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1405),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1449),
.B(n_945),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1369),
.A2(n_1101),
.B(n_823),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1365),
.Y(n_1525)
);

INVx5_ASAP7_75t_L g1526 ( 
.A(n_1367),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1370),
.A2(n_1325),
.B(n_1089),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1370),
.A2(n_1000),
.B(n_971),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1373),
.B(n_1184),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1373),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1464),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1464),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1464),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1393),
.B(n_1272),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1423),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1464),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1406),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1393),
.B(n_1463),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1464),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1408),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1368),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1495),
.B(n_945),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1409),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1414),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1464),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1375),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1376),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1377),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1372),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1415),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1378),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1371),
.A2(n_1416),
.B1(n_1389),
.B2(n_1411),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1418),
.Y(n_1553)
);

INVx6_ASAP7_75t_L g1554 ( 
.A(n_1390),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1379),
.B(n_883),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1371),
.A2(n_970),
.B1(n_987),
.B2(n_956),
.Y(n_1556)
);

CKINVDCx6p67_ASAP7_75t_R g1557 ( 
.A(n_1374),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1381),
.Y(n_1558)
);

AOI22x1_ASAP7_75t_SL g1559 ( 
.A1(n_1461),
.A2(n_1024),
.B1(n_1045),
.B2(n_1020),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1421),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1384),
.Y(n_1561)
);

CKINVDCx6p67_ASAP7_75t_R g1562 ( 
.A(n_1387),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1463),
.B(n_900),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1385),
.A2(n_1388),
.B(n_1386),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1428),
.Y(n_1565)
);

INVx5_ASAP7_75t_L g1566 ( 
.A(n_1427),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1416),
.B(n_907),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1395),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1396),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1431),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1394),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1462),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1392),
.A2(n_1110),
.B1(n_1134),
.B2(n_1077),
.Y(n_1573)
);

INVx5_ASAP7_75t_L g1574 ( 
.A(n_1430),
.Y(n_1574)
);

OA21x2_ASAP7_75t_L g1575 ( 
.A1(n_1432),
.A2(n_1000),
.B(n_971),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1398),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1441),
.B(n_957),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1399),
.A2(n_1401),
.B(n_1400),
.Y(n_1578)
);

BUFx12f_ASAP7_75t_L g1579 ( 
.A(n_1363),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1468),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1490),
.B(n_907),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1433),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1502),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1402),
.B(n_883),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1501),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1434),
.A2(n_1076),
.B(n_1050),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1437),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1403),
.A2(n_1076),
.B(n_1050),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1467),
.B(n_1277),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1439),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1440),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1484),
.A2(n_1229),
.B1(n_1273),
.B2(n_1210),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1404),
.B(n_1004),
.Y(n_1593)
);

OA21x2_ASAP7_75t_L g1594 ( 
.A1(n_1443),
.A2(n_1161),
.B(n_1139),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1444),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1446),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1407),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1419),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1420),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1447),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1448),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1480),
.A2(n_1500),
.B1(n_1417),
.B2(n_1422),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1451),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1452),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1476),
.B(n_1277),
.Y(n_1605)
);

BUFx12f_ASAP7_75t_L g1606 ( 
.A(n_1413),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1435),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1453),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1487),
.B(n_1300),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1455),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1456),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1457),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1404),
.B(n_957),
.Y(n_1613)
);

AND2x6_ASAP7_75t_L g1614 ( 
.A(n_1458),
.B(n_1139),
.Y(n_1614)
);

BUFx8_ASAP7_75t_L g1615 ( 
.A(n_1383),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1460),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1436),
.A2(n_1286),
.B1(n_1141),
.B2(n_1173),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1412),
.B(n_957),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1465),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1466),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1469),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1470),
.Y(n_1622)
);

OAI22x1_ASAP7_75t_L g1623 ( 
.A1(n_1442),
.A2(n_906),
.B1(n_922),
.B2(n_818),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1472),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1412),
.B(n_1194),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1473),
.Y(n_1626)
);

AND2x6_ASAP7_75t_L g1627 ( 
.A(n_1474),
.B(n_1475),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1588),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1512),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1512),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1515),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1546),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1509),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1547),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1515),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1518),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1548),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1505),
.Y(n_1638)
);

AND2x2_ASAP7_75t_SL g1639 ( 
.A(n_1523),
.B(n_1424),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1551),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1520),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1577),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1535),
.Y(n_1643)
);

AND2x6_ASAP7_75t_L g1644 ( 
.A(n_1542),
.B(n_1486),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1538),
.B(n_1574),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1558),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1561),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1531),
.B(n_1425),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1568),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1517),
.Y(n_1650)
);

INVx5_ASAP7_75t_L g1651 ( 
.A(n_1627),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1569),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1556),
.A2(n_1499),
.B1(n_1496),
.B2(n_1169),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1576),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1508),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1596),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1600),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1601),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1530),
.B(n_1425),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1572),
.B(n_1300),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1603),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1531),
.B(n_1429),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1517),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1513),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1611),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1612),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1510),
.A2(n_1478),
.B(n_1477),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1626),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1560),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1532),
.B(n_1429),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1528),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1532),
.B(n_1471),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1513),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1560),
.Y(n_1674)
);

CKINVDCx6p67_ASAP7_75t_R g1675 ( 
.A(n_1579),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1583),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1522),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1522),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1545),
.B(n_1471),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1583),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1574),
.Y(n_1681)
);

INVxp33_ASAP7_75t_L g1682 ( 
.A(n_1552),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1585),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1585),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1590),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1564),
.A2(n_1481),
.B(n_1479),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1574),
.B(n_1445),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1590),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1538),
.B(n_1454),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1591),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1591),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1595),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1522),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1528),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1595),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1593),
.B(n_1483),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1509),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1530),
.B(n_1483),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1545),
.B(n_1485),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1537),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1608),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1608),
.Y(n_1702)
);

AND2x2_ASAP7_75t_SL g1703 ( 
.A(n_1572),
.B(n_1239),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1621),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1621),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1540),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1620),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1537),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1537),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1533),
.B(n_1485),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1543),
.Y(n_1711)
);

INVx6_ASAP7_75t_L g1712 ( 
.A(n_1526),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1624),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1509),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1543),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1543),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1544),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1544),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1544),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1589),
.A2(n_1459),
.B1(n_1040),
.B2(n_986),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1593),
.B(n_1491),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1613),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1541),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1550),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1550),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1550),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1553),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1553),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1605),
.B(n_1353),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1553),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1618),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1565),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1578),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1571),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1565),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1536),
.B(n_1491),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1565),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1625),
.B(n_1482),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1570),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1570),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1570),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1582),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1539),
.B(n_1492),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1582),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1582),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1587),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1587),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1587),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1604),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1604),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1604),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1610),
.Y(n_1752)
);

OA21x2_ASAP7_75t_L g1753 ( 
.A1(n_1529),
.A2(n_1497),
.B(n_1001),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1627),
.B(n_1157),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1566),
.B(n_1194),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1610),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1610),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1616),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1616),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1616),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1567),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1503),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1619),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1503),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1682),
.A2(n_1627),
.B1(n_1580),
.B2(n_1506),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1696),
.B(n_1506),
.Y(n_1766)
);

INVx4_ASAP7_75t_L g1767 ( 
.A(n_1712),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1696),
.B(n_1506),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_L g1769 ( 
.A(n_1644),
.B(n_1627),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1723),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1669),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1734),
.Y(n_1772)
);

INVx5_ASAP7_75t_L g1773 ( 
.A(n_1712),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1677),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1689),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1675),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1674),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1676),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1703),
.B(n_1602),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1645),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1680),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1703),
.B(n_1534),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1683),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1643),
.B(n_1525),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1682),
.A2(n_1527),
.B1(n_1567),
.B2(n_1516),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1641),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1642),
.A2(n_1224),
.B1(n_1607),
.B2(n_885),
.Y(n_1787)
);

BUFx2_ASAP7_75t_L g1788 ( 
.A(n_1643),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1762),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1639),
.B(n_1526),
.Y(n_1790)
);

BUFx10_ASAP7_75t_L g1791 ( 
.A(n_1712),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1753),
.A2(n_1527),
.B1(n_1516),
.B2(n_1524),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1721),
.B(n_1506),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1684),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1762),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1653),
.Y(n_1796)
);

NAND3xp33_ASAP7_75t_L g1797 ( 
.A(n_1642),
.B(n_1729),
.C(n_1720),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1645),
.B(n_1526),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1687),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1721),
.Y(n_1800)
);

INVx4_ASAP7_75t_L g1801 ( 
.A(n_1651),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1685),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1639),
.B(n_1549),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1764),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1659),
.B(n_1698),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1729),
.B(n_1609),
.C(n_1615),
.Y(n_1806)
);

NOR3xp33_ASAP7_75t_L g1807 ( 
.A(n_1660),
.B(n_1573),
.C(n_1597),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1660),
.B(n_1554),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1688),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1764),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1755),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1638),
.Y(n_1812)
);

BUFx3_ASAP7_75t_L g1813 ( 
.A(n_1656),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1677),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1677),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1651),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1753),
.A2(n_1524),
.B1(n_1615),
.B2(n_1586),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1761),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1722),
.B(n_1554),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1659),
.B(n_1581),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1686),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1761),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1722),
.B(n_1566),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1709),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1698),
.B(n_1581),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1638),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1655),
.Y(n_1827)
);

INVxp33_ASAP7_75t_L g1828 ( 
.A(n_1738),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1657),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1731),
.B(n_1566),
.Y(n_1830)
);

BUFx4f_ASAP7_75t_L g1831 ( 
.A(n_1644),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1686),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1731),
.B(n_1555),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1709),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1667),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1648),
.B(n_1619),
.Y(n_1836)
);

AND2x6_ASAP7_75t_L g1837 ( 
.A(n_1733),
.B(n_1563),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1690),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1700),
.B(n_1606),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1700),
.B(n_1514),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1681),
.B(n_1584),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1648),
.B(n_1670),
.C(n_1662),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_L g1843 ( 
.A(n_1644),
.B(n_1157),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1691),
.Y(n_1844)
);

NAND2x1p5_ASAP7_75t_L g1845 ( 
.A(n_1681),
.B(n_1519),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1662),
.B(n_1619),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_SL g1847 ( 
.A(n_1706),
.B(n_1192),
.C(n_1178),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1644),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1711),
.B(n_1521),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1692),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1709),
.Y(n_1851)
);

INVx5_ASAP7_75t_L g1852 ( 
.A(n_1717),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1695),
.Y(n_1853)
);

INVx4_ASAP7_75t_L g1854 ( 
.A(n_1651),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1701),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1658),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1711),
.B(n_1598),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1724),
.B(n_1599),
.Y(n_1858)
);

INVx8_ASAP7_75t_L g1859 ( 
.A(n_1644),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1670),
.B(n_1622),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1655),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1707),
.B(n_1617),
.Y(n_1862)
);

CKINVDCx14_ASAP7_75t_R g1863 ( 
.A(n_1717),
.Y(n_1863)
);

INVx4_ASAP7_75t_L g1864 ( 
.A(n_1651),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1724),
.B(n_1557),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1717),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1735),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1702),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1735),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1664),
.Y(n_1870)
);

AND2x2_ASAP7_75t_SL g1871 ( 
.A(n_1735),
.B(n_1563),
.Y(n_1871)
);

BUFx3_ASAP7_75t_L g1872 ( 
.A(n_1661),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1704),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1672),
.B(n_1622),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1665),
.B(n_1562),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1705),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1713),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1749),
.Y(n_1878)
);

INVx8_ASAP7_75t_L g1879 ( 
.A(n_1749),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1749),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1763),
.B(n_1622),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1763),
.B(n_1507),
.Y(n_1882)
);

NOR2x1p5_ASAP7_75t_L g1883 ( 
.A(n_1629),
.B(n_821),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1666),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1671),
.A2(n_1586),
.B1(n_1594),
.B2(n_1575),
.Y(n_1885)
);

INVx5_ASAP7_75t_L g1886 ( 
.A(n_1671),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1672),
.B(n_1312),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1630),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1679),
.B(n_1614),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1673),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1679),
.B(n_1614),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1632),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1699),
.B(n_1614),
.Y(n_1893)
);

INVx2_ASAP7_75t_SL g1894 ( 
.A(n_1678),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1634),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1699),
.B(n_1312),
.Y(n_1896)
);

NOR2x1p5_ASAP7_75t_L g1897 ( 
.A(n_1668),
.B(n_824),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1710),
.B(n_1353),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1694),
.A2(n_1594),
.B1(n_1575),
.B2(n_1614),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1637),
.B(n_1592),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1631),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1640),
.Y(n_1902)
);

INVx4_ASAP7_75t_L g1903 ( 
.A(n_1633),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1710),
.B(n_963),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1646),
.B(n_1647),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1649),
.B(n_1623),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1652),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1654),
.B(n_997),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1743),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1743),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1694),
.A2(n_1264),
.B1(n_1271),
.B2(n_1252),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1736),
.B(n_824),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1736),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1715),
.B(n_1004),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1716),
.B(n_1013),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1719),
.B(n_1352),
.Y(n_1916)
);

NAND2xp33_ASAP7_75t_L g1917 ( 
.A(n_1650),
.B(n_1157),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1663),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1730),
.B(n_1013),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1635),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1693),
.A2(n_1330),
.B1(n_1346),
.B2(n_1301),
.Y(n_1921)
);

AND2x6_ASAP7_75t_L g1922 ( 
.A(n_1733),
.B(n_1161),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1708),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1718),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1737),
.B(n_1002),
.Y(n_1925)
);

INVxp67_ASAP7_75t_SL g1926 ( 
.A(n_1800),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1805),
.B(n_1739),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_SL g1928 ( 
.A(n_1776),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1904),
.B(n_1740),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1788),
.B(n_1725),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1779),
.A2(n_1742),
.B1(n_1746),
.B2(n_1744),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1784),
.B(n_1726),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1820),
.B(n_1741),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1765),
.B(n_1727),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1871),
.B(n_1728),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1772),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1825),
.B(n_1909),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1771),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1819),
.B(n_1732),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1786),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1879),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1910),
.B(n_1747),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1777),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1778),
.Y(n_1944)
);

AND2x4_ASAP7_75t_SL g1945 ( 
.A(n_1791),
.B(n_1745),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1775),
.B(n_1748),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1811),
.B(n_1770),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1828),
.B(n_1752),
.Y(n_1948)
);

INVx2_ASAP7_75t_SL g1949 ( 
.A(n_1798),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1803),
.B(n_1756),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1913),
.B(n_1757),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1877),
.B(n_1758),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1781),
.B(n_1759),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1783),
.B(n_1794),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1789),
.Y(n_1955)
);

INVxp33_ASAP7_75t_L g1956 ( 
.A(n_1840),
.Y(n_1956)
);

INVx3_ASAP7_75t_L g1957 ( 
.A(n_1851),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1802),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1809),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1818),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1795),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1851),
.Y(n_1962)
);

A2O1A1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1831),
.A2(n_1797),
.B(n_1843),
.C(n_1782),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1838),
.B(n_1844),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1831),
.B(n_1750),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1851),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1850),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1853),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1862),
.B(n_1760),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1804),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1855),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1868),
.B(n_1751),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1822),
.B(n_1559),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1873),
.B(n_1754),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1808),
.B(n_1559),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1876),
.B(n_1754),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1823),
.B(n_1636),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1916),
.B(n_1194),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1810),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1888),
.B(n_1633),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1830),
.B(n_1008),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1773),
.B(n_1697),
.Y(n_1982)
);

INVx8_ASAP7_75t_L g1983 ( 
.A(n_1879),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1848),
.A2(n_887),
.B1(n_959),
.B2(n_881),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1773),
.B(n_1697),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1905),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1812),
.Y(n_1987)
);

O2A1O1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1833),
.A2(n_1787),
.B(n_1912),
.C(n_1896),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1773),
.B(n_1714),
.Y(n_1989)
);

O2A1O1Ixp33_ASAP7_75t_L g1990 ( 
.A1(n_1887),
.A2(n_1235),
.B(n_1248),
.C(n_1211),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1866),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1836),
.B(n_1714),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1826),
.Y(n_1993)
);

BUFx5_ASAP7_75t_L g1994 ( 
.A(n_1821),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1846),
.B(n_1019),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1860),
.B(n_1874),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1767),
.B(n_1628),
.Y(n_1997)
);

INVx4_ASAP7_75t_L g1998 ( 
.A(n_1859),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1769),
.A2(n_1628),
.B(n_1087),
.Y(n_1999)
);

BUFx3_ASAP7_75t_L g2000 ( 
.A(n_1798),
.Y(n_2000)
);

INVxp67_ASAP7_75t_L g2001 ( 
.A(n_1849),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_SL g2002 ( 
.A(n_1767),
.B(n_825),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1766),
.B(n_1019),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1768),
.B(n_1087),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1793),
.B(n_1093),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1799),
.B(n_1074),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1837),
.A2(n_1246),
.B1(n_1270),
.B2(n_1182),
.Y(n_2007)
);

INVx8_ASAP7_75t_L g2008 ( 
.A(n_1859),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1863),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1842),
.B(n_1093),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1807),
.B(n_825),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1827),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1861),
.Y(n_2013)
);

AO22x2_ASAP7_75t_L g2014 ( 
.A1(n_1847),
.A2(n_1349),
.B1(n_1296),
.B2(n_1189),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1785),
.B(n_1146),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1884),
.B(n_826),
.Y(n_2016)
);

BUFx2_ASAP7_75t_L g2017 ( 
.A(n_1780),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1892),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1895),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1837),
.B(n_1146),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1870),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1890),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1837),
.B(n_1189),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_1857),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1791),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1900),
.B(n_1207),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1883),
.B(n_1005),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1858),
.B(n_826),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1837),
.B(n_1190),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1907),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1918),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1790),
.B(n_1875),
.Y(n_2032)
);

OAI22x1_ASAP7_75t_SL g2033 ( 
.A1(n_1796),
.A2(n_831),
.B1(n_832),
.B2(n_830),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1908),
.B(n_1190),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1908),
.B(n_1191),
.Y(n_2035)
);

CKINVDCx20_ASAP7_75t_R g2036 ( 
.A(n_1882),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1852),
.B(n_830),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1852),
.B(n_831),
.Y(n_2038)
);

OAI22x1_ASAP7_75t_R g2039 ( 
.A1(n_1897),
.A2(n_834),
.B1(n_835),
.B2(n_832),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1852),
.B(n_834),
.Y(n_2040)
);

INVx2_ASAP7_75t_SL g2041 ( 
.A(n_1845),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1901),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1920),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1924),
.B(n_1191),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1922),
.A2(n_1216),
.B1(n_1345),
.B2(n_1196),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1914),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1911),
.A2(n_1345),
.B1(n_1196),
.B2(n_1216),
.Y(n_2047)
);

NOR2x1p5_ASAP7_75t_L g2048 ( 
.A(n_1806),
.B(n_1359),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1925),
.B(n_835),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1866),
.B(n_836),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1921),
.B(n_1865),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1866),
.B(n_836),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1839),
.B(n_837),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_L g2054 ( 
.A(n_1922),
.B(n_837),
.Y(n_2054)
);

OAI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1813),
.A2(n_840),
.B1(n_841),
.B2(n_838),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1915),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1903),
.B(n_838),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_1829),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1925),
.B(n_840),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1919),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1856),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1906),
.A2(n_1207),
.B1(n_1318),
.B2(n_1226),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1872),
.B(n_841),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1817),
.A2(n_1207),
.B1(n_1318),
.B2(n_1226),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1903),
.B(n_842),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1902),
.B(n_1318),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1923),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1869),
.B(n_842),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1841),
.B(n_845),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1834),
.B(n_845),
.Y(n_2070)
);

NAND2x1p5_ASAP7_75t_L g2071 ( 
.A(n_1878),
.B(n_1504),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1923),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1894),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1922),
.A2(n_920),
.B1(n_921),
.B2(n_919),
.Y(n_2074)
);

O2A1O1Ixp5_ASAP7_75t_L g2075 ( 
.A1(n_1898),
.A2(n_1835),
.B(n_1881),
.C(n_1832),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1774),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1774),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1878),
.B(n_846),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1814),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1801),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1814),
.Y(n_2081)
);

NOR2xp33_ASAP7_75t_L g2082 ( 
.A(n_1886),
.B(n_1815),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_1886),
.B(n_1356),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1815),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1886),
.B(n_846),
.Y(n_2085)
);

BUFx8_ASAP7_75t_L g2086 ( 
.A(n_1922),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1889),
.B(n_848),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1824),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1824),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1867),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1867),
.B(n_864),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1880),
.B(n_864),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1880),
.B(n_848),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1891),
.B(n_1359),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1893),
.A2(n_853),
.B1(n_854),
.B2(n_850),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1899),
.B(n_1792),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_L g2097 ( 
.A(n_1835),
.B(n_850),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1885),
.B(n_853),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1938),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_1983),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2043),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1937),
.B(n_2001),
.Y(n_2102)
);

AOI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_1947),
.A2(n_1917),
.B1(n_926),
.B2(n_927),
.Y(n_2103)
);

INVx3_ASAP7_75t_L g2104 ( 
.A(n_1983),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_1998),
.B(n_1801),
.Y(n_2105)
);

INVx1_ASAP7_75t_SL g2106 ( 
.A(n_1936),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2024),
.B(n_1986),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1943),
.Y(n_2108)
);

OR2x6_ASAP7_75t_L g2109 ( 
.A(n_2009),
.B(n_1816),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1955),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1956),
.B(n_1816),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1969),
.B(n_854),
.Y(n_2112)
);

OAI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_2075),
.A2(n_1927),
.B(n_1999),
.Y(n_2113)
);

NOR3xp33_ASAP7_75t_L g2114 ( 
.A(n_2053),
.B(n_1011),
.C(n_1010),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_1996),
.A2(n_1832),
.B(n_1821),
.Y(n_2115)
);

NOR3xp33_ASAP7_75t_L g2116 ( 
.A(n_2011),
.B(n_1361),
.C(n_1350),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1983),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1944),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1941),
.B(n_2007),
.Y(n_2119)
);

AOI22xp33_ASAP7_75t_SL g2120 ( 
.A1(n_2051),
.A2(n_858),
.B1(n_863),
.B2(n_856),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1981),
.B(n_856),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1958),
.Y(n_2122)
);

BUFx3_ASAP7_75t_L g2123 ( 
.A(n_1941),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1959),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1961),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1941),
.B(n_1854),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1967),
.Y(n_2127)
);

INVx3_ASAP7_75t_L g2128 ( 
.A(n_1928),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_1998),
.B(n_1854),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1968),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1970),
.Y(n_2131)
);

NAND2x1p5_ASAP7_75t_L g2132 ( 
.A(n_2000),
.B(n_1864),
.Y(n_2132)
);

AOI22xp33_ASAP7_75t_L g2133 ( 
.A1(n_2026),
.A2(n_863),
.B1(n_865),
.B2(n_858),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1971),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1954),
.B(n_865),
.Y(n_2135)
);

AOI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2036),
.A2(n_2032),
.B1(n_2007),
.B2(n_1973),
.Y(n_2136)
);

AOI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_1960),
.A2(n_929),
.B1(n_930),
.B2(n_923),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_1926),
.B(n_866),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_2006),
.B(n_866),
.Y(n_2139)
);

OAI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_2074),
.A2(n_2045),
.B1(n_2059),
.B2(n_2049),
.Y(n_2140)
);

AOI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_1975),
.A2(n_873),
.B1(n_875),
.B2(n_872),
.Y(n_2141)
);

INVx4_ASAP7_75t_L g2142 ( 
.A(n_2008),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1964),
.B(n_1946),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1978),
.B(n_872),
.Y(n_2144)
);

NAND2x1p5_ASAP7_75t_L g2145 ( 
.A(n_1949),
.B(n_1864),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2018),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_2008),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1979),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2031),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_2008),
.Y(n_2150)
);

BUFx6f_ASAP7_75t_L g2151 ( 
.A(n_2077),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_2028),
.B(n_873),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2094),
.A2(n_2087),
.B1(n_1976),
.B2(n_1974),
.Y(n_2153)
);

OR2x2_ASAP7_75t_SL g2154 ( 
.A(n_2033),
.B(n_2039),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_2025),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_L g2156 ( 
.A(n_1994),
.B(n_875),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2019),
.B(n_876),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_SL g2158 ( 
.A1(n_2014),
.A2(n_877),
.B1(n_880),
.B2(n_876),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_SL g2159 ( 
.A(n_1928),
.B(n_2086),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2030),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_2016),
.B(n_877),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_2017),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1929),
.B(n_880),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_2046),
.B(n_884),
.Y(n_2164)
);

AOI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_2083),
.A2(n_936),
.B1(n_938),
.B2(n_932),
.Y(n_2165)
);

AND2x6_ASAP7_75t_SL g2166 ( 
.A(n_2027),
.B(n_1012),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2097),
.A2(n_941),
.B1(n_942),
.B2(n_939),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_L g2168 ( 
.A(n_1994),
.B(n_884),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_2058),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1987),
.Y(n_2170)
);

BUFx3_ASAP7_75t_L g2171 ( 
.A(n_2061),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_1957),
.Y(n_2172)
);

AO22x1_ASAP7_75t_L g2173 ( 
.A1(n_2086),
.A2(n_890),
.B1(n_891),
.B2(n_886),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2021),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_2074),
.B(n_886),
.Y(n_2175)
);

AOI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2047),
.A2(n_891),
.B1(n_892),
.B2(n_890),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1933),
.B(n_892),
.Y(n_2177)
);

OR2x6_ASAP7_75t_L g2178 ( 
.A(n_2041),
.B(n_1172),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1950),
.B(n_894),
.Y(n_2179)
);

CKINVDCx20_ASAP7_75t_R g2180 ( 
.A(n_2066),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_1945),
.B(n_1014),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1993),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2014),
.A2(n_895),
.B1(n_898),
.B2(n_894),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2091),
.B(n_895),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1948),
.B(n_898),
.Y(n_2185)
);

BUFx4f_ASAP7_75t_L g2186 ( 
.A(n_2027),
.Y(n_2186)
);

OR2x6_ASAP7_75t_L g2187 ( 
.A(n_2048),
.B(n_1172),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2012),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2013),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2056),
.B(n_2060),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_SL g2191 ( 
.A1(n_2045),
.A2(n_902),
.B1(n_904),
.B2(n_899),
.Y(n_2191)
);

BUFx3_ASAP7_75t_L g2192 ( 
.A(n_1957),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2022),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_2055),
.B(n_1963),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_2064),
.A2(n_902),
.B1(n_904),
.B2(n_899),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1953),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1972),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_2068),
.Y(n_2198)
);

BUFx6f_ASAP7_75t_L g2199 ( 
.A(n_1962),
.Y(n_2199)
);

A2O1A1Ixp33_ASAP7_75t_L g2200 ( 
.A1(n_1988),
.A2(n_1237),
.B(n_1239),
.C(n_1228),
.Y(n_2200)
);

INVx3_ASAP7_75t_L g2201 ( 
.A(n_1962),
.Y(n_2201)
);

OAI22xp33_ASAP7_75t_L g2202 ( 
.A1(n_2063),
.A2(n_908),
.B1(n_909),
.B2(n_905),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1977),
.B(n_1952),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1940),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1942),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2092),
.B(n_905),
.Y(n_2206)
);

INVx2_ASAP7_75t_SL g2207 ( 
.A(n_1930),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_1966),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_2085),
.B(n_1966),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1951),
.B(n_908),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2042),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2072),
.Y(n_2212)
);

AND2x6_ASAP7_75t_L g2213 ( 
.A(n_2080),
.B(n_1991),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2034),
.B(n_909),
.Y(n_2214)
);

INVx2_ASAP7_75t_SL g2215 ( 
.A(n_2037),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_1939),
.B(n_1080),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2044),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2067),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_1991),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_1984),
.A2(n_947),
.B1(n_951),
.B2(n_943),
.Y(n_2220)
);

HB1xp67_ASAP7_75t_L g2221 ( 
.A(n_1932),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2035),
.B(n_1080),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_2073),
.B(n_1018),
.Y(n_2223)
);

AOI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_1935),
.A2(n_960),
.B1(n_961),
.B2(n_953),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2010),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_1997),
.A2(n_1237),
.B(n_1228),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_R g2227 ( 
.A(n_2054),
.B(n_1081),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1995),
.B(n_1081),
.Y(n_2228)
);

INVx4_ASAP7_75t_L g2229 ( 
.A(n_2080),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_2084),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_2089),
.Y(n_2231)
);

NAND2x1_ASAP7_75t_L g2232 ( 
.A(n_2076),
.B(n_1504),
.Y(n_2232)
);

NOR3xp33_ASAP7_75t_SL g2233 ( 
.A(n_2057),
.B(n_1083),
.C(n_1082),
.Y(n_2233)
);

NOR3xp33_ASAP7_75t_SL g2234 ( 
.A(n_2065),
.B(n_1083),
.C(n_1082),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2090),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_L g2236 ( 
.A(n_2078),
.B(n_1280),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2062),
.B(n_1280),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1980),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_2069),
.Y(n_2239)
);

OR2x2_ASAP7_75t_L g2240 ( 
.A(n_2070),
.B(n_1282),
.Y(n_2240)
);

INVx3_ASAP7_75t_L g2241 ( 
.A(n_2079),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2081),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2095),
.B(n_1282),
.Y(n_2243)
);

A2O1A1Ixp33_ASAP7_75t_L g2244 ( 
.A1(n_1990),
.A2(n_1281),
.B(n_1287),
.C(n_1263),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2088),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1992),
.B(n_1283),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1994),
.Y(n_2247)
);

NOR2xp67_ASAP7_75t_L g2248 ( 
.A(n_2020),
.B(n_1511),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_2038),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1994),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_2136),
.B(n_2082),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_2143),
.B(n_1931),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_2142),
.B(n_1985),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_2140),
.B(n_1994),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2102),
.B(n_2002),
.Y(n_2255)
);

NAND2xp33_ASAP7_75t_SL g2256 ( 
.A(n_2142),
.B(n_2227),
.Y(n_2256)
);

NAND2xp33_ASAP7_75t_SL g2257 ( 
.A(n_2100),
.B(n_2040),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2205),
.B(n_2003),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2153),
.B(n_2023),
.Y(n_2259)
);

NAND2xp33_ASAP7_75t_SL g2260 ( 
.A(n_2147),
.B(n_2050),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_2198),
.B(n_2029),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2196),
.B(n_2071),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2186),
.B(n_2098),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2107),
.B(n_2004),
.Y(n_2264)
);

NAND2xp33_ASAP7_75t_SL g2265 ( 
.A(n_2147),
.B(n_2052),
.Y(n_2265)
);

NAND2xp33_ASAP7_75t_SL g2266 ( 
.A(n_2147),
.B(n_2093),
.Y(n_2266)
);

NAND2xp33_ASAP7_75t_SL g2267 ( 
.A(n_2104),
.B(n_1283),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2239),
.B(n_2005),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2139),
.B(n_2015),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_2229),
.B(n_1965),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2229),
.B(n_1982),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_2172),
.B(n_1989),
.Y(n_2272)
);

NAND2xp33_ASAP7_75t_SL g2273 ( 
.A(n_2233),
.B(n_1284),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2172),
.B(n_1934),
.Y(n_2274)
);

NAND2xp33_ASAP7_75t_SL g2275 ( 
.A(n_2234),
.B(n_1284),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2190),
.B(n_2203),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_2172),
.B(n_2096),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2199),
.B(n_1358),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_2199),
.B(n_1358),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2184),
.B(n_1294),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2199),
.B(n_2208),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2197),
.B(n_1294),
.Y(n_2282)
);

NAND2xp33_ASAP7_75t_SL g2283 ( 
.A(n_2150),
.B(n_1295),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2121),
.B(n_1295),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_2119),
.B(n_1297),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2225),
.B(n_1297),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2201),
.B(n_1339),
.Y(n_2287)
);

NAND2xp33_ASAP7_75t_SL g2288 ( 
.A(n_2150),
.B(n_1298),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_2201),
.B(n_2217),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2171),
.B(n_1339),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_2117),
.B(n_1511),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2207),
.B(n_1340),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_2238),
.B(n_1340),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2151),
.B(n_1343),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2164),
.B(n_1298),
.Y(n_2295)
);

NAND2xp33_ASAP7_75t_SL g2296 ( 
.A(n_2155),
.B(n_1303),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2214),
.B(n_1303),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_2151),
.B(n_1343),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_2151),
.B(n_1344),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2194),
.B(n_1344),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_2180),
.B(n_1347),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2106),
.B(n_1347),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2219),
.B(n_1348),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2249),
.B(n_1348),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2179),
.B(n_1305),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_2223),
.B(n_1351),
.Y(n_2306)
);

NAND2xp33_ASAP7_75t_SL g2307 ( 
.A(n_2191),
.B(n_1305),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2223),
.B(n_1354),
.Y(n_2308)
);

NAND2xp33_ASAP7_75t_SL g2309 ( 
.A(n_2243),
.B(n_2215),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_2162),
.B(n_2169),
.Y(n_2310)
);

NAND2xp33_ASAP7_75t_SL g2311 ( 
.A(n_2135),
.B(n_1308),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2120),
.B(n_1354),
.Y(n_2312)
);

NAND2xp33_ASAP7_75t_SL g2313 ( 
.A(n_2163),
.B(n_1308),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2181),
.B(n_1356),
.Y(n_2314)
);

AND2x4_ASAP7_75t_L g2315 ( 
.A(n_2123),
.B(n_1022),
.Y(n_2315)
);

NAND2xp33_ASAP7_75t_SL g2316 ( 
.A(n_2105),
.B(n_1313),
.Y(n_2316)
);

NAND2xp33_ASAP7_75t_SL g2317 ( 
.A(n_2105),
.B(n_1313),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2177),
.B(n_1314),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_2181),
.B(n_1314),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2192),
.B(n_1328),
.Y(n_2320)
);

NAND2xp33_ASAP7_75t_SL g2321 ( 
.A(n_2129),
.B(n_1315),
.Y(n_2321)
);

NAND2xp33_ASAP7_75t_SL g2322 ( 
.A(n_2129),
.B(n_1315),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2241),
.B(n_1332),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2099),
.B(n_1332),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2108),
.B(n_1333),
.Y(n_2325)
);

NAND2xp33_ASAP7_75t_SL g2326 ( 
.A(n_2210),
.B(n_1320),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2118),
.B(n_2122),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_2124),
.B(n_1333),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_2127),
.B(n_1334),
.Y(n_2329)
);

NAND2xp33_ASAP7_75t_SL g2330 ( 
.A(n_2206),
.B(n_1320),
.Y(n_2330)
);

NAND2xp33_ASAP7_75t_L g2331 ( 
.A(n_2213),
.B(n_1322),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_2130),
.B(n_1334),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_2134),
.B(n_1335),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2146),
.B(n_1335),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_2160),
.B(n_1336),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2230),
.B(n_1336),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2231),
.B(n_1338),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2112),
.B(n_1322),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_2103),
.B(n_1338),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2133),
.B(n_1326),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2138),
.B(n_1351),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2247),
.B(n_2250),
.Y(n_2342)
);

NAND2xp33_ASAP7_75t_SL g2343 ( 
.A(n_2175),
.B(n_2141),
.Y(n_2343)
);

NAND2xp33_ASAP7_75t_SL g2344 ( 
.A(n_2157),
.B(n_1326),
.Y(n_2344)
);

NAND2xp33_ASAP7_75t_SL g2345 ( 
.A(n_2240),
.B(n_1327),
.Y(n_2345)
);

NAND2xp33_ASAP7_75t_SL g2346 ( 
.A(n_2228),
.B(n_1327),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2245),
.B(n_1355),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2158),
.B(n_1355),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2111),
.B(n_1328),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2159),
.B(n_964),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2221),
.B(n_967),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_SL g2352 ( 
.A(n_2235),
.B(n_969),
.Y(n_2352)
);

NAND2xp33_ASAP7_75t_SL g2353 ( 
.A(n_2144),
.B(n_1360),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2218),
.B(n_975),
.Y(n_2354)
);

NAND2xp33_ASAP7_75t_SL g2355 ( 
.A(n_2246),
.B(n_977),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2248),
.B(n_981),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2212),
.B(n_983),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2145),
.B(n_984),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2161),
.B(n_985),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2185),
.B(n_988),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_2242),
.B(n_993),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2236),
.B(n_994),
.Y(n_2362)
);

NAND2xp33_ASAP7_75t_SL g2363 ( 
.A(n_2222),
.B(n_996),
.Y(n_2363)
);

NAND2xp33_ASAP7_75t_SL g2364 ( 
.A(n_2195),
.B(n_998),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_2202),
.B(n_999),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2200),
.B(n_1003),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_2152),
.B(n_1006),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_2109),
.B(n_1027),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2101),
.B(n_2149),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2183),
.B(n_1007),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_2132),
.B(n_1009),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2216),
.B(n_1015),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2113),
.B(n_1016),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2128),
.B(n_1017),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2137),
.B(n_1021),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2237),
.B(n_1023),
.Y(n_2376)
);

NAND2xp33_ASAP7_75t_SL g2377 ( 
.A(n_2126),
.B(n_1025),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_2116),
.B(n_1026),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_2170),
.B(n_1030),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2182),
.B(n_1032),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_2188),
.B(n_1033),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2189),
.B(n_2211),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2178),
.B(n_1034),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2167),
.B(n_1035),
.Y(n_2384)
);

NAND2xp33_ASAP7_75t_SL g2385 ( 
.A(n_2176),
.B(n_1036),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2209),
.B(n_1039),
.Y(n_2386)
);

NAND2xp33_ASAP7_75t_SL g2387 ( 
.A(n_2232),
.B(n_1042),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2114),
.B(n_1044),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_2165),
.B(n_1047),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_2224),
.B(n_1048),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2178),
.B(n_1049),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2174),
.B(n_2193),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_2115),
.B(n_1051),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_2110),
.B(n_1055),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2204),
.B(n_1056),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_2109),
.B(n_1028),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2125),
.B(n_1057),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2131),
.B(n_1058),
.Y(n_2398)
);

NAND2xp33_ASAP7_75t_SL g2399 ( 
.A(n_2156),
.B(n_1062),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2148),
.B(n_2220),
.Y(n_2400)
);

NAND2xp33_ASAP7_75t_SL g2401 ( 
.A(n_2168),
.B(n_1063),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2213),
.B(n_1064),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_2213),
.B(n_1029),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2310),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2392),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2280),
.B(n_2187),
.Y(n_2406)
);

BUFx2_ASAP7_75t_L g2407 ( 
.A(n_2309),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2277),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_2301),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2382),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2276),
.B(n_2166),
.Y(n_2411)
);

HB1xp67_ASAP7_75t_L g2412 ( 
.A(n_2327),
.Y(n_2412)
);

AND2x2_ASAP7_75t_SL g2413 ( 
.A(n_2331),
.B(n_2154),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2269),
.B(n_2173),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2369),
.Y(n_2415)
);

A2O1A1Ixp33_ASAP7_75t_SL g2416 ( 
.A1(n_2295),
.A2(n_2318),
.B(n_2305),
.C(n_2338),
.Y(n_2416)
);

AND2x4_ASAP7_75t_SL g2417 ( 
.A(n_2253),
.B(n_2187),
.Y(n_2417)
);

NAND2xp33_ASAP7_75t_L g2418 ( 
.A(n_2307),
.B(n_2213),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2258),
.B(n_2244),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2289),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_2251),
.B(n_2226),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2297),
.B(n_1302),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2315),
.B(n_1304),
.Y(n_2423)
);

BUFx3_ASAP7_75t_L g2424 ( 
.A(n_2315),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2255),
.B(n_1031),
.Y(n_2425)
);

NOR2xp67_ASAP7_75t_L g2426 ( 
.A(n_2268),
.B(n_788),
.Y(n_2426)
);

AOI21xp33_ASAP7_75t_L g2427 ( 
.A1(n_2259),
.A2(n_1038),
.B(n_1037),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2376),
.B(n_1316),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_2304),
.Y(n_2429)
);

BUFx12f_ASAP7_75t_L g2430 ( 
.A(n_2368),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2400),
.Y(n_2431)
);

INVxp33_ASAP7_75t_L g2432 ( 
.A(n_2261),
.Y(n_2432)
);

AOI22x1_ASAP7_75t_L g2433 ( 
.A1(n_2340),
.A2(n_1066),
.B1(n_1067),
.B2(n_1065),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2281),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2368),
.B(n_1329),
.Y(n_2435)
);

BUFx4f_ASAP7_75t_L g2436 ( 
.A(n_2253),
.Y(n_2436)
);

INVx5_ASAP7_75t_L g2437 ( 
.A(n_2396),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2342),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2396),
.B(n_1331),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2264),
.B(n_1043),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2403),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_2403),
.Y(n_2442)
);

INVx4_ASAP7_75t_L g2443 ( 
.A(n_2291),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2252),
.B(n_1052),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2254),
.Y(n_2445)
);

OAI21x1_ASAP7_75t_L g2446 ( 
.A1(n_2373),
.A2(n_1059),
.B(n_1054),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_2256),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2302),
.Y(n_2448)
);

AND3x1_ASAP7_75t_SL g2449 ( 
.A(n_2345),
.B(n_1061),
.C(n_1060),
.Y(n_2449)
);

CKINVDCx5p33_ASAP7_75t_R g2450 ( 
.A(n_2350),
.Y(n_2450)
);

BUFx12f_ASAP7_75t_L g2451 ( 
.A(n_2291),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2274),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2262),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2272),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2282),
.B(n_1068),
.Y(n_2455)
);

CKINVDCx16_ASAP7_75t_R g2456 ( 
.A(n_2383),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2286),
.B(n_1073),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2316),
.B(n_1069),
.Y(n_2458)
);

NAND2xp33_ASAP7_75t_L g2459 ( 
.A(n_2283),
.B(n_1078),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2393),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2300),
.B(n_1075),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2395),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2285),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2391),
.B(n_2306),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2271),
.B(n_1086),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2270),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2366),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2308),
.B(n_1317),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_SL g2469 ( 
.A(n_2317),
.B(n_1079),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2263),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2394),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2352),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2341),
.B(n_1319),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2397),
.Y(n_2474)
);

OAI22xp5_ASAP7_75t_SL g2475 ( 
.A1(n_2284),
.A2(n_1088),
.B1(n_1097),
.B2(n_1095),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2354),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2398),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2343),
.B(n_1100),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2348),
.B(n_2360),
.Y(n_2479)
);

CKINVDCx8_ASAP7_75t_R g2480 ( 
.A(n_2296),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2314),
.B(n_2319),
.Y(n_2481)
);

BUFx12f_ASAP7_75t_L g2482 ( 
.A(n_2321),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2386),
.Y(n_2483)
);

CKINVDCx16_ASAP7_75t_R g2484 ( 
.A(n_2322),
.Y(n_2484)
);

CKINVDCx20_ASAP7_75t_R g2485 ( 
.A(n_2294),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2290),
.Y(n_2486)
);

AOI22xp5_ASAP7_75t_L g2487 ( 
.A1(n_2364),
.A2(n_1091),
.B1(n_1094),
.B2(n_1092),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2293),
.B(n_1102),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2402),
.B(n_1103),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2399),
.B(n_1084),
.Y(n_2490)
);

CKINVDCx20_ASAP7_75t_R g2491 ( 
.A(n_2298),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2357),
.Y(n_2492)
);

BUFx2_ASAP7_75t_L g2493 ( 
.A(n_2260),
.Y(n_2493)
);

AND2x4_ASAP7_75t_L g2494 ( 
.A(n_2371),
.B(n_1104),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2312),
.B(n_1306),
.Y(n_2495)
);

OR2x6_ASAP7_75t_L g2496 ( 
.A(n_2299),
.B(n_1263),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2361),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2379),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2265),
.Y(n_2499)
);

BUFx12f_ASAP7_75t_L g2500 ( 
.A(n_2267),
.Y(n_2500)
);

AND2x4_ASAP7_75t_L g2501 ( 
.A(n_2358),
.B(n_1108),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_2374),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2347),
.Y(n_2503)
);

BUFx12f_ASAP7_75t_L g2504 ( 
.A(n_2288),
.Y(n_2504)
);

INVx6_ASAP7_75t_L g2505 ( 
.A(n_2266),
.Y(n_2505)
);

AO22x1_ASAP7_75t_L g2506 ( 
.A1(n_2401),
.A2(n_1287),
.B1(n_1311),
.B2(n_1281),
.Y(n_2506)
);

A2O1A1Ixp33_ASAP7_75t_L g2507 ( 
.A1(n_2355),
.A2(n_1311),
.B(n_1342),
.C(n_1341),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2278),
.B(n_1109),
.Y(n_2508)
);

INVx1_ASAP7_75t_SL g2509 ( 
.A(n_2320),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2324),
.B(n_1122),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2325),
.B(n_1269),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2380),
.Y(n_2512)
);

OAI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2362),
.A2(n_1124),
.B1(n_1127),
.B2(n_1123),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2381),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_R g2515 ( 
.A(n_2257),
.B(n_789),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_2387),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2353),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2323),
.Y(n_2518)
);

BUFx6f_ASAP7_75t_L g2519 ( 
.A(n_2336),
.Y(n_2519)
);

AOI22xp5_ASAP7_75t_L g2520 ( 
.A1(n_2385),
.A2(n_1099),
.B1(n_1105),
.B2(n_1096),
.Y(n_2520)
);

NAND2xp33_ASAP7_75t_L g2521 ( 
.A(n_2363),
.B(n_1098),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2328),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2329),
.Y(n_2523)
);

AOI22xp33_ASAP7_75t_L g2524 ( 
.A1(n_2370),
.A2(n_1131),
.B1(n_1133),
.B2(n_1130),
.Y(n_2524)
);

INVxp67_ASAP7_75t_L g2525 ( 
.A(n_2351),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2332),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2333),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2334),
.B(n_1310),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2335),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2356),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2337),
.B(n_1323),
.Y(n_2531)
);

CKINVDCx5p33_ASAP7_75t_R g2532 ( 
.A(n_2346),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2287),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2372),
.B(n_1136),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_2330),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2349),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2292),
.B(n_1147),
.Y(n_2537)
);

NAND2x1_ASAP7_75t_L g2538 ( 
.A(n_2377),
.B(n_1157),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2367),
.B(n_2359),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2279),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2311),
.A2(n_1152),
.B1(n_1154),
.B2(n_1151),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2326),
.B(n_1160),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2303),
.Y(n_2543)
);

INVx4_ASAP7_75t_L g2544 ( 
.A(n_2344),
.Y(n_2544)
);

BUFx3_ASAP7_75t_L g2545 ( 
.A(n_2313),
.Y(n_2545)
);

OAI21x1_ASAP7_75t_L g2546 ( 
.A1(n_2421),
.A2(n_2378),
.B(n_2384),
.Y(n_2546)
);

INVx4_ASAP7_75t_L g2547 ( 
.A(n_2447),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2405),
.Y(n_2548)
);

CKINVDCx20_ASAP7_75t_R g2549 ( 
.A(n_2456),
.Y(n_2549)
);

AOI22x1_ASAP7_75t_L g2550 ( 
.A1(n_2544),
.A2(n_1107),
.B1(n_1111),
.B2(n_1106),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2406),
.B(n_1166),
.Y(n_2551)
);

BUFx2_ASAP7_75t_L g2552 ( 
.A(n_2445),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2410),
.Y(n_2553)
);

AOI22xp5_ASAP7_75t_L g2554 ( 
.A1(n_2505),
.A2(n_2475),
.B1(n_2484),
.B2(n_2449),
.Y(n_2554)
);

BUFx8_ASAP7_75t_L g2555 ( 
.A(n_2500),
.Y(n_2555)
);

OAI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_2478),
.A2(n_2365),
.B(n_2389),
.Y(n_2556)
);

NAND2x1p5_ASAP7_75t_L g2557 ( 
.A(n_2437),
.B(n_2388),
.Y(n_2557)
);

BUFx12f_ASAP7_75t_L g2558 ( 
.A(n_2430),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2410),
.Y(n_2559)
);

INVx5_ASAP7_75t_L g2560 ( 
.A(n_2505),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2412),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_SL g2562 ( 
.A(n_2407),
.B(n_2273),
.Y(n_2562)
);

AND2x4_ASAP7_75t_L g2563 ( 
.A(n_2437),
.B(n_2375),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2415),
.Y(n_2564)
);

OR2x6_ASAP7_75t_L g2565 ( 
.A(n_2451),
.B(n_2339),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2445),
.Y(n_2566)
);

AOI22x1_ASAP7_75t_L g2567 ( 
.A1(n_2544),
.A2(n_1114),
.B1(n_1116),
.B2(n_1113),
.Y(n_2567)
);

INVxp67_ASAP7_75t_L g2568 ( 
.A(n_2411),
.Y(n_2568)
);

BUFx3_ASAP7_75t_L g2569 ( 
.A(n_2424),
.Y(n_2569)
);

CKINVDCx20_ASAP7_75t_R g2570 ( 
.A(n_2485),
.Y(n_2570)
);

OAI21x1_ASAP7_75t_L g2571 ( 
.A1(n_2446),
.A2(n_2438),
.B(n_2408),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2429),
.Y(n_2572)
);

BUFx3_ASAP7_75t_L g2573 ( 
.A(n_2450),
.Y(n_2573)
);

AND2x4_ASAP7_75t_L g2574 ( 
.A(n_2437),
.B(n_2390),
.Y(n_2574)
);

INVx3_ASAP7_75t_L g2575 ( 
.A(n_2454),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2452),
.Y(n_2576)
);

BUFx3_ASAP7_75t_L g2577 ( 
.A(n_2409),
.Y(n_2577)
);

BUFx5_ASAP7_75t_L g2578 ( 
.A(n_2499),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2453),
.Y(n_2579)
);

NOR2x1_ASAP7_75t_SL g2580 ( 
.A(n_2499),
.B(n_1292),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2431),
.Y(n_2581)
);

AO21x2_ASAP7_75t_L g2582 ( 
.A1(n_2460),
.A2(n_1179),
.B(n_1176),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2408),
.Y(n_2583)
);

OAI21x1_ASAP7_75t_SL g2584 ( 
.A1(n_2420),
.A2(n_1183),
.B(n_1180),
.Y(n_2584)
);

OAI21x1_ASAP7_75t_L g2585 ( 
.A1(n_2460),
.A2(n_1197),
.B(n_1188),
.Y(n_2585)
);

OR2x2_ASAP7_75t_L g2586 ( 
.A(n_2404),
.B(n_1199),
.Y(n_2586)
);

INVx1_ASAP7_75t_SL g2587 ( 
.A(n_2509),
.Y(n_2587)
);

BUFx3_ASAP7_75t_L g2588 ( 
.A(n_2519),
.Y(n_2588)
);

INVx4_ASAP7_75t_SL g2589 ( 
.A(n_2482),
.Y(n_2589)
);

BUFx8_ASAP7_75t_L g2590 ( 
.A(n_2504),
.Y(n_2590)
);

BUFx3_ASAP7_75t_L g2591 ( 
.A(n_2519),
.Y(n_2591)
);

AND2x4_ASAP7_75t_L g2592 ( 
.A(n_2443),
.B(n_1157),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2466),
.Y(n_2593)
);

CKINVDCx20_ASAP7_75t_R g2594 ( 
.A(n_2491),
.Y(n_2594)
);

INVx6_ASAP7_75t_SL g2595 ( 
.A(n_2496),
.Y(n_2595)
);

INVx5_ASAP7_75t_L g2596 ( 
.A(n_2516),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2466),
.Y(n_2597)
);

NOR2x1_ASAP7_75t_SL g2598 ( 
.A(n_2470),
.B(n_1285),
.Y(n_2598)
);

OA21x2_ASAP7_75t_L g2599 ( 
.A1(n_2434),
.A2(n_1203),
.B(n_1200),
.Y(n_2599)
);

HB1xp67_ASAP7_75t_L g2600 ( 
.A(n_2470),
.Y(n_2600)
);

AOI22x1_ASAP7_75t_L g2601 ( 
.A1(n_2516),
.A2(n_1209),
.B1(n_1223),
.B2(n_1208),
.Y(n_2601)
);

AND2x4_ASAP7_75t_L g2602 ( 
.A(n_2443),
.B(n_2441),
.Y(n_2602)
);

AND2x4_ASAP7_75t_L g2603 ( 
.A(n_2441),
.B(n_1285),
.Y(n_2603)
);

OAI21x1_ASAP7_75t_L g2604 ( 
.A1(n_2467),
.A2(n_1231),
.B(n_1230),
.Y(n_2604)
);

NAND2x1p5_ASAP7_75t_L g2605 ( 
.A(n_2436),
.B(n_1285),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2463),
.Y(n_2606)
);

INVx2_ASAP7_75t_SL g2607 ( 
.A(n_2417),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2454),
.Y(n_2608)
);

AOI21x1_ASAP7_75t_L g2609 ( 
.A1(n_2444),
.A2(n_2493),
.B(n_2419),
.Y(n_2609)
);

OAI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2427),
.A2(n_2275),
.B(n_1238),
.Y(n_2610)
);

OAI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2487),
.A2(n_1241),
.B(n_1236),
.Y(n_2611)
);

INVx4_ASAP7_75t_L g2612 ( 
.A(n_2486),
.Y(n_2612)
);

BUFx8_ASAP7_75t_L g2613 ( 
.A(n_2422),
.Y(n_2613)
);

AO21x2_ASAP7_75t_L g2614 ( 
.A1(n_2515),
.A2(n_1249),
.B(n_1244),
.Y(n_2614)
);

AO21x2_ASAP7_75t_L g2615 ( 
.A1(n_2414),
.A2(n_1266),
.B(n_1253),
.Y(n_2615)
);

INVx1_ASAP7_75t_SL g2616 ( 
.A(n_2502),
.Y(n_2616)
);

OAI21x1_ASAP7_75t_L g2617 ( 
.A1(n_2467),
.A2(n_1278),
.B(n_1274),
.Y(n_2617)
);

OAI21x1_ASAP7_75t_L g2618 ( 
.A1(n_2538),
.A2(n_1288),
.B(n_1279),
.Y(n_2618)
);

OAI21x1_ASAP7_75t_L g2619 ( 
.A1(n_2442),
.A2(n_1290),
.B(n_1289),
.Y(n_2619)
);

OAI21xp5_ASAP7_75t_L g2620 ( 
.A1(n_2520),
.A2(n_2459),
.B(n_2507),
.Y(n_2620)
);

HB1xp67_ASAP7_75t_L g2621 ( 
.A(n_2463),
.Y(n_2621)
);

AO21x2_ASAP7_75t_L g2622 ( 
.A1(n_2489),
.A2(n_1309),
.B(n_1118),
.Y(n_2622)
);

CKINVDCx20_ASAP7_75t_R g2623 ( 
.A(n_2448),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2540),
.Y(n_2624)
);

HB1xp67_ASAP7_75t_L g2625 ( 
.A(n_2540),
.Y(n_2625)
);

INVx2_ASAP7_75t_SL g2626 ( 
.A(n_2486),
.Y(n_2626)
);

OAI21x1_ASAP7_75t_L g2627 ( 
.A1(n_2442),
.A2(n_798),
.B(n_792),
.Y(n_2627)
);

INVx5_ASAP7_75t_L g2628 ( 
.A(n_2454),
.Y(n_2628)
);

BUFx2_ASAP7_75t_L g2629 ( 
.A(n_2465),
.Y(n_2629)
);

BUFx3_ASAP7_75t_L g2630 ( 
.A(n_2519),
.Y(n_2630)
);

AO21x2_ASAP7_75t_L g2631 ( 
.A1(n_2426),
.A2(n_1119),
.B(n_1117),
.Y(n_2631)
);

HB1xp67_ASAP7_75t_L g2632 ( 
.A(n_2536),
.Y(n_2632)
);

OAI21x1_ASAP7_75t_L g2633 ( 
.A1(n_2440),
.A2(n_802),
.B(n_800),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2464),
.B(n_2423),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2462),
.Y(n_2635)
);

AND2x4_ASAP7_75t_L g2636 ( 
.A(n_2465),
.B(n_1285),
.Y(n_2636)
);

AO21x2_ASAP7_75t_L g2637 ( 
.A1(n_2425),
.A2(n_1121),
.B(n_1120),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2486),
.B(n_1285),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2435),
.B(n_1125),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2536),
.Y(n_2640)
);

OAI21x1_ASAP7_75t_L g2641 ( 
.A1(n_2472),
.A2(n_804),
.B(n_803),
.Y(n_2641)
);

OR2x6_ASAP7_75t_L g2642 ( 
.A(n_2530),
.B(n_1292),
.Y(n_2642)
);

BUFx6f_ASAP7_75t_L g2643 ( 
.A(n_2436),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2471),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2474),
.Y(n_2645)
);

OAI21x1_ASAP7_75t_L g2646 ( 
.A1(n_2476),
.A2(n_809),
.B(n_808),
.Y(n_2646)
);

BUFx2_ASAP7_75t_SL g2647 ( 
.A(n_2545),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2503),
.Y(n_2648)
);

OR3x4_ASAP7_75t_SL g2649 ( 
.A(n_2413),
.B(n_1),
.C(n_3),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2522),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2624),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2564),
.Y(n_2652)
);

NAND2x1p5_ASAP7_75t_L g2653 ( 
.A(n_2560),
.B(n_2477),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2622),
.A2(n_2428),
.B1(n_2479),
.B2(n_2497),
.Y(n_2654)
);

OAI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2620),
.A2(n_2541),
.B1(n_2480),
.B2(n_2432),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2606),
.Y(n_2656)
);

INVx4_ASAP7_75t_SL g2657 ( 
.A(n_2558),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2615),
.A2(n_2498),
.B1(n_2514),
.B2(n_2481),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2640),
.Y(n_2659)
);

INVx6_ASAP7_75t_L g2660 ( 
.A(n_2560),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2621),
.B(n_2439),
.Y(n_2661)
);

AOI22xp33_ASAP7_75t_L g2662 ( 
.A1(n_2637),
.A2(n_2492),
.B1(n_2512),
.B2(n_2495),
.Y(n_2662)
);

CKINVDCx14_ASAP7_75t_R g2663 ( 
.A(n_2549),
.Y(n_2663)
);

BUFx2_ASAP7_75t_SL g2664 ( 
.A(n_2560),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2632),
.Y(n_2665)
);

INVxp67_ASAP7_75t_L g2666 ( 
.A(n_2647),
.Y(n_2666)
);

BUFx6f_ASAP7_75t_L g2667 ( 
.A(n_2569),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2625),
.Y(n_2668)
);

CKINVDCx11_ASAP7_75t_R g2669 ( 
.A(n_2570),
.Y(n_2669)
);

OAI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2554),
.A2(n_2517),
.B1(n_2535),
.B2(n_2532),
.Y(n_2670)
);

BUFx8_ASAP7_75t_SL g2671 ( 
.A(n_2623),
.Y(n_2671)
);

BUFx3_ASAP7_75t_L g2672 ( 
.A(n_2573),
.Y(n_2672)
);

AOI22xp33_ASAP7_75t_L g2673 ( 
.A1(n_2614),
.A2(n_2468),
.B1(n_2483),
.B2(n_2526),
.Y(n_2673)
);

OAI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2601),
.A2(n_2523),
.B1(n_2518),
.B2(n_2496),
.Y(n_2674)
);

BUFx4f_ASAP7_75t_SL g2675 ( 
.A(n_2594),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2577),
.Y(n_2676)
);

OAI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2629),
.A2(n_2525),
.B1(n_2539),
.B2(n_2542),
.Y(n_2677)
);

AOI22xp33_ASAP7_75t_L g2678 ( 
.A1(n_2644),
.A2(n_2527),
.B1(n_2529),
.B2(n_2473),
.Y(n_2678)
);

INVx6_ASAP7_75t_L g2679 ( 
.A(n_2555),
.Y(n_2679)
);

OAI22xp33_ASAP7_75t_L g2680 ( 
.A1(n_2629),
.A2(n_2533),
.B1(n_2543),
.B2(n_2461),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2579),
.Y(n_2681)
);

BUFx8_ASAP7_75t_SL g2682 ( 
.A(n_2572),
.Y(n_2682)
);

INVxp67_ASAP7_75t_SL g2683 ( 
.A(n_2600),
.Y(n_2683)
);

BUFx10_ASAP7_75t_L g2684 ( 
.A(n_2592),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2576),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2583),
.Y(n_2686)
);

INVx5_ASAP7_75t_L g2687 ( 
.A(n_2643),
.Y(n_2687)
);

INVx2_ASAP7_75t_SL g2688 ( 
.A(n_2588),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2593),
.Y(n_2689)
);

CKINVDCx11_ASAP7_75t_R g2690 ( 
.A(n_2589),
.Y(n_2690)
);

INVx4_ASAP7_75t_L g2691 ( 
.A(n_2547),
.Y(n_2691)
);

BUFx12f_ASAP7_75t_L g2692 ( 
.A(n_2555),
.Y(n_2692)
);

BUFx4f_ASAP7_75t_L g2693 ( 
.A(n_2643),
.Y(n_2693)
);

BUFx4f_ASAP7_75t_SL g2694 ( 
.A(n_2590),
.Y(n_2694)
);

BUFx3_ASAP7_75t_L g2695 ( 
.A(n_2590),
.Y(n_2695)
);

INVx3_ASAP7_75t_L g2696 ( 
.A(n_2612),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2591),
.Y(n_2697)
);

INVx5_ASAP7_75t_L g2698 ( 
.A(n_2643),
.Y(n_2698)
);

INVx1_ASAP7_75t_SL g2699 ( 
.A(n_2647),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2597),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2645),
.A2(n_2501),
.B1(n_2494),
.B2(n_2510),
.Y(n_2701)
);

AOI22xp5_ASAP7_75t_L g2702 ( 
.A1(n_2568),
.A2(n_2418),
.B1(n_2636),
.B2(n_2562),
.Y(n_2702)
);

OAI22xp33_ASAP7_75t_L g2703 ( 
.A1(n_2601),
.A2(n_2455),
.B1(n_2457),
.B2(n_2534),
.Y(n_2703)
);

BUFx6f_ASAP7_75t_L g2704 ( 
.A(n_2630),
.Y(n_2704)
);

CKINVDCx20_ASAP7_75t_R g2705 ( 
.A(n_2613),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2551),
.A2(n_2501),
.B1(n_2494),
.B2(n_2511),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2612),
.Y(n_2707)
);

BUFx12f_ASAP7_75t_L g2708 ( 
.A(n_2613),
.Y(n_2708)
);

OAI22xp5_ASAP7_75t_L g2709 ( 
.A1(n_2556),
.A2(n_2524),
.B1(n_2458),
.B2(n_2469),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2648),
.B(n_2416),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_2582),
.A2(n_2528),
.B1(n_2508),
.B2(n_2531),
.Y(n_2711)
);

INVx11_ASAP7_75t_L g2712 ( 
.A(n_2589),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2634),
.B(n_2508),
.Y(n_2713)
);

BUFx6f_ASAP7_75t_L g2714 ( 
.A(n_2607),
.Y(n_2714)
);

OAI21xp5_ASAP7_75t_SL g2715 ( 
.A1(n_2649),
.A2(n_2490),
.B(n_2513),
.Y(n_2715)
);

INVx3_ASAP7_75t_L g2716 ( 
.A(n_2547),
.Y(n_2716)
);

OAI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2596),
.A2(n_2433),
.B1(n_2537),
.B2(n_2488),
.Y(n_2717)
);

INVx6_ASAP7_75t_L g2718 ( 
.A(n_2596),
.Y(n_2718)
);

INVx6_ASAP7_75t_L g2719 ( 
.A(n_2596),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2553),
.Y(n_2720)
);

INVx8_ASAP7_75t_L g2721 ( 
.A(n_2565),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2616),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2559),
.Y(n_2723)
);

CKINVDCx11_ASAP7_75t_R g2724 ( 
.A(n_2587),
.Y(n_2724)
);

NAND2x1p5_ASAP7_75t_L g2725 ( 
.A(n_2628),
.B(n_2506),
.Y(n_2725)
);

CKINVDCx20_ASAP7_75t_R g2726 ( 
.A(n_2626),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2561),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2548),
.Y(n_2728)
);

AOI22xp33_ASAP7_75t_SL g2729 ( 
.A1(n_2599),
.A2(n_2598),
.B1(n_2584),
.B2(n_2580),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2650),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2683),
.B(n_2552),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2669),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2665),
.B(n_2668),
.Y(n_2733)
);

AND2x2_ASAP7_75t_SL g2734 ( 
.A(n_2710),
.B(n_2552),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2661),
.B(n_2566),
.Y(n_2735)
);

A2O1A1Ixp33_ASAP7_75t_L g2736 ( 
.A1(n_2715),
.A2(n_2521),
.B(n_2611),
.C(n_2610),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2703),
.A2(n_2580),
.B(n_2598),
.Y(n_2737)
);

AND2x4_ASAP7_75t_L g2738 ( 
.A(n_2699),
.B(n_2566),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2730),
.Y(n_2739)
);

A2O1A1Ixp33_ASAP7_75t_L g2740 ( 
.A1(n_2655),
.A2(n_2563),
.B(n_2574),
.C(n_2636),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2727),
.B(n_2578),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_L g2742 ( 
.A1(n_2654),
.A2(n_2658),
.B1(n_2662),
.B2(n_2673),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2690),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2651),
.B(n_2578),
.Y(n_2744)
);

OAI21x1_ASAP7_75t_L g2745 ( 
.A1(n_2653),
.A2(n_2609),
.B(n_2571),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2656),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2659),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2686),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2652),
.Y(n_2749)
);

OR2x2_ASAP7_75t_L g2750 ( 
.A(n_2689),
.B(n_2586),
.Y(n_2750)
);

OA21x2_ASAP7_75t_L g2751 ( 
.A1(n_2666),
.A2(n_2609),
.B(n_2581),
.Y(n_2751)
);

OAI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2702),
.A2(n_2602),
.B1(n_2557),
.B2(n_2642),
.Y(n_2752)
);

AOI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2677),
.A2(n_2584),
.B(n_2599),
.Y(n_2753)
);

INVx1_ASAP7_75t_SL g2754 ( 
.A(n_2675),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2663),
.B(n_2602),
.Y(n_2755)
);

OR2x2_ASAP7_75t_L g2756 ( 
.A(n_2700),
.B(n_2635),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2720),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2724),
.B(n_2672),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2723),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2688),
.B(n_2578),
.Y(n_2760)
);

HB1xp67_ASAP7_75t_L g2761 ( 
.A(n_2697),
.Y(n_2761)
);

OAI21x1_ASAP7_75t_L g2762 ( 
.A1(n_2725),
.A2(n_2617),
.B(n_2604),
.Y(n_2762)
);

NAND2x1p5_ASAP7_75t_L g2763 ( 
.A(n_2687),
.B(n_2628),
.Y(n_2763)
);

OA21x2_ASAP7_75t_L g2764 ( 
.A1(n_2678),
.A2(n_2585),
.B(n_2646),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2681),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2717),
.A2(n_2642),
.B(n_2574),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2713),
.B(n_2578),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2696),
.B(n_2575),
.Y(n_2768)
);

AOI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2711),
.A2(n_2595),
.B1(n_2631),
.B2(n_2639),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2701),
.A2(n_2595),
.B1(n_2563),
.B2(n_2575),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2685),
.Y(n_2771)
);

A2O1A1Ixp33_ASAP7_75t_L g2772 ( 
.A1(n_2709),
.A2(n_2546),
.B(n_2641),
.C(n_2633),
.Y(n_2772)
);

OAI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2674),
.A2(n_2592),
.B(n_2567),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2728),
.Y(n_2774)
);

INVx4_ASAP7_75t_L g2775 ( 
.A(n_2712),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2718),
.Y(n_2776)
);

O2A1O1Ixp33_ASAP7_75t_L g2777 ( 
.A1(n_2680),
.A2(n_2565),
.B(n_2638),
.C(n_2603),
.Y(n_2777)
);

A2O1A1Ixp33_ASAP7_75t_L g2778 ( 
.A1(n_2706),
.A2(n_2638),
.B(n_2627),
.C(n_2608),
.Y(n_2778)
);

OAI22xp33_ASAP7_75t_L g2779 ( 
.A1(n_2721),
.A2(n_2628),
.B1(n_2608),
.B2(n_2605),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2707),
.Y(n_2780)
);

BUFx3_ASAP7_75t_L g2781 ( 
.A(n_2692),
.Y(n_2781)
);

A2O1A1Ixp33_ASAP7_75t_L g2782 ( 
.A1(n_2729),
.A2(n_2603),
.B(n_2619),
.C(n_2618),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2716),
.B(n_1292),
.Y(n_2783)
);

AOI21x1_ASAP7_75t_L g2784 ( 
.A1(n_2670),
.A2(n_2550),
.B(n_1357),
.Y(n_2784)
);

AO21x2_ASAP7_75t_L g2785 ( 
.A1(n_2718),
.A2(n_1357),
.B(n_1292),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2704),
.B(n_1292),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2691),
.B(n_1357),
.Y(n_2787)
);

INVx4_ASAP7_75t_L g2788 ( 
.A(n_2679),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2704),
.Y(n_2789)
);

BUFx2_ASAP7_75t_L g2790 ( 
.A(n_2726),
.Y(n_2790)
);

HB1xp67_ASAP7_75t_L g2791 ( 
.A(n_2719),
.Y(n_2791)
);

OAI21x1_ASAP7_75t_L g2792 ( 
.A1(n_2664),
.A2(n_4),
.B(n_5),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2684),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2676),
.B(n_1357),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2719),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2664),
.B(n_1357),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2684),
.Y(n_2797)
);

AOI322xp5_ASAP7_75t_L g2798 ( 
.A1(n_2721),
.A2(n_1137),
.A3(n_1128),
.B1(n_1138),
.B2(n_1140),
.C1(n_1135),
.C2(n_1126),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2667),
.B(n_6),
.Y(n_2799)
);

AOI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2693),
.A2(n_1143),
.B(n_1142),
.Y(n_2800)
);

OAI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2660),
.A2(n_2705),
.B1(n_2679),
.B2(n_2714),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2660),
.Y(n_2802)
);

INVx3_ASAP7_75t_L g2803 ( 
.A(n_2667),
.Y(n_2803)
);

OAI21x1_ASAP7_75t_L g2804 ( 
.A1(n_2687),
.A2(n_6),
.B(n_7),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2738),
.B(n_2657),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_2742),
.A2(n_2708),
.B1(n_2695),
.B2(n_2714),
.Y(n_2806)
);

AOI22xp33_ASAP7_75t_L g2807 ( 
.A1(n_2753),
.A2(n_2694),
.B1(n_2657),
.B2(n_2722),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2765),
.Y(n_2808)
);

HB1xp67_ASAP7_75t_L g2809 ( 
.A(n_2731),
.Y(n_2809)
);

NAND3xp33_ASAP7_75t_L g2810 ( 
.A(n_2741),
.B(n_2698),
.C(n_2687),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2738),
.B(n_2791),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2769),
.A2(n_1145),
.B1(n_1149),
.B2(n_1144),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2734),
.B(n_2698),
.Y(n_2813)
);

INVx3_ASAP7_75t_L g2814 ( 
.A(n_2776),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_SL g2815 ( 
.A1(n_2764),
.A2(n_2698),
.B1(n_1193),
.B2(n_1214),
.Y(n_2815)
);

OAI22xp33_ASAP7_75t_L g2816 ( 
.A1(n_2737),
.A2(n_1158),
.B1(n_1159),
.B2(n_1155),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2751),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_L g2818 ( 
.A1(n_2764),
.A2(n_1163),
.B1(n_1165),
.B2(n_1162),
.Y(n_2818)
);

OAI22xp33_ASAP7_75t_L g2819 ( 
.A1(n_2752),
.A2(n_1168),
.B1(n_1170),
.B2(n_1167),
.Y(n_2819)
);

A2O1A1Ixp33_ASAP7_75t_L g2820 ( 
.A1(n_2736),
.A2(n_1174),
.B(n_1175),
.C(n_1171),
.Y(n_2820)
);

HB1xp67_ASAP7_75t_L g2821 ( 
.A(n_2735),
.Y(n_2821)
);

AOI221xp5_ASAP7_75t_L g2822 ( 
.A1(n_2772),
.A2(n_1187),
.B1(n_1195),
.B2(n_1181),
.C(n_1177),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2765),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2747),
.Y(n_2824)
);

OAI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2740),
.A2(n_1201),
.B1(n_1202),
.B2(n_1198),
.Y(n_2825)
);

AOI22xp33_ASAP7_75t_L g2826 ( 
.A1(n_2773),
.A2(n_1205),
.B1(n_1212),
.B2(n_1204),
.Y(n_2826)
);

INVxp67_ASAP7_75t_L g2827 ( 
.A(n_2761),
.Y(n_2827)
);

AOI22xp33_ASAP7_75t_L g2828 ( 
.A1(n_2750),
.A2(n_1218),
.B1(n_1219),
.B2(n_1215),
.Y(n_2828)
);

BUFx12f_ASAP7_75t_L g2829 ( 
.A(n_2732),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2794),
.B(n_2671),
.Y(n_2830)
);

AOI22xp33_ASAP7_75t_L g2831 ( 
.A1(n_2770),
.A2(n_1221),
.B1(n_1225),
.B2(n_1220),
.Y(n_2831)
);

AND2x4_ASAP7_75t_SL g2832 ( 
.A(n_2788),
.B(n_2682),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2751),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2747),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2755),
.B(n_8),
.Y(n_2835)
);

AOI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_2799),
.A2(n_1232),
.B1(n_1233),
.B2(n_1227),
.Y(n_2836)
);

OAI22xp5_ASAP7_75t_SL g2837 ( 
.A1(n_2743),
.A2(n_2788),
.B1(n_2775),
.B2(n_2801),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2749),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2756),
.Y(n_2839)
);

AOI22xp33_ASAP7_75t_SL g2840 ( 
.A1(n_2766),
.A2(n_1255),
.B1(n_1268),
.B2(n_1234),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2795),
.B(n_9),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_2743),
.A2(n_1242),
.B1(n_1243),
.B2(n_1240),
.Y(n_2842)
);

OR2x6_ASAP7_75t_L g2843 ( 
.A(n_2777),
.B(n_10),
.Y(n_2843)
);

OR2x2_ASAP7_75t_L g2844 ( 
.A(n_2733),
.B(n_10),
.Y(n_2844)
);

OA21x2_ASAP7_75t_L g2845 ( 
.A1(n_2745),
.A2(n_1247),
.B(n_1245),
.Y(n_2845)
);

AOI22xp33_ASAP7_75t_L g2846 ( 
.A1(n_2743),
.A2(n_1254),
.B1(n_1256),
.B2(n_1251),
.Y(n_2846)
);

CKINVDCx5p33_ASAP7_75t_R g2847 ( 
.A(n_2754),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2746),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2814),
.B(n_2776),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2824),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2813),
.Y(n_2851)
);

INVx4_ASAP7_75t_L g2852 ( 
.A(n_2829),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2814),
.B(n_2793),
.Y(n_2853)
);

BUFx2_ASAP7_75t_L g2854 ( 
.A(n_2805),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2817),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2817),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2833),
.Y(n_2857)
);

BUFx3_ASAP7_75t_L g2858 ( 
.A(n_2832),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2811),
.B(n_2797),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2833),
.Y(n_2860)
);

HB1xp67_ASAP7_75t_L g2861 ( 
.A(n_2821),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2834),
.Y(n_2862)
);

BUFx2_ASAP7_75t_L g2863 ( 
.A(n_2809),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2839),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2839),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2848),
.Y(n_2866)
);

HB1xp67_ASAP7_75t_L g2867 ( 
.A(n_2827),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2844),
.B(n_2748),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2808),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2823),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2818),
.B(n_2757),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2845),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2818),
.B(n_2759),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2832),
.B(n_2775),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2847),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2807),
.B(n_2802),
.Y(n_2876)
);

NOR2x1_ASAP7_75t_L g2877 ( 
.A(n_2830),
.B(n_2758),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2845),
.Y(n_2878)
);

OAI221xp5_ASAP7_75t_L g2879 ( 
.A1(n_2826),
.A2(n_2778),
.B1(n_2782),
.B2(n_2786),
.C(n_2798),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2807),
.B(n_2768),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2838),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2835),
.B(n_2768),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2806),
.B(n_2739),
.Y(n_2883)
);

OR2x6_ASAP7_75t_L g2884 ( 
.A(n_2843),
.B(n_2763),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2845),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2854),
.B(n_2830),
.Y(n_2886)
);

OA21x2_ASAP7_75t_L g2887 ( 
.A1(n_2855),
.A2(n_2806),
.B(n_2822),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2872),
.B(n_2828),
.Y(n_2888)
);

AOI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2884),
.A2(n_2837),
.B(n_2871),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2866),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2884),
.A2(n_2879),
.B(n_2878),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2859),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2850),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2850),
.Y(n_2894)
);

AO31x2_ASAP7_75t_L g2895 ( 
.A1(n_2878),
.A2(n_2825),
.A3(n_2820),
.B(n_2789),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2862),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2859),
.Y(n_2897)
);

AND2x2_ASAP7_75t_L g2898 ( 
.A(n_2854),
.B(n_2851),
.Y(n_2898)
);

AO21x2_ASAP7_75t_L g2899 ( 
.A1(n_2885),
.A2(n_2796),
.B(n_2816),
.Y(n_2899)
);

OA21x2_ASAP7_75t_L g2900 ( 
.A1(n_2855),
.A2(n_2810),
.B(n_2790),
.Y(n_2900)
);

INVx4_ASAP7_75t_L g2901 ( 
.A(n_2852),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2861),
.Y(n_2902)
);

INVx4_ASAP7_75t_L g2903 ( 
.A(n_2852),
.Y(n_2903)
);

OAI21x1_ASAP7_75t_L g2904 ( 
.A1(n_2856),
.A2(n_2760),
.B(n_2744),
.Y(n_2904)
);

OAI211xp5_ASAP7_75t_SL g2905 ( 
.A1(n_2877),
.A2(n_2846),
.B(n_2842),
.C(n_2826),
.Y(n_2905)
);

OAI221xp5_ASAP7_75t_L g2906 ( 
.A1(n_2873),
.A2(n_2815),
.B1(n_2812),
.B2(n_2836),
.C(n_2842),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2867),
.Y(n_2907)
);

INVx4_ASAP7_75t_SL g2908 ( 
.A(n_2858),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_L g2909 ( 
.A(n_2852),
.B(n_2781),
.Y(n_2909)
);

OAI211xp5_ASAP7_75t_L g2910 ( 
.A1(n_2863),
.A2(n_2846),
.B(n_2836),
.C(n_2840),
.Y(n_2910)
);

OAI221xp5_ASAP7_75t_L g2911 ( 
.A1(n_2885),
.A2(n_2812),
.B1(n_2828),
.B2(n_2843),
.C(n_2831),
.Y(n_2911)
);

AOI22xp5_ASAP7_75t_L g2912 ( 
.A1(n_2884),
.A2(n_2843),
.B1(n_2819),
.B2(n_2831),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2868),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2856),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2864),
.Y(n_2915)
);

OAI21xp33_ASAP7_75t_L g2916 ( 
.A1(n_2883),
.A2(n_2787),
.B(n_2783),
.Y(n_2916)
);

INVx4_ASAP7_75t_L g2917 ( 
.A(n_2875),
.Y(n_2917)
);

AOI21x1_ASAP7_75t_L g2918 ( 
.A1(n_2884),
.A2(n_2876),
.B(n_2851),
.Y(n_2918)
);

AND2x2_ASAP7_75t_L g2919 ( 
.A(n_2880),
.B(n_2803),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2857),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2865),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2869),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2869),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2857),
.Y(n_2924)
);

OR2x2_ASAP7_75t_L g2925 ( 
.A(n_2913),
.B(n_2907),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2896),
.Y(n_2926)
);

AND2x4_ASAP7_75t_SL g2927 ( 
.A(n_2886),
.B(n_2882),
.Y(n_2927)
);

OAI221xp5_ASAP7_75t_L g2928 ( 
.A1(n_2891),
.A2(n_2888),
.B1(n_2911),
.B2(n_2912),
.C(n_2887),
.Y(n_2928)
);

AOI211xp5_ASAP7_75t_SL g2929 ( 
.A1(n_2910),
.A2(n_2874),
.B(n_2880),
.C(n_2876),
.Y(n_2929)
);

NAND3xp33_ASAP7_75t_L g2930 ( 
.A(n_2888),
.B(n_2860),
.C(n_2863),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2898),
.B(n_2858),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2908),
.B(n_2849),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2899),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2899),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2890),
.Y(n_2935)
);

INVx6_ASAP7_75t_L g2936 ( 
.A(n_2908),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2892),
.Y(n_2937)
);

INVx1_ASAP7_75t_SL g2938 ( 
.A(n_2917),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2893),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2894),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2902),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2919),
.B(n_2849),
.Y(n_2942)
);

AND2x2_ASAP7_75t_L g2943 ( 
.A(n_2897),
.B(n_2853),
.Y(n_2943)
);

AND4x1_ASAP7_75t_L g2944 ( 
.A(n_2912),
.B(n_2841),
.C(n_2882),
.D(n_2800),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2900),
.B(n_2853),
.Y(n_2945)
);

INVx2_ASAP7_75t_SL g2946 ( 
.A(n_2917),
.Y(n_2946)
);

INVx2_ASAP7_75t_SL g2947 ( 
.A(n_2901),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2900),
.B(n_2875),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2918),
.B(n_2780),
.Y(n_2949)
);

INVxp67_ASAP7_75t_L g2950 ( 
.A(n_2909),
.Y(n_2950)
);

BUFx3_ASAP7_75t_L g2951 ( 
.A(n_2901),
.Y(n_2951)
);

OR2x2_ASAP7_75t_L g2952 ( 
.A(n_2915),
.B(n_2860),
.Y(n_2952)
);

BUFx3_ASAP7_75t_L g2953 ( 
.A(n_2903),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2903),
.B(n_2803),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2922),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2895),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2889),
.B(n_2870),
.Y(n_2957)
);

BUFx2_ASAP7_75t_L g2958 ( 
.A(n_2895),
.Y(n_2958)
);

NOR3xp33_ASAP7_75t_L g2959 ( 
.A(n_2911),
.B(n_2784),
.C(n_2792),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2923),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2939),
.Y(n_2961)
);

INVx2_ASAP7_75t_SL g2962 ( 
.A(n_2936),
.Y(n_2962)
);

INVx2_ASAP7_75t_SL g2963 ( 
.A(n_2936),
.Y(n_2963)
);

OAI33xp33_ASAP7_75t_L g2964 ( 
.A1(n_2930),
.A2(n_2905),
.A3(n_2921),
.B1(n_2916),
.B2(n_1260),
.B3(n_1258),
.Y(n_2964)
);

NOR2xp33_ASAP7_75t_L g2965 ( 
.A(n_2936),
.B(n_2906),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2927),
.B(n_2887),
.Y(n_2966)
);

AND2x2_ASAP7_75t_L g2967 ( 
.A(n_2927),
.B(n_2895),
.Y(n_2967)
);

OAI21xp33_ASAP7_75t_L g2968 ( 
.A1(n_2948),
.A2(n_2891),
.B(n_2916),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2958),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2931),
.B(n_2904),
.Y(n_2970)
);

OR2x2_ASAP7_75t_L g2971 ( 
.A(n_2925),
.B(n_2914),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2940),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2931),
.B(n_2920),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2933),
.Y(n_2974)
);

NAND5xp2_ASAP7_75t_L g2975 ( 
.A(n_2948),
.B(n_2906),
.C(n_2767),
.D(n_2804),
.E(n_2779),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2932),
.B(n_2924),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2941),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2929),
.B(n_2870),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2932),
.B(n_2881),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2955),
.Y(n_2980)
);

OR2x2_ASAP7_75t_L g2981 ( 
.A(n_2937),
.B(n_2926),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2960),
.Y(n_2982)
);

AND2x4_ASAP7_75t_L g2983 ( 
.A(n_2946),
.B(n_2881),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2935),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2937),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2952),
.Y(n_2986)
);

NOR2xp67_ASAP7_75t_L g2987 ( 
.A(n_2950),
.B(n_11),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2954),
.B(n_2774),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2954),
.B(n_2785),
.Y(n_2989)
);

INVx4_ASAP7_75t_L g2990 ( 
.A(n_2951),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2938),
.B(n_2785),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2943),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2943),
.Y(n_2993)
);

AND2x2_ASAP7_75t_L g2994 ( 
.A(n_2942),
.B(n_2946),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2959),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2951),
.B(n_11),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2944),
.B(n_1257),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2933),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2934),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2934),
.Y(n_3000)
);

INVx1_ASAP7_75t_SL g3001 ( 
.A(n_2953),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2945),
.B(n_2762),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2947),
.Y(n_3003)
);

INVx1_ASAP7_75t_SL g3004 ( 
.A(n_2953),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2945),
.B(n_12),
.Y(n_3005)
);

AND2x4_ASAP7_75t_L g3006 ( 
.A(n_2947),
.B(n_2771),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2956),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_3005),
.B(n_2957),
.Y(n_3008)
);

INVx2_ASAP7_75t_SL g3009 ( 
.A(n_2973),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2973),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2962),
.Y(n_3011)
);

NOR3xp33_ASAP7_75t_L g3012 ( 
.A(n_2968),
.B(n_2928),
.C(n_2957),
.Y(n_3012)
);

OR2x2_ASAP7_75t_L g3013 ( 
.A(n_2992),
.B(n_2949),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2962),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2969),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2969),
.Y(n_3016)
);

XOR2x2_ASAP7_75t_L g3017 ( 
.A(n_2987),
.B(n_2949),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2963),
.Y(n_3018)
);

INVx3_ASAP7_75t_L g3019 ( 
.A(n_2990),
.Y(n_3019)
);

BUFx2_ASAP7_75t_L g3020 ( 
.A(n_2963),
.Y(n_3020)
);

BUFx2_ASAP7_75t_L g3021 ( 
.A(n_3005),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2993),
.B(n_2986),
.Y(n_3022)
);

XOR2x2_ASAP7_75t_L g3023 ( 
.A(n_2965),
.B(n_2956),
.Y(n_3023)
);

INVx2_ASAP7_75t_SL g3024 ( 
.A(n_2994),
.Y(n_3024)
);

AND2x4_ASAP7_75t_L g3025 ( 
.A(n_2990),
.B(n_12),
.Y(n_3025)
);

NAND4xp75_ASAP7_75t_L g3026 ( 
.A(n_2965),
.B(n_1261),
.C(n_1267),
.D(n_1259),
.Y(n_3026)
);

AND2x2_ASAP7_75t_SL g3027 ( 
.A(n_2966),
.B(n_13),
.Y(n_3027)
);

INVx1_ASAP7_75t_SL g3028 ( 
.A(n_2967),
.Y(n_3028)
);

NAND4xp75_ASAP7_75t_L g3029 ( 
.A(n_2995),
.B(n_2978),
.C(n_2997),
.D(n_2998),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2977),
.Y(n_3030)
);

XOR2x2_ASAP7_75t_L g3031 ( 
.A(n_2975),
.B(n_14),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2977),
.Y(n_3032)
);

NAND4xp75_ASAP7_75t_L g3033 ( 
.A(n_2999),
.B(n_3000),
.C(n_2974),
.D(n_2985),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2981),
.Y(n_3034)
);

INVxp67_ASAP7_75t_SL g3035 ( 
.A(n_2996),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_3003),
.B(n_1275),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2971),
.Y(n_3037)
);

AND2x4_ASAP7_75t_L g3038 ( 
.A(n_2990),
.B(n_15),
.Y(n_3038)
);

INVx6_ASAP7_75t_L g3039 ( 
.A(n_2976),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2984),
.Y(n_3040)
);

NAND4xp75_ASAP7_75t_L g3041 ( 
.A(n_2970),
.B(n_17),
.C(n_15),
.D(n_16),
.Y(n_3041)
);

AOI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2964),
.A2(n_1276),
.B1(n_18),
.B2(n_16),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2979),
.Y(n_3043)
);

XOR2x2_ASAP7_75t_L g3044 ( 
.A(n_2964),
.B(n_17),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2961),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2972),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2980),
.Y(n_3047)
);

INVx1_ASAP7_75t_SL g3048 ( 
.A(n_3001),
.Y(n_3048)
);

NOR2xp33_ASAP7_75t_L g3049 ( 
.A(n_3004),
.B(n_19),
.Y(n_3049)
);

OR2x2_ASAP7_75t_L g3050 ( 
.A(n_2982),
.B(n_20),
.Y(n_3050)
);

AND2x2_ASAP7_75t_L g3051 ( 
.A(n_2983),
.B(n_21),
.Y(n_3051)
);

NOR3xp33_ASAP7_75t_L g3052 ( 
.A(n_2991),
.B(n_22),
.C(n_24),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2983),
.B(n_25),
.Y(n_3053)
);

OR2x2_ASAP7_75t_L g3054 ( 
.A(n_2983),
.B(n_25),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2989),
.Y(n_3055)
);

XNOR2xp5_ASAP7_75t_L g3056 ( 
.A(n_3006),
.B(n_26),
.Y(n_3056)
);

INVxp67_ASAP7_75t_L g3057 ( 
.A(n_3006),
.Y(n_3057)
);

INVx1_ASAP7_75t_SL g3058 ( 
.A(n_3006),
.Y(n_3058)
);

NAND4xp75_ASAP7_75t_L g3059 ( 
.A(n_2974),
.B(n_28),
.C(n_26),
.D(n_27),
.Y(n_3059)
);

XOR2x2_ASAP7_75t_L g3060 ( 
.A(n_3002),
.B(n_29),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_3007),
.Y(n_3061)
);

NAND4xp75_ASAP7_75t_L g3062 ( 
.A(n_3000),
.B(n_33),
.C(n_29),
.D(n_30),
.Y(n_3062)
);

NAND4xp75_ASAP7_75t_SL g3063 ( 
.A(n_3002),
.B(n_34),
.C(n_30),
.D(n_33),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_3007),
.Y(n_3064)
);

XNOR2xp5_ASAP7_75t_L g3065 ( 
.A(n_2988),
.B(n_34),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2969),
.Y(n_3066)
);

INVx1_ASAP7_75t_SL g3067 ( 
.A(n_2966),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2973),
.Y(n_3068)
);

NAND4xp75_ASAP7_75t_SL g3069 ( 
.A(n_3005),
.B(n_39),
.C(n_37),
.D(n_38),
.Y(n_3069)
);

INVxp67_ASAP7_75t_L g3070 ( 
.A(n_2965),
.Y(n_3070)
);

INVx4_ASAP7_75t_L g3071 ( 
.A(n_2990),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_3005),
.B(n_37),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2973),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2969),
.Y(n_3074)
);

XOR2x2_ASAP7_75t_L g3075 ( 
.A(n_2987),
.B(n_39),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3033),
.Y(n_3076)
);

AND2x2_ASAP7_75t_L g3077 ( 
.A(n_3067),
.B(n_40),
.Y(n_3077)
);

NAND2x1p5_ASAP7_75t_L g3078 ( 
.A(n_3048),
.B(n_3051),
.Y(n_3078)
);

NAND4xp25_ASAP7_75t_L g3079 ( 
.A(n_3012),
.B(n_42),
.C(n_40),
.D(n_41),
.Y(n_3079)
);

INVx2_ASAP7_75t_SL g3080 ( 
.A(n_3039),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_3021),
.Y(n_3081)
);

HB1xp67_ASAP7_75t_L g3082 ( 
.A(n_3020),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_3009),
.B(n_41),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_3024),
.B(n_42),
.Y(n_3084)
);

OR2x2_ASAP7_75t_L g3085 ( 
.A(n_3010),
.B(n_43),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3072),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_3030),
.Y(n_3087)
);

OR2x2_ASAP7_75t_L g3088 ( 
.A(n_3068),
.B(n_3073),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_3032),
.Y(n_3089)
);

INVx2_ASAP7_75t_SL g3090 ( 
.A(n_3039),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3015),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_3016),
.Y(n_3092)
);

INVxp67_ASAP7_75t_L g3093 ( 
.A(n_3026),
.Y(n_3093)
);

NAND2xp33_ASAP7_75t_L g3094 ( 
.A(n_3008),
.B(n_43),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_3011),
.B(n_44),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_3075),
.Y(n_3096)
);

OR2x2_ASAP7_75t_L g3097 ( 
.A(n_3034),
.B(n_45),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_3066),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_3074),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_3054),
.Y(n_3100)
);

INVxp67_ASAP7_75t_L g3101 ( 
.A(n_3026),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_3014),
.B(n_45),
.Y(n_3102)
);

A2O1A1Ixp33_ASAP7_75t_L g3103 ( 
.A1(n_3042),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_3061),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_3018),
.B(n_48),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_3049),
.B(n_49),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_3025),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_3064),
.Y(n_3108)
);

OR2x2_ASAP7_75t_L g3109 ( 
.A(n_3013),
.B(n_50),
.Y(n_3109)
);

NOR2xp67_ASAP7_75t_L g3110 ( 
.A(n_3057),
.B(n_50),
.Y(n_3110)
);

OR2x2_ASAP7_75t_L g3111 ( 
.A(n_3035),
.B(n_51),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_3025),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3050),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_3027),
.B(n_53),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_3056),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_3058),
.B(n_53),
.Y(n_3116)
);

HB1xp67_ASAP7_75t_L g3117 ( 
.A(n_3033),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_3022),
.Y(n_3118)
);

INVxp67_ASAP7_75t_L g3119 ( 
.A(n_3059),
.Y(n_3119)
);

INVxp67_ASAP7_75t_L g3120 ( 
.A(n_3062),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_3053),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_3037),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_3028),
.B(n_54),
.Y(n_3123)
);

OR2x6_ASAP7_75t_L g3124 ( 
.A(n_3038),
.B(n_54),
.Y(n_3124)
);

HB1xp67_ASAP7_75t_L g3125 ( 
.A(n_3038),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_3065),
.B(n_55),
.Y(n_3126)
);

INVxp67_ASAP7_75t_SL g3127 ( 
.A(n_3031),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_3040),
.Y(n_3128)
);

INVx2_ASAP7_75t_SL g3129 ( 
.A(n_3043),
.Y(n_3129)
);

INVx1_ASAP7_75t_SL g3130 ( 
.A(n_3069),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_3045),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_3046),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_3047),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_3071),
.B(n_3019),
.Y(n_3134)
);

AOI32xp33_ASAP7_75t_L g3135 ( 
.A1(n_3052),
.A2(n_57),
.A3(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_3017),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_3044),
.B(n_56),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_3036),
.Y(n_3138)
);

AND2x4_ASAP7_75t_L g3139 ( 
.A(n_3055),
.B(n_57),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3060),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_3041),
.B(n_58),
.Y(n_3141)
);

AND2x4_ASAP7_75t_L g3142 ( 
.A(n_3070),
.B(n_59),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3029),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3029),
.Y(n_3144)
);

INVxp67_ASAP7_75t_L g3145 ( 
.A(n_3023),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_3063),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_3067),
.B(n_60),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_3021),
.B(n_61),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_3067),
.B(n_61),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_3067),
.B(n_62),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_3067),
.B(n_62),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3021),
.Y(n_3152)
);

OR2x2_ASAP7_75t_L g3153 ( 
.A(n_3021),
.B(n_64),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_3026),
.B(n_66),
.Y(n_3154)
);

OR2x6_ASAP7_75t_L g3155 ( 
.A(n_3026),
.B(n_67),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_3067),
.B(n_67),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_3021),
.Y(n_3157)
);

OR2x6_ASAP7_75t_L g3158 ( 
.A(n_3026),
.B(n_68),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_3021),
.B(n_68),
.Y(n_3159)
);

OAI22xp33_ASAP7_75t_SL g3160 ( 
.A1(n_3008),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_3160)
);

OAI22xp5_ASAP7_75t_L g3161 ( 
.A1(n_3008),
.A2(n_74),
.B1(n_71),
.B2(n_72),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_3039),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_3021),
.Y(n_3163)
);

OR2x2_ASAP7_75t_SL g3164 ( 
.A(n_3039),
.B(n_72),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_3021),
.B(n_75),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_3067),
.B(n_75),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_3067),
.B(n_76),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_3033),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_3021),
.B(n_76),
.Y(n_3169)
);

AOI22xp33_ASAP7_75t_L g3170 ( 
.A1(n_3117),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_3170)
);

OAI21xp5_ASAP7_75t_L g3171 ( 
.A1(n_3076),
.A2(n_78),
.B(n_80),
.Y(n_3171)
);

AOI21xp33_ASAP7_75t_SL g3172 ( 
.A1(n_3078),
.A2(n_80),
.B(n_81),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_3142),
.B(n_81),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_SL g3174 ( 
.A(n_3160),
.B(n_82),
.Y(n_3174)
);

INVx3_ASAP7_75t_L g3175 ( 
.A(n_3124),
.Y(n_3175)
);

OA22x2_ASAP7_75t_L g3176 ( 
.A1(n_3076),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_3176)
);

OAI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_3168),
.A2(n_84),
.B(n_85),
.Y(n_3177)
);

AOI21xp33_ASAP7_75t_L g3178 ( 
.A1(n_3168),
.A2(n_85),
.B(n_86),
.Y(n_3178)
);

OAI21xp33_ASAP7_75t_L g3179 ( 
.A1(n_3080),
.A2(n_86),
.B(n_88),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3082),
.Y(n_3180)
);

AND2x4_ASAP7_75t_L g3181 ( 
.A(n_3090),
.B(n_89),
.Y(n_3181)
);

NAND3xp33_ASAP7_75t_L g3182 ( 
.A(n_3143),
.B(n_89),
.C(n_90),
.Y(n_3182)
);

INVxp33_ASAP7_75t_L g3183 ( 
.A(n_3125),
.Y(n_3183)
);

OAI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_3144),
.A2(n_90),
.B(n_91),
.Y(n_3184)
);

INVx2_ASAP7_75t_SL g3185 ( 
.A(n_3107),
.Y(n_3185)
);

OAI22xp33_ASAP7_75t_L g3186 ( 
.A1(n_3079),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_3186)
);

NOR2x1_ASAP7_75t_L g3187 ( 
.A(n_3153),
.B(n_94),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3111),
.Y(n_3188)
);

AOI22xp33_ASAP7_75t_L g3189 ( 
.A1(n_3145),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_3189)
);

AOI22xp33_ASAP7_75t_L g3190 ( 
.A1(n_3136),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_3190)
);

NAND3xp33_ASAP7_75t_L g3191 ( 
.A(n_3094),
.B(n_99),
.C(n_100),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3148),
.Y(n_3192)
);

AOI22xp5_ASAP7_75t_SL g3193 ( 
.A1(n_3130),
.A2(n_105),
.B1(n_102),
.B2(n_104),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3159),
.Y(n_3194)
);

INVx2_ASAP7_75t_SL g3195 ( 
.A(n_3112),
.Y(n_3195)
);

AOI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_3137),
.A2(n_106),
.B1(n_102),
.B2(n_104),
.Y(n_3196)
);

OAI21xp33_ASAP7_75t_L g3197 ( 
.A1(n_3162),
.A2(n_106),
.B(n_107),
.Y(n_3197)
);

OAI211xp5_ASAP7_75t_L g3198 ( 
.A1(n_3081),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_3198)
);

AND2x4_ASAP7_75t_L g3199 ( 
.A(n_3095),
.B(n_108),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_3164),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_3124),
.Y(n_3201)
);

OAI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_3122),
.A2(n_114),
.B1(n_111),
.B2(n_113),
.Y(n_3202)
);

NAND3xp33_ASAP7_75t_L g3203 ( 
.A(n_3152),
.B(n_111),
.C(n_113),
.Y(n_3203)
);

OR2x2_ASAP7_75t_L g3204 ( 
.A(n_3157),
.B(n_115),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_3142),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3146),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3165),
.Y(n_3207)
);

OAI21xp33_ASAP7_75t_L g3208 ( 
.A1(n_3127),
.A2(n_3163),
.B(n_3138),
.Y(n_3208)
);

INVxp67_ASAP7_75t_L g3209 ( 
.A(n_3155),
.Y(n_3209)
);

OAI22xp33_ASAP7_75t_SL g3210 ( 
.A1(n_3140),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_3139),
.B(n_119),
.Y(n_3211)
);

AO21x1_ASAP7_75t_L g3212 ( 
.A1(n_3091),
.A2(n_121),
.B(n_122),
.Y(n_3212)
);

OAI22xp33_ASAP7_75t_L g3213 ( 
.A1(n_3100),
.A2(n_124),
.B1(n_121),
.B2(n_123),
.Y(n_3213)
);

OAI22xp33_ASAP7_75t_L g3214 ( 
.A1(n_3085),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_3214)
);

AOI21xp33_ASAP7_75t_SL g3215 ( 
.A1(n_3088),
.A2(n_126),
.B(n_129),
.Y(n_3215)
);

INVx2_ASAP7_75t_SL g3216 ( 
.A(n_3102),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3169),
.Y(n_3217)
);

XOR2x2_ASAP7_75t_L g3218 ( 
.A(n_3110),
.B(n_131),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_3093),
.B(n_3101),
.Y(n_3219)
);

O2A1O1Ixp33_ASAP7_75t_SL g3220 ( 
.A1(n_3129),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_3220)
);

XOR2xp5_ASAP7_75t_L g3221 ( 
.A(n_3096),
.B(n_132),
.Y(n_3221)
);

OAI22xp33_ASAP7_75t_L g3222 ( 
.A1(n_3113),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_3222)
);

OAI21xp33_ASAP7_75t_SL g3223 ( 
.A1(n_3092),
.A2(n_133),
.B(n_134),
.Y(n_3223)
);

XOR2x2_ASAP7_75t_L g3224 ( 
.A(n_3115),
.B(n_3126),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3097),
.Y(n_3225)
);

INVx1_ASAP7_75t_SL g3226 ( 
.A(n_3106),
.Y(n_3226)
);

OAI221xp5_ASAP7_75t_L g3227 ( 
.A1(n_3103),
.A2(n_138),
.B1(n_135),
.B2(n_137),
.C(n_139),
.Y(n_3227)
);

NAND2xp33_ASAP7_75t_SL g3228 ( 
.A(n_3084),
.B(n_139),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3109),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_3119),
.A2(n_3120),
.B1(n_3118),
.B2(n_3141),
.Y(n_3230)
);

INVx2_ASAP7_75t_SL g3231 ( 
.A(n_3105),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3077),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_3155),
.Y(n_3233)
);

O2A1O1Ixp5_ASAP7_75t_L g3234 ( 
.A1(n_3098),
.A2(n_149),
.B(n_161),
.C(n_140),
.Y(n_3234)
);

A2O1A1Ixp33_ASAP7_75t_L g3235 ( 
.A1(n_3135),
.A2(n_785),
.B(n_784),
.C(n_142),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_3086),
.A2(n_3121),
.B1(n_3104),
.B2(n_3108),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3139),
.B(n_140),
.Y(n_3237)
);

NAND4xp25_ASAP7_75t_L g3238 ( 
.A(n_3134),
.B(n_143),
.C(n_141),
.D(n_142),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3114),
.A2(n_141),
.B(n_143),
.Y(n_3239)
);

INVxp67_ASAP7_75t_SL g3240 ( 
.A(n_3154),
.Y(n_3240)
);

OAI22xp5_ASAP7_75t_L g3241 ( 
.A1(n_3161),
.A2(n_147),
.B1(n_144),
.B2(n_146),
.Y(n_3241)
);

OAI22xp33_ASAP7_75t_L g3242 ( 
.A1(n_3116),
.A2(n_147),
.B1(n_144),
.B2(n_146),
.Y(n_3242)
);

OAI221xp5_ASAP7_75t_L g3243 ( 
.A1(n_3158),
.A2(n_151),
.B1(n_148),
.B2(n_150),
.C(n_154),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3147),
.Y(n_3244)
);

O2A1O1Ixp33_ASAP7_75t_R g3245 ( 
.A1(n_3099),
.A2(n_154),
.B(n_148),
.C(n_150),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_3158),
.A2(n_156),
.B(n_157),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3149),
.Y(n_3247)
);

HB1xp67_ASAP7_75t_L g3248 ( 
.A(n_3150),
.Y(n_3248)
);

OAI21xp33_ASAP7_75t_L g3249 ( 
.A1(n_3087),
.A2(n_158),
.B(n_159),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_3083),
.B(n_158),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_3151),
.Y(n_3251)
);

OAI211xp5_ASAP7_75t_SL g3252 ( 
.A1(n_3089),
.A2(n_3128),
.B(n_3131),
.C(n_3132),
.Y(n_3252)
);

AOI22xp5_ASAP7_75t_L g3253 ( 
.A1(n_3167),
.A2(n_163),
.B1(n_159),
.B2(n_162),
.Y(n_3253)
);

AOI211xp5_ASAP7_75t_L g3254 ( 
.A1(n_3156),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_3254)
);

OAI21xp33_ASAP7_75t_L g3255 ( 
.A1(n_3133),
.A2(n_164),
.B(n_165),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3166),
.Y(n_3256)
);

AOI22xp5_ASAP7_75t_L g3257 ( 
.A1(n_3123),
.A2(n_170),
.B1(n_166),
.B2(n_168),
.Y(n_3257)
);

OAI22xp5_ASAP7_75t_L g3258 ( 
.A1(n_3117),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_3258)
);

O2A1O1Ixp33_ASAP7_75t_L g3259 ( 
.A1(n_3117),
.A2(n_174),
.B(n_171),
.C(n_173),
.Y(n_3259)
);

OAI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3117),
.A2(n_174),
.B(n_175),
.Y(n_3260)
);

AOI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_3076),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3164),
.Y(n_3262)
);

OAI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3117),
.A2(n_177),
.B(n_179),
.Y(n_3263)
);

OAI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_3117),
.A2(n_179),
.B(n_180),
.Y(n_3264)
);

OAI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_3117),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_3265)
);

OAI21xp33_ASAP7_75t_L g3266 ( 
.A1(n_3117),
.A2(n_181),
.B(n_182),
.Y(n_3266)
);

OAI22xp33_ASAP7_75t_L g3267 ( 
.A1(n_3076),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_3267)
);

OAI21xp33_ASAP7_75t_L g3268 ( 
.A1(n_3117),
.A2(n_184),
.B(n_187),
.Y(n_3268)
);

AOI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_3076),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_3269)
);

OAI21xp33_ASAP7_75t_L g3270 ( 
.A1(n_3117),
.A2(n_188),
.B(n_189),
.Y(n_3270)
);

AOI21xp5_ASAP7_75t_L g3271 ( 
.A1(n_3117),
.A2(n_190),
.B(n_191),
.Y(n_3271)
);

NOR3xp33_ASAP7_75t_L g3272 ( 
.A(n_3076),
.B(n_190),
.C(n_192),
.Y(n_3272)
);

NAND4xp25_ASAP7_75t_L g3273 ( 
.A(n_3162),
.B(n_196),
.C(n_193),
.D(n_194),
.Y(n_3273)
);

OA22x2_ASAP7_75t_L g3274 ( 
.A1(n_3076),
.A2(n_197),
.B1(n_193),
.B2(n_194),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3082),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3117),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_3276)
);

OAI31xp33_ASAP7_75t_L g3277 ( 
.A1(n_3117),
.A2(n_200),
.A3(n_198),
.B(n_199),
.Y(n_3277)
);

AOI22xp5_ASAP7_75t_L g3278 ( 
.A1(n_3076),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3082),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3164),
.Y(n_3280)
);

OR2x2_ASAP7_75t_L g3281 ( 
.A(n_3082),
.B(n_201),
.Y(n_3281)
);

OAI22xp5_ASAP7_75t_L g3282 ( 
.A1(n_3117),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_3282)
);

OAI22xp33_ASAP7_75t_SL g3283 ( 
.A1(n_3076),
.A2(n_206),
.B1(n_203),
.B2(n_205),
.Y(n_3283)
);

AOI31xp33_ASAP7_75t_L g3284 ( 
.A1(n_3078),
.A2(n_208),
.A3(n_206),
.B(n_207),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3082),
.Y(n_3285)
);

OAI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_3117),
.A2(n_208),
.B(n_209),
.Y(n_3286)
);

AOI22xp5_ASAP7_75t_L g3287 ( 
.A1(n_3076),
.A2(n_213),
.B1(n_210),
.B2(n_211),
.Y(n_3287)
);

OAI31xp33_ASAP7_75t_L g3288 ( 
.A1(n_3117),
.A2(n_214),
.A3(n_210),
.B(n_213),
.Y(n_3288)
);

OAI211xp5_ASAP7_75t_SL g3289 ( 
.A1(n_3076),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_3289)
);

INVx2_ASAP7_75t_SL g3290 ( 
.A(n_3078),
.Y(n_3290)
);

OAI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_3117),
.A2(n_216),
.B(n_218),
.Y(n_3291)
);

CKINVDCx16_ASAP7_75t_R g3292 ( 
.A(n_3082),
.Y(n_3292)
);

AOI22x1_ASAP7_75t_L g3293 ( 
.A1(n_3082),
.A2(n_221),
.B1(n_218),
.B2(n_220),
.Y(n_3293)
);

AOI22xp5_ASAP7_75t_L g3294 ( 
.A1(n_3076),
.A2(n_223),
.B1(n_220),
.B2(n_222),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_3117),
.A2(n_223),
.B(n_224),
.Y(n_3295)
);

OAI22xp5_ASAP7_75t_L g3296 ( 
.A1(n_3117),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_3296)
);

XOR2x2_ASAP7_75t_L g3297 ( 
.A(n_3078),
.B(n_227),
.Y(n_3297)
);

OAI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3076),
.A2(n_229),
.B1(n_226),
.B2(n_228),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3164),
.Y(n_3299)
);

HB1xp67_ASAP7_75t_L g3300 ( 
.A(n_3117),
.Y(n_3300)
);

AO21x1_ASAP7_75t_L g3301 ( 
.A1(n_3076),
.A2(n_228),
.B(n_229),
.Y(n_3301)
);

AOI21xp33_ASAP7_75t_L g3302 ( 
.A1(n_3117),
.A2(n_230),
.B(n_231),
.Y(n_3302)
);

AOI22xp5_ASAP7_75t_L g3303 ( 
.A1(n_3076),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3164),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_3082),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3082),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3082),
.Y(n_3307)
);

NOR2x1_ASAP7_75t_L g3308 ( 
.A(n_3076),
.B(n_233),
.Y(n_3308)
);

AOI22xp33_ASAP7_75t_L g3309 ( 
.A1(n_3117),
.A2(n_237),
.B1(n_234),
.B2(n_235),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3142),
.B(n_234),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3164),
.Y(n_3311)
);

INVxp67_ASAP7_75t_SL g3312 ( 
.A(n_3117),
.Y(n_3312)
);

XOR2x2_ASAP7_75t_L g3313 ( 
.A(n_3078),
.B(n_238),
.Y(n_3313)
);

OAI21xp33_ASAP7_75t_L g3314 ( 
.A1(n_3117),
.A2(n_235),
.B(n_238),
.Y(n_3314)
);

XNOR2xp5_ASAP7_75t_L g3315 ( 
.A(n_3078),
.B(n_239),
.Y(n_3315)
);

AOI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_3076),
.A2(n_242),
.B1(n_239),
.B2(n_240),
.Y(n_3316)
);

OAI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_3117),
.A2(n_243),
.B(n_244),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3164),
.Y(n_3318)
);

A2O1A1Ixp33_ASAP7_75t_L g3319 ( 
.A1(n_3076),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_SL g3320 ( 
.A(n_3160),
.B(n_245),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3117),
.A2(n_250),
.B1(n_246),
.B2(n_249),
.Y(n_3321)
);

O2A1O1Ixp33_ASAP7_75t_SL g3322 ( 
.A1(n_3117),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3082),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3082),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3082),
.Y(n_3325)
);

AOI21xp33_ASAP7_75t_L g3326 ( 
.A1(n_3117),
.A2(n_253),
.B(n_254),
.Y(n_3326)
);

OAI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_3300),
.A2(n_257),
.B1(n_254),
.B2(n_255),
.Y(n_3327)
);

OAI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_3223),
.A2(n_257),
.B(n_258),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3292),
.B(n_259),
.Y(n_3329)
);

INVxp67_ASAP7_75t_L g3330 ( 
.A(n_3248),
.Y(n_3330)
);

AOI222xp33_ASAP7_75t_L g3331 ( 
.A1(n_3312),
.A2(n_3240),
.B1(n_3219),
.B2(n_3308),
.C1(n_3230),
.C2(n_3209),
.Y(n_3331)
);

HB1xp67_ASAP7_75t_L g3332 ( 
.A(n_3315),
.Y(n_3332)
);

OAI221xp5_ASAP7_75t_L g3333 ( 
.A1(n_3271),
.A2(n_262),
.B1(n_259),
.B2(n_261),
.C(n_263),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3176),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3274),
.Y(n_3335)
);

AOI222xp33_ASAP7_75t_L g3336 ( 
.A1(n_3174),
.A2(n_265),
.B1(n_267),
.B2(n_262),
.C1(n_264),
.C2(n_266),
.Y(n_3336)
);

AND2x2_ASAP7_75t_L g3337 ( 
.A(n_3290),
.B(n_264),
.Y(n_3337)
);

AOI21xp5_ASAP7_75t_L g3338 ( 
.A1(n_3322),
.A2(n_266),
.B(n_267),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3183),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_3339)
);

O2A1O1Ixp33_ASAP7_75t_SL g3340 ( 
.A1(n_3180),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_3275),
.B(n_275),
.Y(n_3341)
);

O2A1O1Ixp33_ASAP7_75t_SL g3342 ( 
.A1(n_3279),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_3342)
);

AOI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3220),
.A2(n_3284),
.B(n_3259),
.Y(n_3343)
);

OAI22xp33_ASAP7_75t_SL g3344 ( 
.A1(n_3226),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_3344)
);

AOI22xp5_ASAP7_75t_L g3345 ( 
.A1(n_3200),
.A2(n_281),
.B1(n_278),
.B2(n_279),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_SL g3346 ( 
.A(n_3172),
.B(n_281),
.Y(n_3346)
);

OAI322xp33_ASAP7_75t_L g3347 ( 
.A1(n_3185),
.A2(n_292),
.A3(n_291),
.B1(n_287),
.B2(n_283),
.C1(n_284),
.C2(n_288),
.Y(n_3347)
);

OAI21xp33_ASAP7_75t_L g3348 ( 
.A1(n_3208),
.A2(n_284),
.B(n_288),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3218),
.Y(n_3349)
);

OAI221xp5_ASAP7_75t_L g3350 ( 
.A1(n_3295),
.A2(n_3188),
.B1(n_3263),
.B2(n_3264),
.C(n_3260),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3221),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3212),
.Y(n_3352)
);

OAI21xp5_ASAP7_75t_SL g3353 ( 
.A1(n_3285),
.A2(n_293),
.B(n_294),
.Y(n_3353)
);

AND2x4_ASAP7_75t_L g3354 ( 
.A(n_3195),
.B(n_297),
.Y(n_3354)
);

AOI211xp5_ASAP7_75t_L g3355 ( 
.A1(n_3245),
.A2(n_300),
.B(n_298),
.C(n_299),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3181),
.B(n_298),
.Y(n_3356)
);

INVx1_ASAP7_75t_SL g3357 ( 
.A(n_3297),
.Y(n_3357)
);

NAND3xp33_ASAP7_75t_L g3358 ( 
.A(n_3272),
.B(n_299),
.C(n_300),
.Y(n_3358)
);

OAI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3234),
.A2(n_301),
.B(n_302),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3181),
.B(n_302),
.Y(n_3360)
);

OAI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_3313),
.A2(n_303),
.B(n_304),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3193),
.B(n_303),
.Y(n_3362)
);

OR2x2_ASAP7_75t_L g3363 ( 
.A(n_3281),
.B(n_304),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3301),
.Y(n_3364)
);

BUFx2_ASAP7_75t_L g3365 ( 
.A(n_3305),
.Y(n_3365)
);

NOR2x1_ASAP7_75t_L g3366 ( 
.A(n_3203),
.B(n_305),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3306),
.B(n_305),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3307),
.B(n_306),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_3199),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3199),
.B(n_307),
.Y(n_3370)
);

INVx1_ASAP7_75t_SL g3371 ( 
.A(n_3228),
.Y(n_3371)
);

AOI21xp33_ASAP7_75t_L g3372 ( 
.A1(n_3262),
.A2(n_307),
.B(n_308),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3216),
.B(n_309),
.Y(n_3373)
);

BUFx2_ASAP7_75t_L g3374 ( 
.A(n_3323),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3231),
.B(n_309),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3236),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_3376)
);

NAND3xp33_ASAP7_75t_L g3377 ( 
.A(n_3187),
.B(n_310),
.C(n_311),
.Y(n_3377)
);

AOI211x1_ASAP7_75t_L g3378 ( 
.A1(n_3286),
.A2(n_316),
.B(n_314),
.C(n_315),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3250),
.Y(n_3379)
);

INVxp67_ASAP7_75t_L g3380 ( 
.A(n_3175),
.Y(n_3380)
);

NAND2xp33_ASAP7_75t_SL g3381 ( 
.A(n_3324),
.B(n_315),
.Y(n_3381)
);

OR2x2_ASAP7_75t_L g3382 ( 
.A(n_3325),
.B(n_317),
.Y(n_3382)
);

OAI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_3196),
.A2(n_3269),
.B1(n_3278),
.B2(n_3261),
.Y(n_3383)
);

AOI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3280),
.A2(n_3304),
.B1(n_3311),
.B2(n_3299),
.Y(n_3384)
);

NOR3x1_ASAP7_75t_L g3385 ( 
.A(n_3291),
.B(n_317),
.C(n_318),
.Y(n_3385)
);

INVxp67_ASAP7_75t_L g3386 ( 
.A(n_3175),
.Y(n_3386)
);

AOI22xp5_ASAP7_75t_L g3387 ( 
.A1(n_3318),
.A2(n_3320),
.B1(n_3244),
.B2(n_3247),
.Y(n_3387)
);

CKINVDCx16_ASAP7_75t_R g3388 ( 
.A(n_3232),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3211),
.Y(n_3389)
);

OR2x2_ASAP7_75t_L g3390 ( 
.A(n_3204),
.B(n_319),
.Y(n_3390)
);

HB1xp67_ASAP7_75t_L g3391 ( 
.A(n_3205),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3237),
.Y(n_3392)
);

OAI21xp5_ASAP7_75t_L g3393 ( 
.A1(n_3319),
.A2(n_320),
.B(n_321),
.Y(n_3393)
);

OAI22xp5_ASAP7_75t_L g3394 ( 
.A1(n_3190),
.A2(n_323),
.B1(n_320),
.B2(n_322),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3173),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3310),
.Y(n_3396)
);

AND2x2_ASAP7_75t_SL g3397 ( 
.A(n_3251),
.B(n_322),
.Y(n_3397)
);

INVxp67_ASAP7_75t_L g3398 ( 
.A(n_3233),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3229),
.B(n_324),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3283),
.A2(n_324),
.B(n_326),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3254),
.B(n_326),
.Y(n_3401)
);

OAI22xp5_ASAP7_75t_L g3402 ( 
.A1(n_3191),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3256),
.B(n_327),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3215),
.B(n_328),
.Y(n_3404)
);

O2A1O1Ixp33_ASAP7_75t_SL g3405 ( 
.A1(n_3252),
.A2(n_332),
.B(n_329),
.C(n_331),
.Y(n_3405)
);

OAI221xp5_ASAP7_75t_L g3406 ( 
.A1(n_3317),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_3406)
);

NOR3xp33_ASAP7_75t_L g3407 ( 
.A(n_3302),
.B(n_338),
.C(n_339),
.Y(n_3407)
);

OR2x2_ASAP7_75t_L g3408 ( 
.A(n_3192),
.B(n_339),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3224),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_3210),
.B(n_340),
.Y(n_3410)
);

OR2x2_ASAP7_75t_L g3411 ( 
.A(n_3194),
.B(n_341),
.Y(n_3411)
);

OR2x2_ASAP7_75t_L g3412 ( 
.A(n_3207),
.B(n_341),
.Y(n_3412)
);

AOI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3225),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3239),
.B(n_3246),
.Y(n_3414)
);

NAND2x1_ASAP7_75t_L g3415 ( 
.A(n_3217),
.B(n_342),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3201),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_3416)
);

OAI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_3189),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3417)
);

AOI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_3266),
.A2(n_349),
.B1(n_346),
.B2(n_348),
.Y(n_3418)
);

OAI322xp33_ASAP7_75t_L g3419 ( 
.A1(n_3186),
.A2(n_356),
.A3(n_355),
.B1(n_353),
.B2(n_350),
.C1(n_352),
.C2(n_354),
.Y(n_3419)
);

AOI22xp5_ASAP7_75t_L g3420 ( 
.A1(n_3268),
.A2(n_3270),
.B1(n_3314),
.B2(n_3289),
.Y(n_3420)
);

NOR2xp33_ASAP7_75t_L g3421 ( 
.A(n_3198),
.B(n_352),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3293),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3184),
.B(n_354),
.Y(n_3423)
);

OAI221xp5_ASAP7_75t_L g3424 ( 
.A1(n_3171),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.C(n_358),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3235),
.B(n_357),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3277),
.B(n_358),
.Y(n_3426)
);

AOI211xp5_ASAP7_75t_L g3427 ( 
.A1(n_3326),
.A2(n_362),
.B(n_359),
.C(n_361),
.Y(n_3427)
);

AOI221xp5_ASAP7_75t_L g3428 ( 
.A1(n_3178),
.A2(n_3182),
.B1(n_3276),
.B2(n_3265),
.C(n_3258),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3288),
.B(n_359),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3253),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3243),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_SL g3432 ( 
.A(n_3267),
.B(n_363),
.Y(n_3432)
);

NAND2xp33_ASAP7_75t_L g3433 ( 
.A(n_3179),
.B(n_364),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3257),
.Y(n_3434)
);

OAI31xp33_ASAP7_75t_SL g3435 ( 
.A1(n_3282),
.A2(n_366),
.A3(n_364),
.B(n_365),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3273),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3214),
.B(n_368),
.Y(n_3437)
);

AOI31xp33_ASAP7_75t_L g3438 ( 
.A1(n_3177),
.A2(n_370),
.A3(n_368),
.B(n_369),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3296),
.Y(n_3439)
);

INVx1_ASAP7_75t_SL g3440 ( 
.A(n_3287),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3238),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_3298),
.A2(n_370),
.B(n_371),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3242),
.B(n_372),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3294),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3227),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3303),
.Y(n_3446)
);

AND2x2_ASAP7_75t_L g3447 ( 
.A(n_3249),
.B(n_372),
.Y(n_3447)
);

OAI21xp33_ASAP7_75t_L g3448 ( 
.A1(n_3255),
.A2(n_373),
.B(n_374),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3316),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3241),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_3197),
.B(n_374),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_3170),
.B(n_375),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3391),
.Y(n_3453)
);

NOR2x1p5_ASAP7_75t_L g3454 ( 
.A(n_3422),
.B(n_3309),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_3329),
.B(n_3321),
.Y(n_3455)
);

AOI221x1_ASAP7_75t_L g3456 ( 
.A1(n_3409),
.A2(n_3206),
.B1(n_3202),
.B2(n_3222),
.C(n_3213),
.Y(n_3456)
);

AOI22xp33_ASAP7_75t_L g3457 ( 
.A1(n_3364),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3332),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_SL g3459 ( 
.A(n_3331),
.B(n_377),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3388),
.B(n_378),
.Y(n_3460)
);

OAI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3330),
.A2(n_383),
.B1(n_379),
.B2(n_380),
.Y(n_3461)
);

XOR2x2_ASAP7_75t_L g3462 ( 
.A(n_3357),
.B(n_380),
.Y(n_3462)
);

NOR3xp33_ASAP7_75t_SL g3463 ( 
.A(n_3350),
.B(n_383),
.C(n_384),
.Y(n_3463)
);

OAI221xp5_ASAP7_75t_L g3464 ( 
.A1(n_3352),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.C(n_388),
.Y(n_3464)
);

AND2x4_ASAP7_75t_L g3465 ( 
.A(n_3337),
.B(n_385),
.Y(n_3465)
);

NAND3xp33_ASAP7_75t_L g3466 ( 
.A(n_3381),
.B(n_3387),
.C(n_3386),
.Y(n_3466)
);

CKINVDCx16_ASAP7_75t_R g3467 ( 
.A(n_3361),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3354),
.B(n_386),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3363),
.Y(n_3469)
);

AND2x4_ASAP7_75t_L g3470 ( 
.A(n_3341),
.B(n_387),
.Y(n_3470)
);

OAI211xp5_ASAP7_75t_L g3471 ( 
.A1(n_3365),
.A2(n_390),
.B(n_388),
.C(n_389),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3354),
.B(n_389),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3397),
.B(n_390),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3405),
.A2(n_391),
.B(n_392),
.Y(n_3474)
);

OR2x6_ASAP7_75t_L g3475 ( 
.A(n_3380),
.B(n_392),
.Y(n_3475)
);

AND2x6_ASAP7_75t_L g3476 ( 
.A(n_3367),
.B(n_393),
.Y(n_3476)
);

AOI322xp5_ASAP7_75t_L g3477 ( 
.A1(n_3334),
.A2(n_398),
.A3(n_397),
.B1(n_395),
.B2(n_393),
.C1(n_394),
.C2(n_396),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3390),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3374),
.Y(n_3479)
);

AOI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3335),
.A2(n_397),
.B1(n_394),
.B2(n_396),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3378),
.B(n_398),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3356),
.Y(n_3482)
);

OAI21xp5_ASAP7_75t_SL g3483 ( 
.A1(n_3353),
.A2(n_399),
.B(n_400),
.Y(n_3483)
);

OAI22xp5_ASAP7_75t_L g3484 ( 
.A1(n_3441),
.A2(n_3436),
.B1(n_3420),
.B2(n_3382),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3360),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3340),
.A2(n_399),
.B(n_401),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3399),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3370),
.Y(n_3488)
);

AOI221xp5_ASAP7_75t_L g3489 ( 
.A1(n_3383),
.A2(n_408),
.B1(n_403),
.B2(n_405),
.C(n_410),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3415),
.Y(n_3490)
);

AOI222xp33_ASAP7_75t_L g3491 ( 
.A1(n_3414),
.A2(n_411),
.B1(n_413),
.B2(n_403),
.C1(n_410),
.C2(n_412),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3368),
.B(n_411),
.Y(n_3492)
);

INVxp67_ASAP7_75t_L g3493 ( 
.A(n_3410),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3379),
.Y(n_3494)
);

AOI322xp5_ASAP7_75t_L g3495 ( 
.A1(n_3440),
.A2(n_412),
.A3(n_413),
.B1(n_414),
.B2(n_415),
.C1(n_416),
.C2(n_417),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3378),
.B(n_414),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3408),
.Y(n_3497)
);

OAI21xp33_ASAP7_75t_L g3498 ( 
.A1(n_3348),
.A2(n_415),
.B(n_416),
.Y(n_3498)
);

AOI221xp5_ASAP7_75t_L g3499 ( 
.A1(n_3355),
.A2(n_3359),
.B1(n_3328),
.B2(n_3343),
.C(n_3428),
.Y(n_3499)
);

NOR4xp25_ASAP7_75t_SL g3500 ( 
.A(n_3342),
.B(n_419),
.C(n_417),
.D(n_418),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3338),
.B(n_3371),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3423),
.B(n_418),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3411),
.Y(n_3503)
);

OR2x2_ASAP7_75t_L g3504 ( 
.A(n_3373),
.B(n_420),
.Y(n_3504)
);

AOI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_3346),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_3505)
);

OAI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_3418),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3412),
.Y(n_3507)
);

OR2x2_ASAP7_75t_L g3508 ( 
.A(n_3375),
.B(n_424),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3366),
.B(n_3385),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3369),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3447),
.B(n_426),
.Y(n_3511)
);

OAI22xp33_ASAP7_75t_SL g3512 ( 
.A1(n_3351),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3362),
.Y(n_3513)
);

AOI22xp33_ASAP7_75t_SL g3514 ( 
.A1(n_3349),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_SL g3515 ( 
.A(n_3344),
.B(n_430),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_3433),
.A2(n_430),
.B(n_431),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_3345),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_3517)
);

OAI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_3400),
.A2(n_433),
.B(n_434),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_SL g3519 ( 
.A(n_3336),
.B(n_435),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3404),
.Y(n_3520)
);

OR2x2_ASAP7_75t_L g3521 ( 
.A(n_3403),
.B(n_435),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3401),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3347),
.Y(n_3523)
);

NOR2x1p5_ASAP7_75t_L g3524 ( 
.A(n_3426),
.B(n_436),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3377),
.Y(n_3525)
);

AND2x4_ASAP7_75t_L g3526 ( 
.A(n_3395),
.B(n_436),
.Y(n_3526)
);

OR2x2_ASAP7_75t_L g3527 ( 
.A(n_3376),
.B(n_437),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3450),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3421),
.B(n_437),
.Y(n_3529)
);

O2A1O1Ixp33_ASAP7_75t_L g3530 ( 
.A1(n_3438),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3425),
.Y(n_3531)
);

OR2x2_ASAP7_75t_L g3532 ( 
.A(n_3339),
.B(n_439),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3437),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3429),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3443),
.Y(n_3535)
);

AOI211xp5_ASAP7_75t_L g3536 ( 
.A1(n_3327),
.A2(n_442),
.B(n_440),
.C(n_441),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3419),
.Y(n_3537)
);

INVx1_ASAP7_75t_SL g3538 ( 
.A(n_3452),
.Y(n_3538)
);

NAND4xp25_ASAP7_75t_L g3539 ( 
.A(n_3384),
.B(n_444),
.C(n_442),
.D(n_443),
.Y(n_3539)
);

AOI221xp5_ASAP7_75t_L g3540 ( 
.A1(n_3396),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.C(n_446),
.Y(n_3540)
);

AOI222xp33_ASAP7_75t_L g3541 ( 
.A1(n_3444),
.A2(n_3446),
.B1(n_3449),
.B2(n_3434),
.C1(n_3430),
.C2(n_3398),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_3432),
.A2(n_447),
.B(n_448),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3435),
.B(n_449),
.Y(n_3543)
);

INVx1_ASAP7_75t_SL g3544 ( 
.A(n_3439),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3389),
.Y(n_3545)
);

AND2x2_ASAP7_75t_L g3546 ( 
.A(n_3451),
.B(n_449),
.Y(n_3546)
);

AOI221xp5_ASAP7_75t_L g3547 ( 
.A1(n_3392),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.C(n_453),
.Y(n_3547)
);

INVxp67_ASAP7_75t_L g3548 ( 
.A(n_3333),
.Y(n_3548)
);

AOI221xp5_ASAP7_75t_L g3549 ( 
.A1(n_3393),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.C(n_454),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3427),
.B(n_454),
.Y(n_3550)
);

AOI22xp33_ASAP7_75t_SL g3551 ( 
.A1(n_3431),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3358),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3445),
.Y(n_3553)
);

AOI322xp5_ASAP7_75t_L g3554 ( 
.A1(n_3407),
.A2(n_455),
.A3(n_456),
.B1(n_459),
.B2(n_460),
.C1(n_461),
.C2(n_462),
.Y(n_3554)
);

INVxp67_ASAP7_75t_SL g3555 ( 
.A(n_3416),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3413),
.Y(n_3556)
);

AOI221xp5_ASAP7_75t_L g3557 ( 
.A1(n_3372),
.A2(n_3417),
.B1(n_3448),
.B2(n_3394),
.C(n_3402),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3442),
.B(n_463),
.Y(n_3558)
);

NAND3xp33_ASAP7_75t_L g3559 ( 
.A(n_3406),
.B(n_464),
.C(n_465),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3424),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3391),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3357),
.B(n_464),
.Y(n_3562)
);

OAI211xp5_ASAP7_75t_L g3563 ( 
.A1(n_3330),
.A2(n_467),
.B(n_465),
.C(n_466),
.Y(n_3563)
);

NAND5xp2_ASAP7_75t_L g3564 ( 
.A(n_3331),
.B(n_468),
.C(n_466),
.D(n_467),
.E(n_469),
.Y(n_3564)
);

NOR2xp33_ASAP7_75t_L g3565 ( 
.A(n_3357),
.B(n_468),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3329),
.B(n_469),
.Y(n_3566)
);

BUFx2_ASAP7_75t_SL g3567 ( 
.A(n_3329),
.Y(n_3567)
);

INVxp67_ASAP7_75t_L g3568 ( 
.A(n_3329),
.Y(n_3568)
);

O2A1O1Ixp33_ASAP7_75t_L g3569 ( 
.A1(n_3405),
.A2(n_473),
.B(n_470),
.C(n_472),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3391),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3391),
.Y(n_3571)
);

AOI32xp33_ASAP7_75t_L g3572 ( 
.A1(n_3352),
.A2(n_474),
.A3(n_470),
.B1(n_473),
.B2(n_475),
.Y(n_3572)
);

OAI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3330),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.Y(n_3573)
);

AOI211xp5_ASAP7_75t_L g3574 ( 
.A1(n_3330),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3391),
.Y(n_3575)
);

AOI21xp33_ASAP7_75t_L g3576 ( 
.A1(n_3331),
.A2(n_477),
.B(n_478),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3391),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3391),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3391),
.Y(n_3579)
);

NOR3xp33_ASAP7_75t_L g3580 ( 
.A(n_3409),
.B(n_479),
.C(n_480),
.Y(n_3580)
);

AND2x4_ASAP7_75t_L g3581 ( 
.A(n_3329),
.B(n_481),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3329),
.B(n_481),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_L g3583 ( 
.A(n_3357),
.B(n_482),
.Y(n_3583)
);

AOI22xp33_ASAP7_75t_L g3584 ( 
.A1(n_3364),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_3584)
);

NOR4xp25_ASAP7_75t_L g3585 ( 
.A(n_3364),
.B(n_485),
.C(n_483),
.D(n_484),
.Y(n_3585)
);

OAI221xp5_ASAP7_75t_L g3586 ( 
.A1(n_3409),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.C(n_488),
.Y(n_3586)
);

OAI21xp33_ASAP7_75t_L g3587 ( 
.A1(n_3409),
.A2(n_486),
.B(n_487),
.Y(n_3587)
);

INVxp33_ASAP7_75t_L g3588 ( 
.A(n_3329),
.Y(n_3588)
);

INVxp67_ASAP7_75t_L g3589 ( 
.A(n_3329),
.Y(n_3589)
);

AO32x1_ASAP7_75t_L g3590 ( 
.A1(n_3376),
.A2(n_494),
.A3(n_491),
.B1(n_492),
.B2(n_495),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3391),
.Y(n_3591)
);

OR2x2_ASAP7_75t_L g3592 ( 
.A(n_3388),
.B(n_491),
.Y(n_3592)
);

AOI221xp5_ASAP7_75t_L g3593 ( 
.A1(n_3352),
.A2(n_496),
.B1(n_492),
.B2(n_495),
.C(n_497),
.Y(n_3593)
);

OR2x2_ASAP7_75t_L g3594 ( 
.A(n_3388),
.B(n_496),
.Y(n_3594)
);

AOI211xp5_ASAP7_75t_L g3595 ( 
.A1(n_3330),
.A2(n_500),
.B(n_498),
.C(n_499),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3391),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_SL g3597 ( 
.A(n_3331),
.B(n_499),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3391),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3354),
.B(n_500),
.Y(n_3599)
);

AOI21xp33_ASAP7_75t_L g3600 ( 
.A1(n_3331),
.A2(n_501),
.B(n_502),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3354),
.B(n_501),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3391),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3329),
.B(n_502),
.Y(n_3603)
);

OR2x2_ASAP7_75t_L g3604 ( 
.A(n_3388),
.B(n_503),
.Y(n_3604)
);

AOI321xp33_ASAP7_75t_L g3605 ( 
.A1(n_3409),
.A2(n_503),
.A3(n_504),
.B1(n_505),
.B2(n_506),
.C(n_507),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3391),
.Y(n_3606)
);

INVx1_ASAP7_75t_SL g3607 ( 
.A(n_3329),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3391),
.Y(n_3608)
);

NOR3xp33_ASAP7_75t_L g3609 ( 
.A(n_3576),
.B(n_504),
.C(n_505),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3460),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3476),
.B(n_506),
.Y(n_3611)
);

CKINVDCx20_ASAP7_75t_R g3612 ( 
.A(n_3462),
.Y(n_3612)
);

AOI211xp5_ASAP7_75t_L g3613 ( 
.A1(n_3600),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3567),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3476),
.B(n_510),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3476),
.B(n_510),
.Y(n_3616)
);

INVxp67_ASAP7_75t_L g3617 ( 
.A(n_3564),
.Y(n_3617)
);

OR2x2_ASAP7_75t_L g3618 ( 
.A(n_3592),
.B(n_511),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3594),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3476),
.B(n_511),
.Y(n_3620)
);

AOI221xp5_ASAP7_75t_L g3621 ( 
.A1(n_3459),
.A2(n_514),
.B1(n_512),
.B2(n_513),
.C(n_515),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3604),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_SL g3623 ( 
.A(n_3466),
.B(n_512),
.Y(n_3623)
);

NOR2xp33_ASAP7_75t_L g3624 ( 
.A(n_3588),
.B(n_513),
.Y(n_3624)
);

NOR2xp33_ASAP7_75t_L g3625 ( 
.A(n_3607),
.B(n_516),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3581),
.B(n_516),
.Y(n_3626)
);

NOR2x1_ASAP7_75t_L g3627 ( 
.A(n_3453),
.B(n_517),
.Y(n_3627)
);

INVx1_ASAP7_75t_SL g3628 ( 
.A(n_3566),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3470),
.B(n_517),
.Y(n_3629)
);

NOR3x1_ASAP7_75t_L g3630 ( 
.A(n_3483),
.B(n_518),
.C(n_519),
.Y(n_3630)
);

AOI211xp5_ASAP7_75t_L g3631 ( 
.A1(n_3458),
.A2(n_523),
.B(n_520),
.C(n_522),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3582),
.B(n_520),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3590),
.Y(n_3633)
);

INVxp67_ASAP7_75t_L g3634 ( 
.A(n_3509),
.Y(n_3634)
);

AOI221xp5_ASAP7_75t_L g3635 ( 
.A1(n_3597),
.A2(n_526),
.B1(n_522),
.B2(n_524),
.C(n_527),
.Y(n_3635)
);

NOR3xp33_ASAP7_75t_L g3636 ( 
.A(n_3568),
.B(n_527),
.C(n_528),
.Y(n_3636)
);

NAND3xp33_ASAP7_75t_SL g3637 ( 
.A(n_3500),
.B(n_530),
.C(n_531),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3603),
.B(n_530),
.Y(n_3638)
);

OAI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3474),
.A2(n_531),
.B(n_532),
.Y(n_3639)
);

INVx1_ASAP7_75t_SL g3640 ( 
.A(n_3492),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3590),
.Y(n_3641)
);

INVx1_ASAP7_75t_SL g3642 ( 
.A(n_3544),
.Y(n_3642)
);

NAND4xp25_ASAP7_75t_SL g3643 ( 
.A(n_3479),
.B(n_535),
.C(n_533),
.D(n_534),
.Y(n_3643)
);

NAND3xp33_ASAP7_75t_SL g3644 ( 
.A(n_3585),
.B(n_534),
.C(n_536),
.Y(n_3644)
);

OAI211xp5_ASAP7_75t_L g3645 ( 
.A1(n_3561),
.A2(n_538),
.B(n_536),
.C(n_537),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_3501),
.A2(n_540),
.B(n_541),
.Y(n_3646)
);

NOR2xp33_ASAP7_75t_L g3647 ( 
.A(n_3589),
.B(n_3539),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3570),
.Y(n_3648)
);

AOI21xp5_ASAP7_75t_L g3649 ( 
.A1(n_3486),
.A2(n_540),
.B(n_541),
.Y(n_3649)
);

NOR2x1_ASAP7_75t_L g3650 ( 
.A(n_3571),
.B(n_542),
.Y(n_3650)
);

OAI221xp5_ASAP7_75t_SL g3651 ( 
.A1(n_3499),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.C(n_545),
.Y(n_3651)
);

AOI21xp5_ASAP7_75t_L g3652 ( 
.A1(n_3569),
.A2(n_546),
.B(n_547),
.Y(n_3652)
);

INVxp67_ASAP7_75t_SL g3653 ( 
.A(n_3490),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3575),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3577),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3578),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3579),
.Y(n_3657)
);

OA22x2_ASAP7_75t_L g3658 ( 
.A1(n_3456),
.A2(n_550),
.B1(n_547),
.B2(n_549),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3591),
.Y(n_3659)
);

NAND3xp33_ASAP7_75t_SL g3660 ( 
.A(n_3541),
.B(n_549),
.C(n_550),
.Y(n_3660)
);

NOR2xp67_ASAP7_75t_L g3661 ( 
.A(n_3596),
.B(n_551),
.Y(n_3661)
);

O2A1O1Ixp33_ASAP7_75t_L g3662 ( 
.A1(n_3580),
.A2(n_554),
.B(n_552),
.C(n_553),
.Y(n_3662)
);

NOR2xp33_ASAP7_75t_SL g3663 ( 
.A(n_3598),
.B(n_552),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3465),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3602),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3502),
.B(n_553),
.Y(n_3666)
);

OAI322xp33_ASAP7_75t_L g3667 ( 
.A1(n_3493),
.A2(n_555),
.A3(n_557),
.B1(n_558),
.B2(n_559),
.C1(n_560),
.C2(n_561),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3475),
.Y(n_3668)
);

INVxp67_ASAP7_75t_SL g3669 ( 
.A(n_3606),
.Y(n_3669)
);

NOR2xp67_ASAP7_75t_L g3670 ( 
.A(n_3608),
.B(n_555),
.Y(n_3670)
);

HB1xp67_ASAP7_75t_L g3671 ( 
.A(n_3475),
.Y(n_3671)
);

NAND3xp33_ASAP7_75t_L g3672 ( 
.A(n_3463),
.B(n_558),
.C(n_561),
.Y(n_3672)
);

AOI221xp5_ASAP7_75t_L g3673 ( 
.A1(n_3513),
.A2(n_562),
.B1(n_563),
.B2(n_564),
.C(n_565),
.Y(n_3673)
);

NOR2xp67_ASAP7_75t_L g3674 ( 
.A(n_3494),
.B(n_562),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_SL g3675 ( 
.A(n_3605),
.B(n_563),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3524),
.Y(n_3676)
);

AOI211xp5_ASAP7_75t_L g3677 ( 
.A1(n_3484),
.A2(n_566),
.B(n_564),
.C(n_565),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3468),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3526),
.B(n_567),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3487),
.B(n_568),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3514),
.B(n_568),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_SL g3682 ( 
.A(n_3512),
.B(n_569),
.Y(n_3682)
);

AOI221xp5_ASAP7_75t_L g3683 ( 
.A1(n_3531),
.A2(n_569),
.B1(n_570),
.B2(n_571),
.C(n_572),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3455),
.B(n_570),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3471),
.B(n_571),
.Y(n_3685)
);

NAND2x1_ASAP7_75t_L g3686 ( 
.A(n_3545),
.B(n_572),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_L g3687 ( 
.A(n_3563),
.B(n_573),
.Y(n_3687)
);

OAI211xp5_ASAP7_75t_L g3688 ( 
.A1(n_3587),
.A2(n_578),
.B(n_576),
.C(n_577),
.Y(n_3688)
);

OR2x2_ASAP7_75t_L g3689 ( 
.A(n_3523),
.B(n_576),
.Y(n_3689)
);

OAI221xp5_ASAP7_75t_L g3690 ( 
.A1(n_3518),
.A2(n_578),
.B1(n_579),
.B2(n_580),
.C(n_581),
.Y(n_3690)
);

INVx1_ASAP7_75t_SL g3691 ( 
.A(n_3521),
.Y(n_3691)
);

NOR2x1_ASAP7_75t_L g3692 ( 
.A(n_3472),
.B(n_579),
.Y(n_3692)
);

NOR2xp33_ASAP7_75t_L g3693 ( 
.A(n_3515),
.B(n_580),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3599),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3601),
.Y(n_3695)
);

OAI211xp5_ASAP7_75t_SL g3696 ( 
.A1(n_3537),
.A2(n_584),
.B(n_581),
.C(n_582),
.Y(n_3696)
);

OAI22xp5_ASAP7_75t_L g3697 ( 
.A1(n_3505),
.A2(n_587),
.B1(n_584),
.B2(n_585),
.Y(n_3697)
);

NOR3x1_ASAP7_75t_L g3698 ( 
.A(n_3559),
.B(n_585),
.C(n_588),
.Y(n_3698)
);

NOR3xp33_ASAP7_75t_L g3699 ( 
.A(n_3562),
.B(n_588),
.C(n_589),
.Y(n_3699)
);

NOR2xp33_ASAP7_75t_L g3700 ( 
.A(n_3467),
.B(n_590),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_SL g3701 ( 
.A(n_3565),
.B(n_590),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3481),
.Y(n_3702)
);

OAI322xp33_ASAP7_75t_SL g3703 ( 
.A1(n_3614),
.A2(n_3535),
.A3(n_3534),
.B1(n_3510),
.B2(n_3533),
.C1(n_3528),
.C2(n_3522),
.Y(n_3703)
);

OAI31xp33_ASAP7_75t_L g3704 ( 
.A1(n_3610),
.A2(n_3520),
.A3(n_3454),
.B(n_3525),
.Y(n_3704)
);

AOI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_3642),
.A2(n_3686),
.B(n_3653),
.Y(n_3705)
);

A2O1A1Ixp33_ASAP7_75t_L g3706 ( 
.A1(n_3649),
.A2(n_3583),
.B(n_3542),
.C(n_3530),
.Y(n_3706)
);

AOI221xp5_ASAP7_75t_L g3707 ( 
.A1(n_3644),
.A2(n_3485),
.B1(n_3482),
.B2(n_3488),
.C(n_3497),
.Y(n_3707)
);

NAND2x1_ASAP7_75t_L g3708 ( 
.A(n_3633),
.B(n_3552),
.Y(n_3708)
);

AOI221xp5_ASAP7_75t_L g3709 ( 
.A1(n_3639),
.A2(n_3507),
.B1(n_3503),
.B2(n_3519),
.C(n_3469),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3617),
.B(n_3511),
.Y(n_3710)
);

NAND3xp33_ASAP7_75t_L g3711 ( 
.A(n_3677),
.B(n_3572),
.C(n_3551),
.Y(n_3711)
);

OAI211xp5_ASAP7_75t_L g3712 ( 
.A1(n_3634),
.A2(n_3669),
.B(n_3641),
.C(n_3654),
.Y(n_3712)
);

AOI322xp5_ASAP7_75t_L g3713 ( 
.A1(n_3637),
.A2(n_3555),
.A3(n_3538),
.B1(n_3478),
.B2(n_3556),
.C1(n_3553),
.C2(n_3557),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_SL g3714 ( 
.A(n_3677),
.B(n_3491),
.Y(n_3714)
);

OAI221xp5_ASAP7_75t_L g3715 ( 
.A1(n_3646),
.A2(n_3498),
.B1(n_3480),
.B2(n_3532),
.C(n_3516),
.Y(n_3715)
);

NOR3xp33_ASAP7_75t_L g3716 ( 
.A(n_3660),
.B(n_3586),
.C(n_3464),
.Y(n_3716)
);

AOI222xp33_ASAP7_75t_L g3717 ( 
.A1(n_3628),
.A2(n_3622),
.B1(n_3619),
.B2(n_3640),
.C1(n_3670),
.C2(n_3661),
.Y(n_3717)
);

AOI21xp33_ASAP7_75t_SL g3718 ( 
.A1(n_3658),
.A2(n_3496),
.B(n_3504),
.Y(n_3718)
);

OAI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3648),
.A2(n_3584),
.B1(n_3457),
.B2(n_3527),
.Y(n_3719)
);

OAI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3652),
.A2(n_3548),
.B(n_3560),
.Y(n_3720)
);

NAND2x1_ASAP7_75t_L g3721 ( 
.A(n_3627),
.B(n_3546),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3611),
.Y(n_3722)
);

AOI22xp33_ASAP7_75t_L g3723 ( 
.A1(n_3702),
.A2(n_3676),
.B1(n_3612),
.B2(n_3692),
.Y(n_3723)
);

AOI221xp5_ASAP7_75t_L g3724 ( 
.A1(n_3678),
.A2(n_3543),
.B1(n_3517),
.B2(n_3549),
.C(n_3506),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3615),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_3643),
.A2(n_3675),
.B(n_3623),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_SL g3727 ( 
.A(n_3650),
.B(n_3593),
.Y(n_3727)
);

OAI211xp5_ASAP7_75t_L g3728 ( 
.A1(n_3655),
.A2(n_3574),
.B(n_3595),
.C(n_3477),
.Y(n_3728)
);

AOI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3682),
.A2(n_3473),
.B(n_3550),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_SL g3730 ( 
.A(n_3663),
.B(n_3489),
.Y(n_3730)
);

AOI211xp5_ASAP7_75t_L g3731 ( 
.A1(n_3647),
.A2(n_3461),
.B(n_3573),
.C(n_3529),
.Y(n_3731)
);

A2O1A1Ixp33_ASAP7_75t_SL g3732 ( 
.A1(n_3656),
.A2(n_3536),
.B(n_3558),
.C(n_3495),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_3681),
.A2(n_3508),
.B(n_3540),
.Y(n_3733)
);

OR2x2_ASAP7_75t_L g3734 ( 
.A(n_3657),
.B(n_3554),
.Y(n_3734)
);

AOI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_3645),
.A2(n_3547),
.B(n_591),
.Y(n_3735)
);

NOR2xp33_ASAP7_75t_SL g3736 ( 
.A(n_3651),
.B(n_592),
.Y(n_3736)
);

OAI211xp5_ASAP7_75t_L g3737 ( 
.A1(n_3659),
.A2(n_3665),
.B(n_3635),
.C(n_3621),
.Y(n_3737)
);

OAI221xp5_ASAP7_75t_SL g3738 ( 
.A1(n_3689),
.A2(n_594),
.B1(n_596),
.B2(n_597),
.C(n_598),
.Y(n_3738)
);

AOI21xp33_ASAP7_75t_L g3739 ( 
.A1(n_3691),
.A2(n_3671),
.B(n_3668),
.Y(n_3739)
);

NOR3xp33_ASAP7_75t_L g3740 ( 
.A(n_3700),
.B(n_597),
.C(n_599),
.Y(n_3740)
);

NOR2xp33_ASAP7_75t_L g3741 ( 
.A(n_3696),
.B(n_600),
.Y(n_3741)
);

AOI22xp5_ASAP7_75t_L g3742 ( 
.A1(n_3693),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_3742)
);

AOI221xp5_ASAP7_75t_L g3743 ( 
.A1(n_3694),
.A2(n_601),
.B1(n_602),
.B2(n_603),
.C(n_605),
.Y(n_3743)
);

NOR2xp33_ASAP7_75t_L g3744 ( 
.A(n_3672),
.B(n_3616),
.Y(n_3744)
);

OAI321xp33_ASAP7_75t_L g3745 ( 
.A1(n_3695),
.A2(n_603),
.A3(n_605),
.B1(n_606),
.B2(n_608),
.C(n_609),
.Y(n_3745)
);

NOR2xp33_ASAP7_75t_L g3746 ( 
.A(n_3620),
.B(n_609),
.Y(n_3746)
);

NAND2xp33_ASAP7_75t_SL g3747 ( 
.A(n_3618),
.B(n_610),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3674),
.Y(n_3748)
);

OAI21xp33_ASAP7_75t_SL g3749 ( 
.A1(n_3625),
.A2(n_610),
.B(n_611),
.Y(n_3749)
);

OAI22xp33_ASAP7_75t_L g3750 ( 
.A1(n_3701),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_SL g3751 ( 
.A(n_3631),
.B(n_613),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3680),
.A2(n_3697),
.B(n_3690),
.Y(n_3752)
);

AOI222xp33_ASAP7_75t_L g3753 ( 
.A1(n_3684),
.A2(n_614),
.B1(n_615),
.B2(n_616),
.C1(n_617),
.C2(n_618),
.Y(n_3753)
);

NAND4xp25_ASAP7_75t_SL g3754 ( 
.A(n_3609),
.B(n_617),
.C(n_614),
.D(n_615),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3624),
.A2(n_619),
.B(n_621),
.Y(n_3755)
);

NAND4xp25_ASAP7_75t_L g3756 ( 
.A(n_3698),
.B(n_3630),
.C(n_3613),
.D(n_3664),
.Y(n_3756)
);

OAI211xp5_ASAP7_75t_L g3757 ( 
.A1(n_3688),
.A2(n_622),
.B(n_619),
.C(n_621),
.Y(n_3757)
);

AOI21xp5_ASAP7_75t_L g3758 ( 
.A1(n_3679),
.A2(n_622),
.B(n_623),
.Y(n_3758)
);

AOI221xp5_ASAP7_75t_L g3759 ( 
.A1(n_3685),
.A2(n_624),
.B1(n_625),
.B2(n_626),
.C(n_627),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3632),
.Y(n_3760)
);

OAI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3687),
.A2(n_3662),
.B(n_3636),
.Y(n_3761)
);

NOR3xp33_ASAP7_75t_L g3762 ( 
.A(n_3638),
.B(n_3666),
.C(n_3699),
.Y(n_3762)
);

OAI21xp5_ASAP7_75t_SL g3763 ( 
.A1(n_3683),
.A2(n_625),
.B(n_626),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3708),
.Y(n_3764)
);

A2O1A1Ixp33_ASAP7_75t_SL g3765 ( 
.A1(n_3712),
.A2(n_3626),
.B(n_3629),
.C(n_3667),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3721),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3710),
.Y(n_3767)
);

OAI22xp5_ASAP7_75t_L g3768 ( 
.A1(n_3705),
.A2(n_3673),
.B1(n_628),
.B2(n_629),
.Y(n_3768)
);

AOI22xp5_ASAP7_75t_L g3769 ( 
.A1(n_3744),
.A2(n_627),
.B1(n_629),
.B2(n_630),
.Y(n_3769)
);

AOI22xp5_ASAP7_75t_L g3770 ( 
.A1(n_3719),
.A2(n_631),
.B1(n_632),
.B2(n_633),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3748),
.Y(n_3771)
);

A2O1A1Ixp33_ASAP7_75t_SL g3772 ( 
.A1(n_3704),
.A2(n_631),
.B(n_632),
.C(n_634),
.Y(n_3772)
);

INVx3_ASAP7_75t_L g3773 ( 
.A(n_3734),
.Y(n_3773)
);

BUFx2_ASAP7_75t_L g3774 ( 
.A(n_3749),
.Y(n_3774)
);

O2A1O1Ixp33_ASAP7_75t_SL g3775 ( 
.A1(n_3732),
.A2(n_634),
.B(n_635),
.C(n_637),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3741),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3760),
.Y(n_3777)
);

INVxp33_ASAP7_75t_L g3778 ( 
.A(n_3756),
.Y(n_3778)
);

AOI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_3717),
.A2(n_638),
.B1(n_639),
.B2(n_640),
.Y(n_3779)
);

AND4x1_ASAP7_75t_L g3780 ( 
.A(n_3707),
.B(n_638),
.C(n_639),
.D(n_641),
.Y(n_3780)
);

AOI22xp5_ASAP7_75t_L g3781 ( 
.A1(n_3723),
.A2(n_641),
.B1(n_642),
.B2(n_643),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3722),
.Y(n_3782)
);

AOI22xp5_ASAP7_75t_L g3783 ( 
.A1(n_3762),
.A2(n_643),
.B1(n_644),
.B2(n_645),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3714),
.Y(n_3784)
);

AND4x1_ASAP7_75t_L g3785 ( 
.A(n_3709),
.B(n_644),
.C(n_645),
.D(n_646),
.Y(n_3785)
);

INVxp67_ASAP7_75t_SL g3786 ( 
.A(n_3746),
.Y(n_3786)
);

AOI22xp5_ASAP7_75t_L g3787 ( 
.A1(n_3716),
.A2(n_646),
.B1(n_647),
.B2(n_648),
.Y(n_3787)
);

OAI22xp5_ASAP7_75t_L g3788 ( 
.A1(n_3711),
.A2(n_647),
.B1(n_648),
.B2(n_649),
.Y(n_3788)
);

OAI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3742),
.A2(n_649),
.B1(n_650),
.B2(n_652),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3747),
.Y(n_3790)
);

AOI22xp5_ASAP7_75t_L g3791 ( 
.A1(n_3728),
.A2(n_652),
.B1(n_653),
.B2(n_654),
.Y(n_3791)
);

OAI22xp5_ASAP7_75t_L g3792 ( 
.A1(n_3737),
.A2(n_3738),
.B1(n_3715),
.B2(n_3731),
.Y(n_3792)
);

AOI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3725),
.A2(n_654),
.B1(n_655),
.B2(n_656),
.Y(n_3793)
);

INVx1_ASAP7_75t_SL g3794 ( 
.A(n_3727),
.Y(n_3794)
);

O2A1O1Ixp33_ASAP7_75t_SL g3795 ( 
.A1(n_3706),
.A2(n_3751),
.B(n_3730),
.C(n_3750),
.Y(n_3795)
);

OAI22xp5_ASAP7_75t_L g3796 ( 
.A1(n_3726),
.A2(n_655),
.B1(n_656),
.B2(n_658),
.Y(n_3796)
);

O2A1O1Ixp33_ASAP7_75t_L g3797 ( 
.A1(n_3739),
.A2(n_660),
.B(n_662),
.C(n_663),
.Y(n_3797)
);

AOI221xp5_ASAP7_75t_L g3798 ( 
.A1(n_3718),
.A2(n_663),
.B1(n_664),
.B2(n_665),
.C(n_667),
.Y(n_3798)
);

O2A1O1Ixp33_ASAP7_75t_SL g3799 ( 
.A1(n_3757),
.A2(n_668),
.B(n_670),
.C(n_671),
.Y(n_3799)
);

NOR4xp25_ASAP7_75t_L g3800 ( 
.A(n_3720),
.B(n_668),
.C(n_671),
.D(n_672),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3740),
.Y(n_3801)
);

NOR4xp25_ASAP7_75t_SL g3802 ( 
.A(n_3764),
.B(n_3763),
.C(n_3724),
.D(n_3759),
.Y(n_3802)
);

O2A1O1Ixp33_ASAP7_75t_L g3803 ( 
.A1(n_3772),
.A2(n_3761),
.B(n_3735),
.C(n_3758),
.Y(n_3803)
);

OAI211xp5_ASAP7_75t_L g3804 ( 
.A1(n_3766),
.A2(n_3781),
.B(n_3767),
.C(n_3779),
.Y(n_3804)
);

XOR2xp5_ASAP7_75t_L g3805 ( 
.A(n_3778),
.B(n_3754),
.Y(n_3805)
);

AOI22xp5_ASAP7_75t_L g3806 ( 
.A1(n_3771),
.A2(n_3736),
.B1(n_3729),
.B2(n_3733),
.Y(n_3806)
);

AOI211xp5_ASAP7_75t_L g3807 ( 
.A1(n_3775),
.A2(n_3752),
.B(n_3755),
.C(n_3745),
.Y(n_3807)
);

AOI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3765),
.A2(n_3703),
.B(n_3743),
.Y(n_3808)
);

AOI221xp5_ASAP7_75t_L g3809 ( 
.A1(n_3774),
.A2(n_3773),
.B1(n_3784),
.B2(n_3782),
.C(n_3768),
.Y(n_3809)
);

AOI321xp33_ASAP7_75t_L g3810 ( 
.A1(n_3792),
.A2(n_3713),
.A3(n_3753),
.B1(n_675),
.B2(n_676),
.C(n_677),
.Y(n_3810)
);

NOR3xp33_ASAP7_75t_L g3811 ( 
.A(n_3773),
.B(n_673),
.C(n_674),
.Y(n_3811)
);

AOI211xp5_ASAP7_75t_L g3812 ( 
.A1(n_3797),
.A2(n_675),
.B(n_678),
.C(n_679),
.Y(n_3812)
);

OAI21xp5_ASAP7_75t_SL g3813 ( 
.A1(n_3791),
.A2(n_678),
.B(n_679),
.Y(n_3813)
);

OAI222xp33_ASAP7_75t_L g3814 ( 
.A1(n_3794),
.A2(n_681),
.B1(n_682),
.B2(n_683),
.C1(n_684),
.C2(n_685),
.Y(n_3814)
);

AOI221xp5_ASAP7_75t_L g3815 ( 
.A1(n_3799),
.A2(n_682),
.B1(n_683),
.B2(n_685),
.C(n_687),
.Y(n_3815)
);

OAI221xp5_ASAP7_75t_L g3816 ( 
.A1(n_3798),
.A2(n_687),
.B1(n_688),
.B2(n_689),
.C(n_691),
.Y(n_3816)
);

AOI221xp5_ASAP7_75t_L g3817 ( 
.A1(n_3800),
.A2(n_689),
.B1(n_691),
.B2(n_692),
.C(n_693),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_3786),
.B(n_693),
.Y(n_3818)
);

AOI221xp5_ASAP7_75t_SL g3819 ( 
.A1(n_3777),
.A2(n_695),
.B1(n_696),
.B2(n_697),
.C(n_698),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3785),
.B(n_695),
.Y(n_3820)
);

AOI221x1_ASAP7_75t_L g3821 ( 
.A1(n_3808),
.A2(n_3788),
.B1(n_3796),
.B2(n_3776),
.C(n_3790),
.Y(n_3821)
);

INVxp67_ASAP7_75t_L g3822 ( 
.A(n_3805),
.Y(n_3822)
);

NAND5xp2_ASAP7_75t_L g3823 ( 
.A(n_3810),
.B(n_3795),
.C(n_3801),
.D(n_3770),
.E(n_3787),
.Y(n_3823)
);

INVx1_ASAP7_75t_SL g3824 ( 
.A(n_3818),
.Y(n_3824)
);

OAI22xp33_ASAP7_75t_L g3825 ( 
.A1(n_3806),
.A2(n_3783),
.B1(n_3793),
.B2(n_3769),
.Y(n_3825)
);

AOI221x1_ASAP7_75t_L g3826 ( 
.A1(n_3811),
.A2(n_3789),
.B1(n_3809),
.B2(n_3804),
.C(n_3802),
.Y(n_3826)
);

NAND4xp25_ASAP7_75t_L g3827 ( 
.A(n_3807),
.B(n_3803),
.C(n_3815),
.D(n_3812),
.Y(n_3827)
);

INVxp67_ASAP7_75t_SL g3828 ( 
.A(n_3820),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3814),
.A2(n_3780),
.B(n_696),
.Y(n_3829)
);

NOR2x1_ASAP7_75t_L g3830 ( 
.A(n_3813),
.B(n_697),
.Y(n_3830)
);

OAI221xp5_ASAP7_75t_SL g3831 ( 
.A1(n_3817),
.A2(n_3819),
.B1(n_3816),
.B2(n_700),
.C(n_701),
.Y(n_3831)
);

NOR3xp33_ASAP7_75t_L g3832 ( 
.A(n_3809),
.B(n_698),
.C(n_699),
.Y(n_3832)
);

NOR3xp33_ASAP7_75t_SL g3833 ( 
.A(n_3804),
.B(n_699),
.C(n_702),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3822),
.A2(n_702),
.B(n_703),
.Y(n_3834)
);

AOI21xp33_ASAP7_75t_L g3835 ( 
.A1(n_3824),
.A2(n_703),
.B(n_704),
.Y(n_3835)
);

OAI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3829),
.A2(n_705),
.B(n_706),
.Y(n_3836)
);

CKINVDCx16_ASAP7_75t_R g3837 ( 
.A(n_3830),
.Y(n_3837)
);

A2O1A1Ixp33_ASAP7_75t_L g3838 ( 
.A1(n_3828),
.A2(n_706),
.B(n_707),
.C(n_708),
.Y(n_3838)
);

OAI221xp5_ASAP7_75t_L g3839 ( 
.A1(n_3827),
.A2(n_707),
.B1(n_708),
.B2(n_709),
.C(n_710),
.Y(n_3839)
);

CKINVDCx5p33_ASAP7_75t_R g3840 ( 
.A(n_3833),
.Y(n_3840)
);

INVxp67_ASAP7_75t_L g3841 ( 
.A(n_3823),
.Y(n_3841)
);

INVx1_ASAP7_75t_SL g3842 ( 
.A(n_3826),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3821),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3843),
.B(n_3832),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3842),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3840),
.Y(n_3846)
);

CKINVDCx20_ASAP7_75t_R g3847 ( 
.A(n_3841),
.Y(n_3847)
);

INVxp33_ASAP7_75t_L g3848 ( 
.A(n_3836),
.Y(n_3848)
);

NAND4xp25_ASAP7_75t_L g3849 ( 
.A(n_3845),
.B(n_3831),
.C(n_3834),
.D(n_3835),
.Y(n_3849)
);

NOR3xp33_ASAP7_75t_SL g3850 ( 
.A(n_3846),
.B(n_3837),
.C(n_3825),
.Y(n_3850)
);

AOI221xp5_ASAP7_75t_SL g3851 ( 
.A1(n_3847),
.A2(n_3839),
.B1(n_3838),
.B2(n_713),
.C(n_714),
.Y(n_3851)
);

HB1xp67_ASAP7_75t_L g3852 ( 
.A(n_3849),
.Y(n_3852)
);

OAI22xp5_ASAP7_75t_L g3853 ( 
.A1(n_3852),
.A2(n_3844),
.B1(n_3850),
.B2(n_3848),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3853),
.Y(n_3854)
);

AOI22xp5_ASAP7_75t_L g3855 ( 
.A1(n_3854),
.A2(n_3851),
.B1(n_712),
.B2(n_714),
.Y(n_3855)
);

AOI31xp33_ASAP7_75t_L g3856 ( 
.A1(n_3855),
.A2(n_711),
.A3(n_715),
.B(n_716),
.Y(n_3856)
);

OAI22xp5_ASAP7_75t_SL g3857 ( 
.A1(n_3856),
.A2(n_711),
.B1(n_716),
.B2(n_717),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3857),
.B(n_718),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3858),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3859),
.Y(n_3860)
);

AOI22x1_ASAP7_75t_L g3861 ( 
.A1(n_3860),
.A2(n_719),
.B1(n_720),
.B2(n_722),
.Y(n_3861)
);

AOI221xp5_ASAP7_75t_L g3862 ( 
.A1(n_3861),
.A2(n_719),
.B1(n_720),
.B2(n_722),
.C(n_723),
.Y(n_3862)
);

AOI211xp5_ASAP7_75t_L g3863 ( 
.A1(n_3862),
.A2(n_723),
.B(n_724),
.C(n_725),
.Y(n_3863)
);


endmodule