module fake_jpeg_16985_n_172 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_1),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_35),
.A2(n_44),
.B(n_28),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_5),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_23),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_6),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_6),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_27),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_31),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_31),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_68),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_42),
.B(n_24),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_77),
.B(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_28),
.B1(n_27),
.B2(n_20),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_89)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_15),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_73),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_70),
.B1(n_79),
.B2(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_92),
.B1(n_99),
.B2(n_106),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_58),
.A2(n_26),
.B(n_29),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_97),
.B(n_82),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_90),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_85),
.B(n_66),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_32),
.B1(n_30),
.B2(n_11),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_11),
.B(n_74),
.C(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_101),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_81),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_73),
.B1(n_80),
.B2(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_83),
.B1(n_60),
.B2(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_64),
.B1(n_57),
.B2(n_78),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_102),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_92),
.B(n_91),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_84),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_81),
.C(n_82),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_108),
.C(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_105),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_81),
.C(n_84),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_127),
.B(n_125),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_115),
.B1(n_122),
.B2(n_113),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_95),
.B(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_91),
.B(n_87),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_103),
.C(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_96),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_95),
.B1(n_94),
.B2(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_139),
.B1(n_112),
.B2(n_120),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_143),
.B(n_144),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_142),
.C(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_124),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_120),
.B1(n_112),
.B2(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_118),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_117),
.C(n_126),
.Y(n_142)
);

INVxp33_ASAP7_75t_SL g145 ( 
.A(n_111),
.Y(n_145)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_139),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_135),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_158),
.B(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_163),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_133),
.B(n_148),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_153),
.C(n_147),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_159),
.C(n_160),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_154),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_151),
.B(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_170),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_SL g170 ( 
.A(n_165),
.B(n_151),
.C(n_150),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_169),
.Y(n_172)
);


endmodule