module fake_jpeg_2417_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_42),
.Y(n_95)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_55),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_27),
.B(n_8),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_37),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_30),
.B(n_1),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_27),
.B(n_8),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_16),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_67),
.B(n_71),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_24),
.B1(n_30),
.B2(n_20),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_68),
.A2(n_84),
.B1(n_26),
.B2(n_5),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_39),
.B1(n_18),
.B2(n_38),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_89),
.B1(n_106),
.B2(n_25),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_24),
.B1(n_30),
.B2(n_29),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_40),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_75),
.A2(n_77),
.B(n_105),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_42),
.A2(n_25),
.B1(n_33),
.B2(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_38),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_58),
.B1(n_41),
.B2(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_31),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_15),
.Y(n_91)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_91),
.A2(n_10),
.A3(n_12),
.B1(n_14),
.B2(n_74),
.Y(n_142)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_51),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_53),
.B(n_32),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_33),
.B1(n_21),
.B2(n_40),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_100),
.B1(n_92),
.B2(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_44),
.A2(n_33),
.B1(n_40),
.B2(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_62),
.B(n_18),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_63),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_22),
.B1(n_23),
.B2(n_17),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_33),
.C(n_22),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_14),
.C(n_92),
.Y(n_146)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_118),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_26),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_146),
.C(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_25),
.B1(n_26),
.B2(n_3),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_136),
.B1(n_98),
.B2(n_94),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_145),
.B1(n_87),
.B2(n_69),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_127),
.B(n_141),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_2),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_73),
.B(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_100),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_138)
);

OAI22x1_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_116),
.B1(n_143),
.B2(n_135),
.Y(n_183)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_88),
.A2(n_110),
.B1(n_102),
.B2(n_99),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_102),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_148),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_153),
.B1(n_162),
.B2(n_179),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_117),
.C(n_123),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_88),
.B1(n_65),
.B2(n_85),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_96),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_105),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_122),
.B1(n_130),
.B2(n_141),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_164),
.B(n_173),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_107),
.B1(n_65),
.B2(n_85),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_183),
.B1(n_125),
.B2(n_131),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_166),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_81),
.B(n_111),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_103),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_114),
.B(n_81),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_182),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_69),
.B(n_101),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_79),
.B1(n_101),
.B2(n_147),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_120),
.A2(n_79),
.B1(n_101),
.B2(n_127),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_153),
.B1(n_152),
.B2(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_133),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_113),
.B1(n_140),
.B2(n_121),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_187),
.A2(n_201),
.B1(n_205),
.B2(n_208),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_188),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_209),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_191),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_138),
.B1(n_125),
.B2(n_134),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_194),
.A2(n_149),
.B1(n_170),
.B2(n_177),
.Y(n_236)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_150),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_167),
.A2(n_117),
.B1(n_121),
.B2(n_162),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_166),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_217),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_168),
.B1(n_156),
.B2(n_151),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_161),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_178),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_210),
.B(n_212),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_154),
.B(n_173),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_172),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_171),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_213),
.A2(n_215),
.B(n_199),
.Y(n_222)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_241),
.B(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_197),
.C(n_233),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_176),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_226),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_154),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_183),
.Y(n_231)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_182),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_238),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_200),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_205),
.B1(n_194),
.B2(n_188),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_177),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_193),
.A2(n_166),
.B1(n_213),
.B2(n_198),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_240),
.A2(n_188),
.B1(n_195),
.B2(n_216),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_211),
.A2(n_192),
.B1(n_207),
.B2(n_205),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_203),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_211),
.B(n_207),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_250),
.B(n_230),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_248),
.C(n_256),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_206),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_191),
.B(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_255),
.A2(n_229),
.B1(n_227),
.B2(n_232),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_243),
.C(n_231),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_245),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_263),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_205),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_260),
.C(n_265),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_204),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_227),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_244),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_216),
.C(n_202),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_220),
.A2(n_208),
.B(n_240),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_226),
.B(n_234),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_239),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_239),
.C(n_242),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_247),
.CI(n_249),
.CON(n_269),
.SN(n_269)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_272),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_264),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_274),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_255),
.B(n_246),
.C(n_265),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_280),
.Y(n_298)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_282),
.B(n_257),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_244),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_261),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_250),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_259),
.C(n_252),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_294),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_295),
.C(n_299),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_249),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_297),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_257),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_251),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_280),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_273),
.CI(n_269),
.CON(n_301),
.SN(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_303),
.Y(n_315)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_295),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_305),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_270),
.C(n_277),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_270),
.C(n_271),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_298),
.C(n_291),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_251),
.B(n_272),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_306),
.C(n_310),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_279),
.B1(n_276),
.B2(n_283),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_293),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_282),
.B(n_269),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_312),
.B(n_301),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_289),
.B1(n_252),
.B2(n_275),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_312),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_305),
.C(n_309),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_324),
.Y(n_333)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_323),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_325),
.B(n_326),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_281),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_321),
.A3(n_301),
.B1(n_306),
.B2(n_314),
.C1(n_225),
.C2(n_266),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_328),
.A2(n_315),
.B(n_320),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_322),
.C(n_321),
.Y(n_334)
);

AOI21xp33_ASAP7_75t_L g337 ( 
.A1(n_334),
.A2(n_336),
.B(n_332),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_324),
.C(n_285),
.Y(n_336)
);

AO21x1_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_335),
.B(n_278),
.Y(n_338)
);

AOI321xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_329),
.A3(n_288),
.B1(n_242),
.B2(n_219),
.C(n_237),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_288),
.B(n_219),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_288),
.Y(n_341)
);


endmodule