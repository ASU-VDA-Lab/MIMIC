module real_jpeg_33349_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_18),
.Y(n_23)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NAND2x1p5_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_24),
.B(n_34),
.C(n_37),
.Y(n_33)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_15),
.Y(n_14)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

OAI221xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_24),
.B1(n_30),
.B2(n_32),
.C(n_33),
.Y(n_7)
);

AOI22xp33_ASAP7_75t_SL g8 ( 
.A1(n_9),
.A2(n_10),
.B1(n_20),
.B2(n_23),
.Y(n_8)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_9),
.A2(n_10),
.B1(n_22),
.B2(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_9),
.A2(n_10),
.B1(n_22),
.B2(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NAND2x1_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_19),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_18),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_18),
.Y(n_19)
);

OA21x2_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_14),
.B(n_16),
.Y(n_12)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

OA21x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);


endmodule