module real_aes_9306_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1301;
wire n_1632;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_1584;
wire n_466;
wire n_1277;
wire n_559;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
XNOR2xp5_ASAP7_75t_L g750 ( .A(n_0), .B(n_751), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_1), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_2), .A2(n_78), .B1(n_516), .B2(n_518), .Y(n_515) );
INVx1_ASAP7_75t_L g597 ( .A(n_2), .Y(n_597) );
INVxp67_ASAP7_75t_SL g1609 ( .A(n_3), .Y(n_1609) );
AOI22xp33_ASAP7_75t_L g1627 ( .A1(n_3), .A2(n_44), .B1(n_1628), .B2(n_1629), .Y(n_1627) );
AO22x2_ASAP7_75t_L g1230 ( .A1(n_4), .A2(n_1231), .B1(n_1272), .B2(n_1273), .Y(n_1230) );
INVxp67_ASAP7_75t_L g1272 ( .A(n_4), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_5), .A2(n_238), .B1(n_1073), .B2(n_1075), .Y(n_1072) );
INVx1_ASAP7_75t_L g1114 ( .A(n_5), .Y(n_1114) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_6), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_7), .A2(n_74), .B1(n_1301), .B2(n_1313), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_8), .Y(n_296) );
AND2x2_ASAP7_75t_L g323 ( .A(n_8), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_8), .B(n_217), .Y(n_352) );
INVx1_ASAP7_75t_L g398 ( .A(n_8), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_9), .A2(n_168), .B1(n_832), .B2(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g871 ( .A(n_9), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g780 ( .A1(n_10), .A2(n_197), .B1(n_497), .B2(n_503), .Y(n_780) );
INVx1_ASAP7_75t_L g799 ( .A(n_10), .Y(n_799) );
INVx1_ASAP7_75t_L g1193 ( .A(n_11), .Y(n_1193) );
OAI22xp33_ASAP7_75t_L g1218 ( .A1(n_11), .A2(n_149), .B1(n_971), .B2(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1535 ( .A(n_12), .Y(n_1535) );
OAI221xp5_ASAP7_75t_L g1547 ( .A1(n_12), .A2(n_589), .B1(n_652), .B2(n_1548), .C(n_1550), .Y(n_1547) );
CKINVDCx5p33_ASAP7_75t_R g1085 ( .A(n_13), .Y(n_1085) );
XNOR2x2_ASAP7_75t_L g1136 ( .A(n_14), .B(n_1137), .Y(n_1136) );
AOI22xp5_ASAP7_75t_L g1342 ( .A1(n_14), .A2(n_83), .B1(n_1297), .B2(n_1301), .Y(n_1342) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_15), .Y(n_331) );
AOI21xp33_ASAP7_75t_L g1152 ( .A1(n_16), .A2(n_796), .B(n_797), .Y(n_1152) );
INVx1_ASAP7_75t_L g1175 ( .A(n_16), .Y(n_1175) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_17), .A2(n_236), .B1(n_327), .B2(n_796), .C(n_797), .Y(n_795) );
OAI22xp33_ASAP7_75t_L g804 ( .A1(n_17), .A2(n_95), .B1(n_805), .B2(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g932 ( .A(n_18), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_18), .A2(n_214), .B1(n_524), .B2(n_526), .Y(n_961) );
XNOR2xp5_ASAP7_75t_L g963 ( .A(n_19), .B(n_964), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_20), .A2(n_222), .B1(n_578), .B2(n_657), .C(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g721 ( .A(n_20), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_21), .A2(n_52), .B1(n_1034), .B2(n_1036), .Y(n_1088) );
INVx1_ASAP7_75t_L g1130 ( .A(n_21), .Y(n_1130) );
INVxp67_ASAP7_75t_SL g1185 ( .A(n_22), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_22), .A2(n_255), .B1(n_1207), .B2(n_1214), .Y(n_1213) );
INVx2_ASAP7_75t_L g411 ( .A(n_23), .Y(n_411) );
OR2x2_ASAP7_75t_L g425 ( .A(n_23), .B(n_409), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_24), .A2(n_147), .B1(n_537), .B2(n_541), .Y(n_636) );
INVx1_ASAP7_75t_L g665 ( .A(n_24), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_25), .A2(n_232), .B1(n_524), .B2(n_526), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_25), .A2(n_232), .B1(n_610), .B2(n_612), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_26), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_27), .A2(n_179), .B1(n_612), .B2(n_785), .Y(n_1160) );
INVx1_ASAP7_75t_L g1171 ( .A(n_27), .Y(n_1171) );
AOI22xp33_ASAP7_75t_SL g1200 ( .A1(n_28), .A2(n_87), .B1(n_990), .B2(n_1201), .Y(n_1200) );
INVxp33_ASAP7_75t_L g1226 ( .A(n_28), .Y(n_1226) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_29), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g1341 ( .A1(n_30), .A2(n_141), .B1(n_1285), .B2(n_1293), .Y(n_1341) );
INVx1_ASAP7_75t_L g322 ( .A(n_31), .Y(n_322) );
OR2x2_ASAP7_75t_L g351 ( .A(n_31), .B(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g363 ( .A(n_31), .Y(n_363) );
BUFx2_ASAP7_75t_L g405 ( .A(n_31), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g1051 ( .A1(n_32), .A2(n_209), .B1(n_712), .B2(n_992), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_32), .A2(n_209), .B1(n_510), .B2(n_747), .Y(n_1055) );
INVx1_ASAP7_75t_L g977 ( .A(n_33), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_33), .A2(n_208), .B1(n_990), .B2(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g1333 ( .A(n_34), .Y(n_1333) );
AOI221xp5_ASAP7_75t_L g1559 ( .A1(n_35), .A2(n_138), .B1(n_699), .B2(n_796), .C(n_797), .Y(n_1559) );
OAI22xp33_ASAP7_75t_L g1565 ( .A1(n_35), .A2(n_103), .B1(n_805), .B2(n_807), .Y(n_1565) );
INVx1_ASAP7_75t_L g1190 ( .A(n_36), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_36), .A2(n_72), .B1(n_837), .B2(n_1211), .Y(n_1210) );
OAI221xp5_ASAP7_75t_L g1239 ( .A1(n_37), .A2(n_245), .B1(n_971), .B2(n_1240), .C(n_1241), .Y(n_1239) );
INVx1_ASAP7_75t_L g1248 ( .A(n_37), .Y(n_1248) );
INVx1_ASAP7_75t_L g774 ( .A(n_38), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_38), .A2(n_82), .B1(n_612), .B2(n_785), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_39), .A2(n_69), .B1(n_297), .B2(n_940), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_39), .A2(n_184), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_40), .A2(n_66), .B1(n_361), .B2(n_709), .C(n_710), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_40), .A2(n_66), .B1(n_518), .B2(n_741), .Y(n_740) );
OAI22xp33_ASAP7_75t_L g1161 ( .A1(n_41), .A2(n_48), .B1(n_563), .B2(n_589), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_41), .A2(n_48), .B1(n_840), .B2(n_982), .C(n_1169), .Y(n_1168) );
OAI22xp33_ASAP7_75t_L g1542 ( .A1(n_42), .A2(n_65), .B1(n_497), .B2(n_503), .Y(n_1542) );
INVx1_ASAP7_75t_L g1562 ( .A(n_42), .Y(n_1562) );
INVx1_ASAP7_75t_L g1391 ( .A(n_43), .Y(n_1391) );
INVxp67_ASAP7_75t_SL g1612 ( .A(n_44), .Y(n_1612) );
INVx1_ASAP7_75t_L g794 ( .A(n_45), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_45), .A2(n_236), .B1(n_541), .B2(n_803), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_46), .A2(n_239), .B1(n_981), .B2(n_982), .Y(n_980) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_46), .A2(n_239), .B1(n_996), .B2(n_1002), .Y(n_1001) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_47), .B(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_49), .A2(n_256), .B1(n_1079), .B2(n_1614), .Y(n_1613) );
AOI221xp5_ASAP7_75t_SL g1623 ( .A1(n_49), .A2(n_506), .B1(n_1624), .B2(n_1625), .C(n_1630), .Y(n_1623) );
CKINVDCx5p33_ASAP7_75t_R g1141 ( .A(n_50), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_51), .A2(n_277), .B1(n_712), .B2(n_713), .Y(n_948) );
AOI22xp33_ASAP7_75t_SL g957 ( .A1(n_51), .A2(n_277), .B1(n_512), .B2(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g1080 ( .A(n_52), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_53), .A2(n_89), .B1(n_990), .B2(n_1199), .Y(n_1198) );
AOI22xp33_ASAP7_75t_SL g1206 ( .A1(n_53), .A2(n_89), .B1(n_1207), .B2(n_1208), .Y(n_1206) );
OAI211xp5_ASAP7_75t_L g1583 ( .A1(n_54), .A2(n_1029), .B(n_1584), .C(n_1586), .Y(n_1583) );
INVx1_ASAP7_75t_L g1606 ( .A(n_54), .Y(n_1606) );
CKINVDCx5p33_ASAP7_75t_R g1099 ( .A(n_55), .Y(n_1099) );
INVx1_ASAP7_75t_L g889 ( .A(n_56), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_56), .A2(n_156), .B1(n_606), .B2(n_950), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_57), .A2(n_240), .B1(n_904), .B2(n_971), .Y(n_970) );
OAI22xp33_ASAP7_75t_L g1011 ( .A1(n_57), .A2(n_240), .B1(n_927), .B2(n_1012), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_58), .A2(n_173), .B1(n_610), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_58), .A2(n_173), .B1(n_682), .B2(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g628 ( .A(n_59), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g1143 ( .A(n_60), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_61), .A2(n_110), .B1(n_1285), .B2(n_1293), .Y(n_1284) );
INVx1_ASAP7_75t_L g782 ( .A(n_62), .Y(n_782) );
INVx1_ASAP7_75t_L g1538 ( .A(n_63), .Y(n_1538) );
OAI211xp5_ASAP7_75t_L g1554 ( .A1(n_63), .A2(n_563), .B(n_1555), .C(n_1560), .Y(n_1554) );
INVx1_ASAP7_75t_L g823 ( .A(n_64), .Y(n_823) );
AOI221xp5_ASAP7_75t_L g854 ( .A1(n_64), .A2(n_67), .B1(n_657), .B2(n_855), .C(n_857), .Y(n_854) );
INVx1_ASAP7_75t_L g1561 ( .A(n_65), .Y(n_1561) );
INVx1_ASAP7_75t_L g821 ( .A(n_67), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_68), .A2(n_100), .B1(n_996), .B2(n_1203), .Y(n_1202) );
INVxp67_ASAP7_75t_SL g1217 ( .A(n_68), .Y(n_1217) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_69), .A2(n_235), .B1(n_1034), .B2(n_1036), .Y(n_1033) );
INVx1_ASAP7_75t_L g901 ( .A(n_70), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_70), .A2(n_123), .B1(n_710), .B2(n_953), .Y(n_952) );
CKINVDCx5p33_ASAP7_75t_R g1148 ( .A(n_71), .Y(n_1148) );
INVxp33_ASAP7_75t_L g1187 ( .A(n_72), .Y(n_1187) );
CKINVDCx16_ASAP7_75t_R g689 ( .A(n_73), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_75), .A2(n_589), .B1(n_641), .B2(n_646), .C(n_652), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_75), .A2(n_278), .B1(n_516), .B2(n_522), .Y(n_680) );
INVx1_ASAP7_75t_L g314 ( .A(n_76), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_76), .A2(n_140), .B1(n_438), .B2(n_439), .C(n_444), .Y(n_437) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_77), .Y(n_547) );
INVx1_ASAP7_75t_L g594 ( .A(n_78), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_79), .A2(n_249), .B1(n_521), .B2(n_522), .Y(n_520) );
OAI211xp5_ASAP7_75t_SL g562 ( .A1(n_79), .A2(n_563), .B(n_568), .C(n_583), .Y(n_562) );
INVx1_ASAP7_75t_L g1246 ( .A(n_80), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_80), .A2(n_224), .B1(n_549), .B2(n_739), .Y(n_1271) );
AOI22xp5_ASAP7_75t_L g1315 ( .A1(n_81), .A2(n_122), .B1(n_1285), .B2(n_1293), .Y(n_1315) );
INVx1_ASAP7_75t_L g777 ( .A(n_82), .Y(n_777) );
INVx1_ASAP7_75t_L g645 ( .A(n_84), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_84), .A2(n_219), .B1(n_677), .B2(n_678), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_85), .A2(n_233), .B1(n_990), .B2(n_1259), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_85), .A2(n_233), .B1(n_739), .B2(n_1207), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_86), .A2(n_129), .B1(n_587), .B2(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g733 ( .A(n_86), .Y(n_733) );
INVxp67_ASAP7_75t_SL g1227 ( .A(n_87), .Y(n_1227) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_88), .A2(n_130), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g1052 ( .A1(n_88), .A2(n_130), .B1(n_694), .B2(n_992), .Y(n_1052) );
XNOR2x2_ASAP7_75t_L g880 ( .A(n_90), .B(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g1028 ( .A(n_91), .Y(n_1028) );
OAI222xp33_ASAP7_75t_L g1040 ( .A1(n_91), .A2(n_184), .B1(n_198), .B2(n_1041), .C1(n_1042), .C2(n_1043), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_92), .A2(n_177), .B1(n_843), .B2(n_844), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_92), .A2(n_177), .B1(n_610), .B2(n_669), .Y(n_876) );
INVx1_ASAP7_75t_L g539 ( .A(n_93), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_93), .A2(n_193), .B1(n_578), .B2(n_580), .C(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g1541 ( .A(n_94), .Y(n_1541) );
OAI22xp5_ASAP7_75t_L g1546 ( .A1(n_94), .A2(n_154), .B1(n_612), .B2(n_785), .Y(n_1546) );
INVx1_ASAP7_75t_L g793 ( .A(n_95), .Y(n_793) );
INVx1_ASAP7_75t_L g368 ( .A(n_96), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_96), .A2(n_274), .B1(n_468), .B2(n_472), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g1107 ( .A(n_97), .Y(n_1107) );
INVx1_ASAP7_75t_L g409 ( .A(n_98), .Y(n_409) );
INVx1_ASAP7_75t_L g455 ( .A(n_98), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_99), .A2(n_171), .B1(n_982), .B2(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1018 ( .A(n_99), .Y(n_1018) );
INVxp33_ASAP7_75t_L g1223 ( .A(n_100), .Y(n_1223) );
INVx1_ASAP7_75t_L g1587 ( .A(n_101), .Y(n_1587) );
AOI22xp33_ASAP7_75t_SL g984 ( .A1(n_102), .A2(n_143), .B1(n_833), .B2(n_843), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_102), .A2(n_143), .B1(n_694), .B2(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1556 ( .A(n_103), .Y(n_1556) );
INVx1_ASAP7_75t_L g705 ( .A(n_104), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_104), .A2(n_105), .B1(n_438), .B2(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g706 ( .A(n_105), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_106), .A2(n_244), .B1(n_694), .B2(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g724 ( .A(n_106), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_107), .A2(n_126), .B1(n_1285), .B2(n_1293), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_108), .A2(n_221), .B1(n_1285), .B2(n_1293), .Y(n_1304) );
AOI22xp5_ASAP7_75t_L g1296 ( .A1(n_109), .A2(n_146), .B1(n_1297), .B2(n_1301), .Y(n_1296) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_111), .Y(n_1106) );
INVx1_ASAP7_75t_L g1321 ( .A(n_112), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_113), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_114), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_115), .A2(n_190), .B1(n_510), .B2(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g601 ( .A(n_115), .Y(n_601) );
INVx1_ASAP7_75t_L g700 ( .A(n_116), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_116), .A2(n_262), .B1(n_741), .B2(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g967 ( .A(n_117), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_117), .A2(n_203), .B1(n_699), .B2(n_996), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g1087 ( .A(n_118), .B(n_1032), .Y(n_1087) );
INVx1_ASAP7_75t_L g1128 ( .A(n_118), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_119), .A2(n_273), .B1(n_996), .B2(n_1197), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_119), .A2(n_273), .B1(n_969), .B2(n_981), .Y(n_1209) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_120), .Y(n_828) );
OAI211xp5_ASAP7_75t_L g1592 ( .A1(n_121), .A2(n_369), .B(n_1077), .C(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g1620 ( .A(n_121), .Y(n_1620) );
INVx1_ASAP7_75t_L g884 ( .A(n_123), .Y(n_884) );
INVx1_ASAP7_75t_L g288 ( .A(n_124), .Y(n_288) );
OA22x2_ASAP7_75t_L g1067 ( .A1(n_125), .A2(n_1068), .B1(n_1134), .B2(n_1135), .Y(n_1067) );
INVxp67_ASAP7_75t_SL g1135 ( .A(n_125), .Y(n_1135) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_127), .Y(n_974) );
AO22x1_ASAP7_75t_SL g1318 ( .A1(n_128), .A2(n_229), .B1(n_1285), .B2(n_1293), .Y(n_1318) );
INVx1_ASAP7_75t_L g734 ( .A(n_129), .Y(n_734) );
INVx1_ASAP7_75t_L g1389 ( .A(n_131), .Y(n_1389) );
AO221x2_ASAP7_75t_L g1327 ( .A1(n_132), .A2(n_267), .B1(n_1313), .B2(n_1328), .C(n_1329), .Y(n_1327) );
OAI22xp5_ASAP7_75t_L g1589 ( .A1(n_133), .A2(n_206), .B1(n_1031), .B2(n_1034), .Y(n_1589) );
INVx1_ASAP7_75t_L g1600 ( .A(n_133), .Y(n_1600) );
INVx1_ASAP7_75t_L g1242 ( .A(n_134), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_134), .A2(n_151), .B1(n_918), .B2(n_996), .Y(n_1264) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_135), .Y(n_417) );
XNOR2xp5_ASAP7_75t_L g814 ( .A(n_136), .B(n_815), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_137), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g1564 ( .A1(n_138), .A2(n_167), .B1(n_541), .B2(n_803), .Y(n_1564) );
INVx1_ASAP7_75t_L g920 ( .A(n_139), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_139), .A2(n_218), .B1(n_516), .B2(n_518), .Y(n_960) );
INVx1_ASAP7_75t_L g336 ( .A(n_140), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_142), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g1158 ( .A(n_144), .Y(n_1158) );
OAI221xp5_ASAP7_75t_L g1172 ( .A1(n_144), .A2(n_497), .B1(n_503), .B2(n_530), .C(n_1173), .Y(n_1172) );
XOR2xp5_ASAP7_75t_L g624 ( .A(n_145), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g655 ( .A(n_147), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g1528 ( .A(n_148), .Y(n_1528) );
INVxp67_ASAP7_75t_SL g1191 ( .A(n_149), .Y(n_1191) );
INVx1_ASAP7_75t_L g1255 ( .A(n_150), .Y(n_1255) );
AOI22xp33_ASAP7_75t_SL g1269 ( .A1(n_150), .A2(n_153), .B1(n_982), .B2(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1234 ( .A(n_151), .Y(n_1234) );
INVx1_ASAP7_75t_L g635 ( .A(n_152), .Y(n_635) );
INVx1_ASAP7_75t_L g1250 ( .A(n_153), .Y(n_1250) );
INVx1_ASAP7_75t_L g1540 ( .A(n_154), .Y(n_1540) );
INVx1_ASAP7_75t_L g634 ( .A(n_155), .Y(n_634) );
INVx1_ASAP7_75t_L g898 ( .A(n_156), .Y(n_898) );
INVx1_ASAP7_75t_L g629 ( .A(n_157), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_158), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_159), .A2(n_246), .B1(n_844), .B2(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1014 ( .A(n_159), .Y(n_1014) );
AOI22xp5_ASAP7_75t_L g1305 ( .A1(n_160), .A2(n_259), .B1(n_1297), .B2(n_1301), .Y(n_1305) );
INVx1_ASAP7_75t_L g1046 ( .A(n_161), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_161), .A2(n_166), .B1(n_524), .B2(n_526), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_162), .A2(n_196), .B1(n_857), .B2(n_918), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_162), .A2(n_196), .B1(n_981), .B2(n_982), .Y(n_1267) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_163), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_164), .A2(n_194), .B1(n_697), .B2(n_947), .Y(n_946) );
AOI22xp33_ASAP7_75t_SL g959 ( .A1(n_164), .A2(n_194), .B1(n_518), .B2(n_673), .Y(n_959) );
XOR2xp5_ASAP7_75t_L g1521 ( .A(n_165), .B(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1047 ( .A(n_166), .Y(n_1047) );
INVx1_ASAP7_75t_L g1558 ( .A(n_167), .Y(n_1558) );
INVx1_ASAP7_75t_L g873 ( .A(n_168), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g1529 ( .A(n_169), .Y(n_1529) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_170), .A2(n_227), .B1(n_837), .B2(n_838), .Y(n_836) );
INVx1_ASAP7_75t_L g864 ( .A(n_170), .Y(n_864) );
INVx1_ASAP7_75t_L g1010 ( .A(n_171), .Y(n_1010) );
INVx1_ASAP7_75t_L g649 ( .A(n_172), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_172), .A2(n_200), .B1(n_673), .B2(n_675), .Y(n_672) );
AOI22x1_ASAP7_75t_SL g1020 ( .A1(n_174), .A2(n_1021), .B1(n_1061), .B2(n_1062), .Y(n_1020) );
INVx1_ASAP7_75t_L g1061 ( .A(n_174), .Y(n_1061) );
INVx1_ASAP7_75t_L g552 ( .A(n_175), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_176), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_178), .Y(n_824) );
INVx1_ASAP7_75t_L g1170 ( .A(n_179), .Y(n_1170) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_180), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_181), .A2(n_250), .B1(n_1301), .B2(n_1313), .Y(n_1316) );
INVx1_ASAP7_75t_L g1025 ( .A(n_182), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_182), .A2(n_235), .B1(n_918), .B2(n_947), .Y(n_1053) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_183), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_183), .B(n_288), .Y(n_1292) );
AND3x2_ASAP7_75t_L g1298 ( .A(n_183), .B(n_288), .C(n_1289), .Y(n_1298) );
OAI22xp33_ASAP7_75t_L g1582 ( .A1(n_185), .A2(n_234), .B1(n_1032), .B2(n_1036), .Y(n_1582) );
OAI22xp33_ASAP7_75t_L g1596 ( .A1(n_185), .A2(n_215), .B1(n_297), .B2(n_940), .Y(n_1596) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_186), .Y(n_1081) );
INVx2_ASAP7_75t_L g301 ( .A(n_187), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_188), .Y(n_1237) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_189), .Y(n_760) );
INVx1_ASAP7_75t_L g604 ( .A(n_190), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_191), .A2(n_213), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_191), .A2(n_213), .B1(n_737), .B2(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g1531 ( .A(n_192), .Y(n_1531) );
AOI21xp33_ASAP7_75t_L g1552 ( .A1(n_192), .A2(n_361), .B(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g544 ( .A(n_193), .Y(n_544) );
INVx1_ASAP7_75t_L g1323 ( .A(n_195), .Y(n_1323) );
INVx1_ASAP7_75t_L g800 ( .A(n_197), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_198), .Y(n_1027) );
INVx1_ASAP7_75t_L g902 ( .A(n_199), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_199), .A2(n_231), .B1(n_925), .B2(n_927), .Y(n_924) );
INVx1_ASAP7_75t_L g651 ( .A(n_200), .Y(n_651) );
INVx1_ASAP7_75t_L g1289 ( .A(n_201), .Y(n_1289) );
INVx1_ASAP7_75t_L g846 ( .A(n_202), .Y(n_846) );
INVx1_ASAP7_75t_L g973 ( .A(n_203), .Y(n_973) );
CKINVDCx16_ASAP7_75t_R g1179 ( .A(n_204), .Y(n_1179) );
INVx1_ASAP7_75t_L g1544 ( .A(n_205), .Y(n_1544) );
INVx1_ASAP7_75t_L g1605 ( .A(n_206), .Y(n_1605) );
INVx1_ASAP7_75t_L g769 ( .A(n_207), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g786 ( .A1(n_207), .A2(n_589), .B1(n_652), .B2(n_787), .C(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g976 ( .A(n_208), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g1591 ( .A1(n_210), .A2(n_271), .B1(n_1073), .B2(n_1075), .Y(n_1591) );
AOI22xp33_ASAP7_75t_L g1621 ( .A1(n_210), .A2(n_271), .B1(n_1207), .B2(n_1622), .Y(n_1621) );
AOI22xp33_ASAP7_75t_SL g1050 ( .A1(n_211), .A2(n_253), .B1(n_918), .B2(n_955), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_211), .A2(n_253), .B1(n_516), .B2(n_522), .Y(n_1056) );
INVx1_ASAP7_75t_L g375 ( .A(n_212), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_212), .A2(n_272), .B1(n_438), .B2(n_463), .C(n_465), .Y(n_462) );
INVx1_ASAP7_75t_L g935 ( .A(n_214), .Y(n_935) );
INVx1_ASAP7_75t_L g1617 ( .A(n_215), .Y(n_1617) );
CKINVDCx20_ASAP7_75t_R g1330 ( .A(n_216), .Y(n_1330) );
INVx1_ASAP7_75t_L g303 ( .A(n_217), .Y(n_303) );
INVx2_ASAP7_75t_L g324 ( .A(n_217), .Y(n_324) );
INVx1_ASAP7_75t_L g938 ( .A(n_218), .Y(n_938) );
INVx1_ASAP7_75t_L g643 ( .A(n_219), .Y(n_643) );
INVx1_ASAP7_75t_L g1145 ( .A(n_220), .Y(n_1145) );
AOI221xp5_ASAP7_75t_L g1164 ( .A1(n_220), .A2(n_247), .B1(n_982), .B2(n_1165), .C(n_1167), .Y(n_1164) );
INVx1_ASAP7_75t_L g725 ( .A(n_222), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g1071 ( .A(n_223), .Y(n_1071) );
INVx1_ASAP7_75t_L g1245 ( .A(n_224), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1385 ( .A1(n_225), .A2(n_226), .B1(n_1386), .B2(n_1387), .C(n_1388), .Y(n_1385) );
XNOR2x1_ASAP7_75t_L g309 ( .A(n_226), .B(n_310), .Y(n_309) );
XNOR2xp5_ASAP7_75t_L g617 ( .A(n_226), .B(n_310), .Y(n_617) );
INVx1_ASAP7_75t_L g867 ( .A(n_227), .Y(n_867) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_228), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1571 ( .A1(n_229), .A2(n_1572), .B1(n_1577), .B2(n_1634), .Y(n_1571) );
OAI22xp5_ASAP7_75t_L g1579 ( .A1(n_229), .A2(n_1580), .B1(n_1632), .B2(n_1633), .Y(n_1579) );
INVxp67_ASAP7_75t_SL g1633 ( .A(n_229), .Y(n_1633) );
INVx1_ASAP7_75t_L g1588 ( .A(n_230), .Y(n_1588) );
INVx1_ASAP7_75t_L g908 ( .A(n_231), .Y(n_908) );
INVx1_ASAP7_75t_L g1601 ( .A(n_234), .Y(n_1601) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_237), .Y(n_1151) );
INVx1_ASAP7_75t_L g1115 ( .A(n_238), .Y(n_1115) );
OAI211xp5_ASAP7_75t_L g1089 ( .A1(n_241), .A2(n_1029), .B(n_1090), .C(n_1092), .Y(n_1089) );
INVx1_ASAP7_75t_L g1133 ( .A(n_241), .Y(n_1133) );
INVx1_ASAP7_75t_L g1157 ( .A(n_242), .Y(n_1157) );
HB1xp67_ASAP7_75t_L g1173 ( .A(n_242), .Y(n_1173) );
INVx1_ASAP7_75t_L g1188 ( .A(n_243), .Y(n_1188) );
INVx1_ASAP7_75t_L g722 ( .A(n_244), .Y(n_722) );
INVx1_ASAP7_75t_L g1249 ( .A(n_245), .Y(n_1249) );
INVx1_ASAP7_75t_L g1016 ( .A(n_246), .Y(n_1016) );
AOI21xp33_ASAP7_75t_L g1146 ( .A1(n_247), .A2(n_361), .B(n_560), .Y(n_1146) );
INVx1_ASAP7_75t_L g1290 ( .A(n_248), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_248), .B(n_1288), .Y(n_1295) );
OAI221xp5_ASAP7_75t_L g588 ( .A1(n_249), .A2(n_589), .B1(n_592), .B2(n_600), .C(n_607), .Y(n_588) );
INVx1_ASAP7_75t_L g638 ( .A(n_251), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_252), .Y(n_820) );
OAI211xp5_ASAP7_75t_L g1076 ( .A1(n_254), .A2(n_862), .B(n_1077), .C(n_1078), .Y(n_1076) );
INVx1_ASAP7_75t_L g1112 ( .A(n_254), .Y(n_1112) );
INVx1_ASAP7_75t_L g1184 ( .A(n_255), .Y(n_1184) );
INVxp67_ASAP7_75t_SL g1626 ( .A(n_256), .Y(n_1626) );
INVx2_ASAP7_75t_L g300 ( .A(n_257), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_258), .B(n_727), .Y(n_726) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_260), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g343 ( .A1(n_261), .A2(n_263), .B1(n_344), .B2(n_353), .C(n_357), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_261), .A2(n_263), .B1(n_427), .B2(n_432), .Y(n_426) );
INVx1_ASAP7_75t_L g715 ( .A(n_262), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_264), .A2(n_265), .B1(n_838), .B2(n_840), .Y(n_839) );
OAI221xp5_ASAP7_75t_L g860 ( .A1(n_264), .A2(n_589), .B1(n_607), .B2(n_861), .C(n_870), .Y(n_860) );
OAI211xp5_ASAP7_75t_SL g848 ( .A1(n_265), .A2(n_563), .B(n_849), .C(n_859), .Y(n_848) );
INVx1_ASAP7_75t_L g1238 ( .A(n_266), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_266), .A2(n_269), .B1(n_990), .B2(n_1263), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g1532 ( .A(n_268), .Y(n_1532) );
INVx1_ASAP7_75t_L g1235 ( .A(n_269), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_270), .Y(n_1102) );
INVx1_ASAP7_75t_L g377 ( .A(n_272), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_274), .Y(n_381) );
BUFx3_ASAP7_75t_L g414 ( .A(n_275), .Y(n_414) );
INVx1_ASAP7_75t_L g443 ( .A(n_275), .Y(n_443) );
BUFx3_ASAP7_75t_L g416 ( .A(n_276), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_276), .Y(n_423) );
OAI221xp5_ASAP7_75t_L g653 ( .A1(n_278), .A2(n_563), .B1(n_654), .B2(n_658), .C(n_666), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_279), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g1094 ( .A(n_280), .Y(n_1094) );
INVx1_ASAP7_75t_L g771 ( .A(n_281), .Y(n_771) );
OAI211xp5_ASAP7_75t_L g790 ( .A1(n_281), .A2(n_563), .B(n_791), .C(n_798), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_304), .B(n_1277), .Y(n_282) );
BUFx12f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
AND2x4_ASAP7_75t_L g1576 ( .A(n_286), .B(n_292), .Y(n_1576) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g1570 ( .A(n_287), .Y(n_1570) );
NAND2xp5_ASAP7_75t_L g1637 ( .A(n_287), .B(n_289), .Y(n_1637) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_289), .B(n_1570), .Y(n_1569) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x6_ASAP7_75t_L g941 ( .A(n_294), .B(n_405), .Y(n_941) );
OR2x2_ASAP7_75t_L g1069 ( .A(n_294), .B(n_405), .Y(n_1069) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g599 ( .A(n_295), .B(n_303), .Y(n_599) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g361 ( .A(n_296), .B(n_362), .Y(n_361) );
INVx8_ASAP7_75t_L g937 ( .A(n_297), .Y(n_937) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
INVx2_ASAP7_75t_SL g367 ( .A(n_298), .Y(n_367) );
OR2x2_ASAP7_75t_L g402 ( .A(n_298), .B(n_351), .Y(n_402) );
INVx1_ASAP7_75t_L g596 ( .A(n_298), .Y(n_596) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_298), .Y(n_650) );
OR2x6_ASAP7_75t_L g940 ( .A(n_298), .B(n_931), .Y(n_940) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x4_ASAP7_75t_L g319 ( .A(n_300), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g329 ( .A(n_300), .Y(n_329) );
AND2x2_ASAP7_75t_L g335 ( .A(n_300), .B(n_301), .Y(n_335) );
INVx2_ASAP7_75t_L g340 ( .A(n_300), .Y(n_340) );
INVx1_ASAP7_75t_L g374 ( .A(n_300), .Y(n_374) );
INVx2_ASAP7_75t_L g320 ( .A(n_301), .Y(n_320) );
INVx1_ASAP7_75t_L g342 ( .A(n_301), .Y(n_342) );
INVx1_ASAP7_75t_L g349 ( .A(n_301), .Y(n_349) );
INVx1_ASAP7_75t_L g373 ( .A(n_301), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_301), .B(n_340), .Y(n_380) );
AND2x4_ASAP7_75t_L g926 ( .A(n_302), .B(n_349), .Y(n_926) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g927 ( .A(n_303), .B(n_928), .Y(n_927) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_303), .B(n_928), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_811), .B2(n_1276), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
XNOR2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_618), .Y(n_306) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_487), .B1(n_488), .B2(n_617), .Y(n_307) );
INVx3_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_399), .Y(n_310) );
NOR3xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_343), .C(n_359), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_330), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_325), .B2(n_326), .Y(n_313) );
BUFx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_321), .Y(n_316) );
INVx1_ASAP7_75t_L g1549 ( .A(n_317), .Y(n_1549) );
INVx3_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_318), .Y(n_664) );
INVx3_ASAP7_75t_L g994 ( .A(n_318), .Y(n_994) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_319), .Y(n_383) );
INVx1_ASAP7_75t_L g576 ( .A(n_319), .Y(n_576) );
INVx1_ASAP7_75t_L g875 ( .A(n_319), .Y(n_875) );
AND2x4_ASAP7_75t_L g328 ( .A(n_320), .B(n_329), .Y(n_328) );
AND2x6_ASAP7_75t_L g326 ( .A(n_321), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g332 ( .A(n_321), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g337 ( .A(n_321), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g395 ( .A(n_322), .Y(n_395) );
OR2x2_ASAP7_75t_L g538 ( .A(n_322), .B(n_425), .Y(n_538) );
INVx2_ASAP7_75t_L g566 ( .A(n_323), .Y(n_566) );
AND2x4_ASAP7_75t_L g590 ( .A(n_323), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g611 ( .A(n_323), .B(n_339), .Y(n_611) );
INVx1_ASAP7_75t_L g362 ( .A(n_324), .Y(n_362) );
INVx1_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g444 ( .A1(n_325), .A2(n_331), .B1(n_445), .B2(n_450), .C(n_452), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_327), .B(n_350), .Y(n_358) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx3_ASAP7_75t_L g567 ( .A(n_328), .Y(n_567) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_328), .Y(n_580) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_328), .Y(n_699) );
AND2x4_ASAP7_75t_L g921 ( .A(n_328), .B(n_922), .Y(n_921) );
BUFx2_ASAP7_75t_L g1253 ( .A(n_328), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B1(n_336), .B2(n_337), .Y(n_330) );
INVx1_ASAP7_75t_L g579 ( .A(n_333), .Y(n_579) );
BUFx2_ASAP7_75t_L g709 ( .A(n_333), .Y(n_709) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_SL g560 ( .A(n_334), .Y(n_560) );
INVx2_ASAP7_75t_L g796 ( .A(n_334), .Y(n_796) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_335), .Y(n_591) );
INVx2_ASAP7_75t_SL g951 ( .A(n_338), .Y(n_951) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx2_ASAP7_75t_L g694 ( .A(n_339), .Y(n_694) );
BUFx2_ASAP7_75t_L g712 ( .A(n_339), .Y(n_712) );
AND2x4_ASAP7_75t_L g930 ( .A(n_339), .B(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g991 ( .A(n_339), .Y(n_991) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g356 ( .A(n_340), .Y(n_356) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2x1_ASAP7_75t_SL g346 ( .A(n_347), .B(n_350), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g702 ( .A(n_347), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_349), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g1156 ( .A1(n_349), .A2(n_355), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_350), .B(n_355), .Y(n_354) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g559 ( .A(n_352), .Y(n_559) );
BUFx4f_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x6_ASAP7_75t_L g587 ( .A(n_356), .B(n_558), .Y(n_587) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI33xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_364), .A3(n_376), .B1(n_384), .B2(n_388), .B3(n_392), .Y(n_359) );
OAI33xp33_ASAP7_75t_L g1118 ( .A1(n_360), .A2(n_392), .A3(n_1119), .B1(n_1122), .B2(n_1125), .B3(n_1129), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g1607 ( .A1(n_360), .A2(n_1608), .B1(n_1615), .B2(n_1616), .Y(n_1607) );
OR2x6_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g931 ( .A(n_362), .Y(n_931) );
BUFx2_ASAP7_75t_L g486 ( .A(n_363), .Y(n_486) );
INVx2_ASAP7_75t_L g508 ( .A(n_363), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B1(n_369), .B2(n_375), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_365), .A2(n_389), .B1(n_390), .B2(n_391), .Y(n_388) );
BUFx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g390 ( .A(n_370), .Y(n_390) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g593 ( .A(n_371), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g654 ( .A1(n_371), .A2(n_635), .B1(n_650), .B2(n_655), .C(n_656), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g1144 ( .A1(n_371), .A2(n_1145), .B(n_1146), .Y(n_1144) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g608 ( .A(n_372), .Y(n_608) );
BUFx2_ASAP7_75t_L g863 ( .A(n_372), .Y(n_863) );
INVx2_ASAP7_75t_L g1042 ( .A(n_372), .Y(n_1042) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_373), .B(n_374), .Y(n_648) );
INVx1_ASAP7_75t_L g928 ( .A(n_374), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B1(n_381), .B2(n_382), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_378), .A2(n_385), .B1(n_386), .B2(n_387), .Y(n_384) );
BUFx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_379), .B(n_1074), .Y(n_1073) );
INVx2_ASAP7_75t_L g1124 ( .A(n_379), .Y(n_1124) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g571 ( .A(n_380), .Y(n_571) );
INVx1_ASAP7_75t_L g661 ( .A(n_380), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g791 ( .A1(n_382), .A2(n_792), .B1(n_793), .B2(n_794), .C(n_795), .Y(n_791) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_SL g386 ( .A(n_383), .Y(n_386) );
BUFx3_ASAP7_75t_L g606 ( .A(n_383), .Y(n_606) );
INVx2_ASAP7_75t_SL g644 ( .A(n_383), .Y(n_644) );
INVx4_ASAP7_75t_L g714 ( .A(n_383), .Y(n_714) );
INVx2_ASAP7_75t_SL g1557 ( .A(n_383), .Y(n_1557) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_385), .A2(n_420), .B(n_426), .C(n_437), .Y(n_419) );
INVx1_ASAP7_75t_L g695 ( .A(n_386), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_387), .A2(n_389), .B1(n_479), .B2(n_481), .Y(n_478) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_391), .A2(n_457), .B1(n_462), .B2(n_467), .C(n_474), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g1598 ( .A(n_392), .B(n_1599), .C(n_1604), .Y(n_1598) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI33xp33_ASAP7_75t_L g943 ( .A1(n_393), .A2(n_944), .A3(n_946), .B1(n_948), .B2(n_949), .B3(n_952), .Y(n_943) );
AOI33xp33_ASAP7_75t_L g1048 ( .A1(n_393), .A2(n_1049), .A3(n_1050), .B1(n_1051), .B2(n_1052), .B3(n_1053), .Y(n_1048) );
AOI33xp33_ASAP7_75t_L g1195 ( .A1(n_393), .A2(n_1049), .A3(n_1196), .B1(n_1198), .B2(n_1200), .B3(n_1202), .Y(n_1195) );
INVx6_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx5_ASAP7_75t_L g997 ( .A(n_394), .Y(n_997) );
OR2x6_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_395), .B(n_407), .Y(n_500) );
INVx2_ASAP7_75t_L g582 ( .A(n_396), .Y(n_582) );
BUFx2_ASAP7_75t_L g797 ( .A(n_396), .Y(n_797) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g923 ( .A(n_397), .Y(n_923) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_417), .B(n_418), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OR2x6_ASAP7_75t_L g553 ( .A(n_404), .B(n_554), .Y(n_553) );
AOI222xp33_ASAP7_75t_L g1174 ( .A1(n_404), .A2(n_545), .B1(n_548), .B2(n_1148), .C1(n_1154), .C2(n_1175), .Y(n_1174) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AND2x4_ASAP7_75t_L g529 ( .A(n_405), .B(n_454), .Y(n_529) );
AND2x4_ASAP7_75t_L g779 ( .A(n_405), .B(n_454), .Y(n_779) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_412), .Y(n_406) );
AND2x4_ASAP7_75t_L g428 ( .A(n_407), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_407), .Y(n_433) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g454 ( .A(n_410), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g466 ( .A(n_411), .B(n_455), .Y(n_466) );
INVx1_ASAP7_75t_L g887 ( .A(n_411), .Y(n_887) );
INVx1_ASAP7_75t_L g892 ( .A(n_411), .Y(n_892) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_411), .Y(n_897) );
INVx6_ASAP7_75t_L g471 ( .A(n_412), .Y(n_471) );
INVx2_ASAP7_75t_L g517 ( .A(n_412), .Y(n_517) );
BUFx2_ASAP7_75t_L g837 ( .A(n_412), .Y(n_837) );
AND2x4_ASAP7_75t_L g895 ( .A(n_412), .B(n_896), .Y(n_895) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g436 ( .A(n_413), .Y(n_436) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g422 ( .A(n_414), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g461 ( .A(n_414), .B(n_416), .Y(n_461) );
INVx1_ASAP7_75t_L g431 ( .A(n_415), .Y(n_431) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g442 ( .A(n_416), .B(n_443), .Y(n_442) );
AOI31xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_456), .A3(n_478), .B(n_484), .Y(n_418) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
BUFx3_ASAP7_75t_L g438 ( .A(n_421), .Y(n_438) );
INVx2_ASAP7_75t_SL g511 ( .A(n_421), .Y(n_511) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_422), .Y(n_525) );
INVx2_ASAP7_75t_SL g550 ( .A(n_422), .Y(n_550) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_422), .Y(n_684) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_422), .Y(n_738) );
BUFx3_ASAP7_75t_L g757 ( .A(n_422), .Y(n_757) );
BUFx2_ASAP7_75t_L g832 ( .A(n_422), .Y(n_832) );
AND2x6_ASAP7_75t_L g890 ( .A(n_422), .B(n_891), .Y(n_890) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_422), .Y(n_1207) );
INVx1_ASAP7_75t_L g449 ( .A(n_423), .Y(n_449) );
AND2x4_ASAP7_75t_L g459 ( .A(n_424), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g480 ( .A(n_425), .B(n_451), .Y(n_480) );
OR2x2_ASAP7_75t_L g482 ( .A(n_425), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g498 ( .A(n_430), .Y(n_498) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g907 ( .A(n_431), .Y(n_907) );
OR2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_SL g475 ( .A(n_433), .Y(n_475) );
OR2x6_ASAP7_75t_L g503 ( .A(n_434), .B(n_500), .Y(n_503) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g1629 ( .A(n_435), .Y(n_1629) );
BUFx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x6_ASAP7_75t_L g909 ( .A(n_436), .B(n_892), .Y(n_909) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g679 ( .A(n_441), .Y(n_679) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_441), .Y(n_739) );
INVx1_ASAP7_75t_L g759 ( .A(n_441), .Y(n_759) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g473 ( .A(n_442), .Y(n_473) );
INVx2_ASAP7_75t_L g483 ( .A(n_442), .Y(n_483) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_442), .Y(n_514) );
INVx1_ASAP7_75t_L g527 ( .A(n_442), .Y(n_527) );
INVx1_ASAP7_75t_L g448 ( .A(n_443), .Y(n_448) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g770 ( .A(n_446), .Y(n_770) );
BUFx4f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g542 ( .A(n_447), .Y(n_542) );
BUFx2_ASAP7_75t_L g766 ( .A(n_447), .Y(n_766) );
INVx1_ASAP7_75t_L g1109 ( .A(n_447), .Y(n_1109) );
INVx1_ASAP7_75t_L g1585 ( .A(n_447), .Y(n_1585) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
OR2x2_ASAP7_75t_L g451 ( .A(n_448), .B(n_449), .Y(n_451) );
BUFx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g763 ( .A(n_451), .Y(n_763) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_451), .B(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1631 ( .A(n_451), .Y(n_1631) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g915 ( .A(n_455), .Y(n_915) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g464 ( .A(n_460), .Y(n_464) );
INVx2_ASAP7_75t_SL g519 ( .A(n_460), .Y(n_519) );
BUFx3_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_460), .Y(n_531) );
BUFx4f_ASAP7_75t_L g675 ( .A(n_460), .Y(n_675) );
INVx1_ASAP7_75t_L g1212 ( .A(n_460), .Y(n_1212) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_461), .Y(n_477) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g507 ( .A(n_466), .Y(n_507) );
INVx1_ASAP7_75t_L g987 ( .A(n_466), .Y(n_987) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g981 ( .A(n_470), .Y(n_981) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g674 ( .A(n_471), .Y(n_674) );
INVx1_ASAP7_75t_L g743 ( .A(n_471), .Y(n_743) );
BUFx6f_ASAP7_75t_L g841 ( .A(n_471), .Y(n_841) );
INVx2_ASAP7_75t_L g888 ( .A(n_471), .Y(n_888) );
HB1xp67_ASAP7_75t_L g1166 ( .A(n_471), .Y(n_1166) );
INVx1_ASAP7_75t_L g1270 ( .A(n_471), .Y(n_1270) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x6_ASAP7_75t_L g537 ( .A(n_473), .B(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g803 ( .A(n_473), .B(n_538), .Y(n_803) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
BUFx6f_ASAP7_75t_L g1059 ( .A(n_476), .Y(n_1059) );
OAI21xp33_ASAP7_75t_L g1241 ( .A1(n_476), .A2(n_912), .B(n_1242), .Y(n_1241) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g632 ( .A(n_477), .Y(n_632) );
AND2x4_ASAP7_75t_L g911 ( .A(n_477), .B(n_912), .Y(n_911) );
BUFx6f_ASAP7_75t_L g969 ( .A(n_477), .Y(n_969) );
INVx2_ASAP7_75t_L g983 ( .A(n_477), .Y(n_983) );
INVx6_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g835 ( .A(n_483), .Y(n_835) );
INVx1_ASAP7_75t_L g1104 ( .A(n_483), .Y(n_1104) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g616 ( .A(n_486), .Y(n_616) );
AND2x4_ASAP7_75t_L g914 ( .A(n_486), .B(n_915), .Y(n_914) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_486), .B(n_915), .Y(n_1037) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND3x1_ASAP7_75t_L g491 ( .A(n_492), .B(n_551), .C(n_561), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_533), .Y(n_492) );
NAND3xp33_ASAP7_75t_SL g493 ( .A(n_494), .B(n_504), .C(n_530), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_501), .B2(n_502), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_495), .A2(n_501), .B1(n_584), .B2(n_586), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_496), .A2(n_502), .B1(n_628), .B2(n_629), .C(n_630), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_496), .A2(n_502), .B1(n_827), .B2(n_828), .Y(n_826) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g732 ( .A(n_497), .Y(n_732) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g1628 ( .A(n_498), .Y(n_1628) );
INVx2_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g532 ( .A(n_500), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g731 ( .A1(n_502), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AOI33xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_509), .A3(n_515), .B1(n_520), .B2(n_523), .B3(n_528), .Y(n_504) );
AOI33xp33_ASAP7_75t_L g735 ( .A1(n_505), .A2(n_528), .A3(n_736), .B1(n_740), .B2(n_744), .B3(n_746), .Y(n_735) );
AOI33xp33_ASAP7_75t_L g956 ( .A1(n_505), .A2(n_528), .A3(n_957), .B1(n_959), .B2(n_960), .B3(n_961), .Y(n_956) );
AOI33xp33_ASAP7_75t_L g1054 ( .A1(n_505), .A2(n_529), .A3(n_1055), .B1(n_1056), .B2(n_1057), .B3(n_1060), .Y(n_1054) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_506), .Y(n_671) );
INVx2_ASAP7_75t_L g830 ( .A(n_506), .Y(n_830) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
OR2x2_ASAP7_75t_L g754 ( .A(n_507), .B(n_508), .Y(n_754) );
INVx2_ASAP7_75t_L g555 ( .A(n_508), .Y(n_555) );
BUFx2_ASAP7_75t_L g718 ( .A(n_508), .Y(n_718) );
AND2x4_ASAP7_75t_L g945 ( .A(n_508), .B(n_599), .Y(n_945) );
OR2x2_ASAP7_75t_L g986 ( .A(n_508), .B(n_987), .Y(n_986) );
AND2x4_ASAP7_75t_L g1049 ( .A(n_508), .B(n_599), .Y(n_1049) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g677 ( .A(n_511), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g1167 ( .A1(n_511), .A2(n_527), .B1(n_1141), .B2(n_1143), .Y(n_1167) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g685 ( .A(n_513), .Y(n_685) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_514), .Y(n_776) );
AND2x6_ASAP7_75t_L g899 ( .A(n_514), .B(n_886), .Y(n_899) );
INVx1_ASAP7_75t_L g1116 ( .A(n_514), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1208 ( .A(n_514), .Y(n_1208) );
BUFx6f_ASAP7_75t_L g1214 ( .A(n_514), .Y(n_1214) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_SL g521 ( .A(n_517), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_518), .B(n_1025), .Y(n_1024) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g838 ( .A(n_519), .Y(n_838) );
AND2x2_ASAP7_75t_L g545 ( .A(n_521), .B(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g808 ( .A(n_525), .Y(n_808) );
BUFx4f_ASAP7_75t_L g843 ( .A(n_525), .Y(n_843) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g747 ( .A(n_527), .Y(n_747) );
OAI22xp33_ASAP7_75t_L g1526 ( .A1(n_527), .A2(n_1527), .B1(n_1528), .B2(n_1529), .Y(n_1526) );
BUFx4f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx4f_ASAP7_75t_L g686 ( .A(n_529), .Y(n_686) );
INVx4_ASAP7_75t_L g1117 ( .A(n_529), .Y(n_1117) );
AOI221xp5_ASAP7_75t_L g1163 ( .A1(n_529), .A2(n_830), .B1(n_1164), .B2(n_1168), .C(n_1172), .Y(n_1163) );
INVx1_ASAP7_75t_L g730 ( .A(n_530), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_531), .Y(n_745) );
AND2x2_ASAP7_75t_L g630 ( .A(n_532), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_543), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B1(n_539), .B2(n_540), .Y(n_534) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_535), .A2(n_547), .B1(n_569), .B2(n_572), .C(n_577), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_536), .A2(n_540), .B1(n_724), .B2(n_725), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_536), .A2(n_540), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_536), .A2(n_540), .B1(n_1149), .B2(n_1151), .Y(n_1176) );
CKINVDCx6p67_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
OR2x6_ASAP7_75t_L g541 ( .A(n_538), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g546 ( .A(n_538), .Y(n_546) );
OR2x2_ASAP7_75t_L g805 ( .A(n_538), .B(n_806), .Y(n_805) );
OR2x2_ASAP7_75t_L g807 ( .A(n_538), .B(n_808), .Y(n_807) );
CKINVDCx6p67_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
BUFx3_ASAP7_75t_L g1111 ( .A(n_542), .Y(n_1111) );
INVx1_ASAP7_75t_L g1619 ( .A(n_542), .Y(n_1619) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B1(n_547), .B2(n_548), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_545), .A2(n_548), .B1(n_634), .B2(n_635), .C(n_636), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_545), .A2(n_548), .B1(n_721), .B2(n_722), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_545), .A2(n_548), .B1(n_823), .B2(n_824), .Y(n_822) );
AND2x2_ASAP7_75t_L g548 ( .A(n_546), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g1007 ( .A(n_550), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_550), .A2(n_1114), .B1(n_1115), .B2(n_1116), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_553), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g727 ( .A(n_553), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_553), .B(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_553), .B(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_553), .B(n_1544), .Y(n_1543) );
NOR2xp67_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g1162 ( .A(n_555), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
AND2x2_ASAP7_75t_L g584 ( .A(n_557), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g667 ( .A(n_557), .B(n_585), .Y(n_667) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OR2x2_ASAP7_75t_L g607 ( .A(n_558), .B(n_608), .Y(n_607) );
OR2x6_ASAP7_75t_L g652 ( .A(n_558), .B(n_608), .Y(n_652) );
INVx1_ASAP7_75t_L g703 ( .A(n_558), .Y(n_703) );
INVx1_ASAP7_75t_L g1159 ( .A(n_558), .Y(n_1159) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
BUFx2_ASAP7_75t_L g996 ( .A(n_560), .Y(n_996) );
OAI31xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_588), .A3(n_609), .B(n_615), .Y(n_561) );
INVx8_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_564), .A2(n_693), .B1(n_696), .B2(n_700), .C(n_701), .Y(n_692) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
AND2x4_ASAP7_75t_L g613 ( .A(n_565), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g856 ( .A(n_567), .Y(n_856) );
BUFx6f_ASAP7_75t_L g1614 ( .A(n_567), .Y(n_1614) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g603 ( .A(n_571), .Y(n_603) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g614 ( .A(n_576), .Y(n_614) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_SL g919 ( .A(n_580), .Y(n_919) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_580), .Y(n_1002) );
BUFx2_ASAP7_75t_L g1203 ( .A(n_580), .Y(n_1203) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g657 ( .A(n_582), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_584), .A2(n_586), .B1(n_799), .B2(n_800), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_584), .A2(n_586), .B1(n_1561), .B2(n_1562), .Y(n_1560) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_586), .A2(n_628), .B1(n_629), .B2(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_586), .A2(n_667), .B1(n_827), .B2(n_828), .Y(n_859) );
CKINVDCx11_ASAP7_75t_R g586 ( .A(n_587), .Y(n_586) );
CKINVDCx6p67_ASAP7_75t_R g589 ( .A(n_590), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_590), .A2(n_708), .B1(n_711), .B2(n_715), .C(n_716), .Y(n_707) );
INVx3_ASAP7_75t_L g858 ( .A(n_591), .Y(n_858) );
BUFx6f_ASAP7_75t_L g955 ( .A(n_591), .Y(n_955) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_595), .B2(n_597), .C(n_598), .Y(n_592) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g789 ( .A(n_596), .Y(n_789) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_598), .A2(n_647), .B1(n_649), .B2(n_650), .C(n_651), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g788 ( .A1(n_598), .A2(n_647), .B1(n_764), .B2(n_767), .C(n_789), .Y(n_788) );
BUFx2_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g869 ( .A(n_599), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_600) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_SL g642 ( .A(n_603), .Y(n_642) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g1121 ( .A(n_608), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_608), .B(n_1156), .Y(n_1155) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_611), .A2(n_613), .B1(n_705), .B2(n_706), .Y(n_704) );
INVx3_ASAP7_75t_L g785 ( .A(n_611), .Y(n_785) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx3_ASAP7_75t_L g669 ( .A(n_613), .Y(n_669) );
INVx1_ASAP7_75t_L g853 ( .A(n_614), .Y(n_853) );
OAI31xp33_ASAP7_75t_L g639 ( .A1(n_615), .A2(n_640), .A3(n_653), .B(n_668), .Y(n_639) );
OAI31xp33_ASAP7_75t_L g783 ( .A1(n_615), .A2(n_784), .A3(n_786), .B(n_790), .Y(n_783) );
OAI31xp33_ASAP7_75t_L g1545 ( .A1(n_615), .A2(n_1546), .A3(n_1547), .B(n_1554), .Y(n_1545) );
BUFx8_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_748), .B1(n_749), .B2(n_809), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_622), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_687), .B2(n_688), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND4xp75_ASAP7_75t_SL g625 ( .A(n_626), .B(n_637), .C(n_639), .D(n_670), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_633), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_630), .B(n_753), .C(n_780), .Y(n_752) );
NOR3xp33_ASAP7_75t_L g1524 ( .A(n_630), .B(n_1525), .C(n_1542), .Y(n_1524) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_634), .A2(n_659), .B1(n_662), .B2(n_665), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_644), .B2(n_645), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_642), .A2(n_714), .B1(n_758), .B2(n_760), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g1125 ( .A1(n_642), .A2(n_1094), .B1(n_1126), .B2(n_1128), .Y(n_1125) );
INVx2_ASAP7_75t_L g1132 ( .A(n_647), .Y(n_1132) );
BUFx3_ASAP7_75t_L g1551 ( .A(n_647), .Y(n_1551) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g866 ( .A(n_650), .Y(n_866) );
OAI22xp33_ASAP7_75t_L g1119 ( .A1(n_650), .A2(n_1106), .B1(n_1107), .B2(n_1120), .Y(n_1119) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_650), .A2(n_1130), .B1(n_1131), .B2(n_1133), .Y(n_1129) );
OAI22xp33_ASAP7_75t_SL g1604 ( .A1(n_650), .A2(n_862), .B1(n_1605), .B2(n_1606), .Y(n_1604) );
INVx2_ASAP7_75t_L g716 ( .A(n_652), .Y(n_716) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g850 ( .A(n_660), .Y(n_850) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g792 ( .A(n_661), .Y(n_792) );
INVx2_ASAP7_75t_L g872 ( .A(n_661), .Y(n_872) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx3_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_SL g1127 ( .A(n_664), .Y(n_1127) );
INVx2_ASAP7_75t_L g1263 ( .A(n_664), .Y(n_1263) );
INVx2_ASAP7_75t_L g1603 ( .A(n_664), .Y(n_1603) );
INVx2_ASAP7_75t_L g1611 ( .A(n_664), .Y(n_1611) );
AOI33xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .A3(n_676), .B1(n_680), .B2(n_681), .B3(n_686), .Y(n_670) );
BUFx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_674), .Y(n_1058) );
AOI222xp33_ASAP7_75t_L g900 ( .A1(n_675), .A2(n_901), .B1(n_902), .B2(n_903), .C1(n_908), .C2(n_909), .Y(n_900) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g1101 ( .A(n_683), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1169 ( .A1(n_683), .A2(n_834), .B1(n_1170), .B2(n_1171), .Y(n_1169) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g773 ( .A(n_684), .Y(n_773) );
AOI322xp5_ASAP7_75t_L g1092 ( .A1(n_684), .A2(n_909), .A3(n_1081), .B1(n_1085), .B2(n_1093), .C1(n_1094), .C2(n_1095), .Y(n_1092) );
INVx2_ASAP7_75t_SL g1527 ( .A(n_684), .Y(n_1527) );
CKINVDCx5p33_ASAP7_75t_R g1615 ( .A(n_686), .Y(n_1615) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
XNOR2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NOR4xp75_ASAP7_75t_L g690 ( .A(n_691), .B(n_719), .C(n_726), .D(n_728), .Y(n_690) );
AOI31xp33_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_704), .A3(n_707), .B(n_717), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g1009 ( .A1(n_697), .A2(n_921), .B(n_1010), .C(n_1011), .Y(n_1009) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g710 ( .A(n_698), .Y(n_710) );
INVx2_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
BUFx6f_ASAP7_75t_L g1197 ( .A(n_699), .Y(n_1197) );
AOI222xp33_ASAP7_75t_L g1189 ( .A1(n_710), .A2(n_1082), .B1(n_1190), .B2(n_1191), .C1(n_1192), .C2(n_1193), .Y(n_1189) );
INVx2_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g877 ( .A(n_717), .Y(n_877) );
CKINVDCx8_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_723), .Y(n_719) );
NAND3xp33_ASAP7_75t_SL g728 ( .A(n_729), .B(n_731), .C(n_735), .Y(n_728) );
NAND3xp33_ASAP7_75t_L g825 ( .A(n_729), .B(n_826), .C(n_829), .Y(n_825) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
BUFx3_ASAP7_75t_L g958 ( .A(n_738), .Y(n_958) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AND4x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_781), .C(n_783), .D(n_801), .Y(n_751) );
OAI33xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .A3(n_761), .B1(n_768), .B2(n_772), .B3(n_778), .Y(n_753) );
OAI33xp33_ASAP7_75t_L g1097 ( .A1(n_754), .A2(n_1098), .A3(n_1105), .B1(n_1110), .B2(n_1113), .B3(n_1117), .Y(n_1097) );
INVx1_ASAP7_75t_SL g1205 ( .A(n_754), .Y(n_1205) );
OAI33xp33_ASAP7_75t_L g1525 ( .A1(n_754), .A2(n_778), .A3(n_1526), .B1(n_1530), .B2(n_1533), .B3(n_1539), .Y(n_1525) );
OAI22xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_755) );
INVx2_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_759), .A2(n_773), .B1(n_1540), .B2(n_1541), .Y(n_1539) );
OAI22xp33_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_764), .B1(n_765), .B2(n_767), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g768 ( .A1(n_762), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
OAI22xp33_ASAP7_75t_SL g1105 ( .A1(n_762), .A2(n_1106), .B1(n_1107), .B2(n_1108), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1110 ( .A1(n_762), .A2(n_1071), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g1530 ( .A1(n_762), .A2(n_765), .B1(n_1531), .B2(n_1532), .Y(n_1530) );
OAI221xp5_ASAP7_75t_L g1616 ( .A1(n_762), .A2(n_1617), .B1(n_1618), .B2(n_1620), .C(n_1621), .Y(n_1616) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g806 ( .A(n_763), .Y(n_806) );
INVx2_ASAP7_75t_L g1534 ( .A(n_763), .Y(n_1534) );
INVx2_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B1(n_775), .B2(n_777), .Y(n_772) );
INVx2_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AOI33xp33_ASAP7_75t_L g829 ( .A1(n_779), .A2(n_830), .A3(n_831), .B1(n_836), .B2(n_839), .B3(n_842), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g1003 ( .A(n_779), .B(n_1004), .C(n_1006), .Y(n_1003) );
AOI33xp33_ASAP7_75t_L g1204 ( .A1(n_779), .A2(n_1205), .A3(n_1206), .B1(n_1209), .B2(n_1210), .B3(n_1213), .Y(n_1204) );
NAND3xp33_ASAP7_75t_L g1268 ( .A(n_779), .B(n_1269), .C(n_1271), .Y(n_1268) );
OAI221xp5_ASAP7_75t_L g1555 ( .A1(n_792), .A2(n_1556), .B1(n_1557), .B2(n_1558), .C(n_1559), .Y(n_1555) );
BUFx3_ASAP7_75t_L g947 ( .A(n_796), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_804), .Y(n_801) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g1276 ( .A(n_811), .Y(n_1276) );
AO22x2_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_1063), .B1(n_1064), .B2(n_1275), .Y(n_811) );
INVx1_ASAP7_75t_L g1275 ( .A(n_812), .Y(n_1275) );
XOR2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_878), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_845), .C(n_847), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_825), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_822), .Y(n_818) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_820), .A2(n_824), .B1(n_850), .B2(n_851), .C(n_854), .Y(n_849) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g844 ( .A(n_834), .Y(n_844) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
HB1xp67_ASAP7_75t_L g1624 ( .A(n_837), .Y(n_1624) );
INVx4_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g1005 ( .A(n_841), .Y(n_1005) );
OAI31xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_860), .A3(n_876), .B(n_877), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g1599 ( .A1(n_850), .A2(n_1600), .B1(n_1601), .B2(n_1602), .Y(n_1599) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g1000 ( .A(n_853), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_853), .A2(n_1099), .B1(n_1102), .B2(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g1079 ( .A(n_858), .Y(n_1079) );
INVx2_ASAP7_75t_SL g1553 ( .A(n_858), .Y(n_1553) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_864), .B1(n_865), .B2(n_867), .C(n_868), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_872), .A2(n_1141), .B1(n_1142), .B2(n_1143), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_872), .A2(n_993), .B1(n_1148), .B2(n_1149), .Y(n_1147) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g934 ( .A(n_875), .Y(n_934) );
XNOR2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_962), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
AOI211x1_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_913), .B(n_916), .C(n_942), .Y(n_881) );
NAND4xp25_ASAP7_75t_SL g882 ( .A(n_883), .B(n_893), .C(n_900), .D(n_910), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_889), .B2(n_890), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_885), .A2(n_895), .B1(n_973), .B2(n_974), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_885), .A2(n_899), .B1(n_1234), .B2(n_1235), .Y(n_1233) );
AND2x4_ASAP7_75t_L g885 ( .A(n_886), .B(n_888), .Y(n_885) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_886), .B(n_888), .Y(n_1224) );
INVx1_ASAP7_75t_SL g886 ( .A(n_887), .Y(n_886) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_887), .B(n_1221), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_890), .A2(n_899), .B1(n_976), .B2(n_977), .Y(n_975) );
CKINVDCx6p67_ASAP7_75t_R g1031 ( .A(n_890), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_890), .A2(n_899), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
AOI221xp5_ASAP7_75t_L g1236 ( .A1(n_890), .A2(n_895), .B1(n_1237), .B2(n_1238), .C(n_1239), .Y(n_1236) );
INVx1_ASAP7_75t_L g912 ( .A(n_891), .Y(n_912) );
INVx1_ASAP7_75t_L g1035 ( .A(n_891), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_891), .B(n_969), .Y(n_1091) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_895), .B1(n_898), .B2(n_899), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_894), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_936) );
INVx4_ASAP7_75t_L g1036 ( .A(n_895), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_895), .A2(n_1188), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
AND2x4_ASAP7_75t_L g905 ( .A(n_896), .B(n_906), .Y(n_905) );
AND2x2_ASAP7_75t_SL g1095 ( .A(n_896), .B(n_906), .Y(n_1095) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx4_ASAP7_75t_L g1032 ( .A(n_899), .Y(n_1032) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_905), .A2(n_909), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1586 ( .A1(n_905), .A2(n_909), .B1(n_1587), .B2(n_1588), .Y(n_1586) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g1221 ( .A(n_907), .Y(n_1221) );
INVx3_ASAP7_75t_L g971 ( .A(n_909), .Y(n_971) );
INVx5_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
AOI211xp5_ASAP7_75t_L g966 ( .A1(n_911), .A2(n_967), .B(n_968), .C(n_970), .Y(n_966) );
CKINVDCx8_ASAP7_75t_R g1029 ( .A(n_911), .Y(n_1029) );
AOI211xp5_ASAP7_75t_L g1216 ( .A1(n_911), .A2(n_1091), .B(n_1217), .C(n_1218), .Y(n_1216) );
AOI221x1_ASAP7_75t_L g1231 ( .A1(n_913), .A2(n_1181), .B1(n_1232), .B2(n_1243), .C(n_1256), .Y(n_1231) );
OAI31xp33_ASAP7_75t_L g1581 ( .A1(n_913), .A2(n_1582), .A3(n_1583), .B(n_1589), .Y(n_1581) );
BUFx6f_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
AO211x2_ASAP7_75t_L g964 ( .A1(n_914), .A2(n_965), .B(n_978), .C(n_1008), .Y(n_964) );
AOI31xp33_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_929), .A3(n_936), .B(n_941), .Y(n_916) );
AOI211xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_920), .B(n_921), .C(n_924), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NOR3xp33_ASAP7_75t_L g1039 ( .A(n_921), .B(n_1040), .C(n_1044), .Y(n_1039) );
CKINVDCx11_ASAP7_75t_R g1077 ( .A(n_921), .Y(n_1077) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVxp67_ASAP7_75t_L g1084 ( .A(n_923), .Y(n_1084) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx2_ASAP7_75t_L g1012 ( .A(n_926), .Y(n_1012) );
INVx2_ASAP7_75t_L g1041 ( .A(n_926), .Y(n_1041) );
AOI322xp5_ASAP7_75t_L g1078 ( .A1(n_926), .A2(n_1074), .A3(n_1079), .B1(n_1080), .B2(n_1081), .C1(n_1082), .C2(n_1085), .Y(n_1078) );
AOI222xp33_ASAP7_75t_L g1247 ( .A1(n_926), .A2(n_1082), .B1(n_1248), .B2(n_1249), .C1(n_1250), .C2(n_1251), .Y(n_1247) );
INVx1_ASAP7_75t_L g1083 ( .A(n_928), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_932), .B1(n_933), .B2(n_935), .Y(n_929) );
AOI22xp33_ASAP7_75t_SL g1013 ( .A1(n_930), .A2(n_1014), .B1(n_1015), .B2(n_1016), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1045 ( .A1(n_930), .A2(n_1015), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_930), .A2(n_933), .B1(n_1184), .B2(n_1185), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_930), .A2(n_933), .B1(n_1245), .B2(n_1246), .Y(n_1244) );
AND2x4_ASAP7_75t_L g933 ( .A(n_931), .B(n_934), .Y(n_933) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_931), .B(n_934), .Y(n_1015) );
INVx1_ASAP7_75t_L g1074 ( .A(n_931), .Y(n_1074) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_937), .A2(n_974), .B1(n_1018), .B2(n_1019), .Y(n_1017) );
AOI211xp5_ASAP7_75t_L g1070 ( .A1(n_937), .A2(n_1071), .B(n_1072), .C(n_1076), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_937), .A2(n_939), .B1(n_1187), .B2(n_1188), .Y(n_1186) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_937), .A2(n_939), .B1(n_1237), .B2(n_1255), .Y(n_1254) );
INVx4_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx5_ASAP7_75t_L g1019 ( .A(n_940), .Y(n_1019) );
AOI31xp33_ASAP7_75t_L g1008 ( .A1(n_941), .A2(n_1009), .A3(n_1013), .B(n_1017), .Y(n_1008) );
AO21x1_ASAP7_75t_SL g1038 ( .A1(n_941), .A2(n_1039), .B(n_1045), .Y(n_1038) );
CKINVDCx16_ASAP7_75t_R g1181 ( .A(n_941), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_943), .B(n_956), .Y(n_942) );
BUFx3_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
NAND3xp33_ASAP7_75t_L g998 ( .A(n_945), .B(n_999), .C(n_1001), .Y(n_998) );
INVx3_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
A2O1A1Ixp33_ASAP7_75t_L g1153 ( .A1(n_955), .A2(n_1154), .B(n_1155), .C(n_1159), .Y(n_1153) );
XNOR2x1_ASAP7_75t_L g962 ( .A(n_963), .B(n_1020), .Y(n_962) );
NAND3xp33_ASAP7_75t_L g965 ( .A(n_966), .B(n_972), .C(n_975), .Y(n_965) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NAND4xp25_ASAP7_75t_L g978 ( .A(n_979), .B(n_988), .C(n_998), .D(n_1003), .Y(n_978) );
NAND3xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_984), .C(n_985), .Y(n_979) );
INVx3_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
NAND3xp33_ASAP7_75t_L g1265 ( .A(n_985), .B(n_1266), .C(n_1267), .Y(n_1265) );
INVx3_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
NAND3xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_995), .C(n_997), .Y(n_988) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx1_ASAP7_75t_L g1199 ( .A(n_993), .Y(n_1199) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx2_ASAP7_75t_L g1142 ( .A(n_994), .Y(n_1142) );
NAND3xp33_ASAP7_75t_L g1261 ( .A(n_997), .B(n_1262), .C(n_1264), .Y(n_1261) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1012), .Y(n_1192) );
INVx5_ASAP7_75t_SL g1075 ( .A(n_1015), .Y(n_1075) );
AND4x1_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1038), .C(n_1048), .D(n_1054), .Y(n_1021) );
NAND4xp25_ASAP7_75t_L g1062 ( .A(n_1022), .B(n_1038), .C(n_1048), .D(n_1054), .Y(n_1062) );
OAI31xp33_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1030), .A3(n_1033), .B(n_1037), .Y(n_1022) );
NAND3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1026), .C(n_1029), .Y(n_1023) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1035), .Y(n_1093) );
OAI31xp33_ASAP7_75t_SL g1086 ( .A1(n_1037), .A2(n_1087), .A3(n_1088), .B(n_1089), .Y(n_1086) );
INVx1_ASAP7_75t_SL g1228 ( .A(n_1037), .Y(n_1228) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1041), .Y(n_1594) );
OAI21xp33_ASAP7_75t_L g1150 ( .A1(n_1042), .A2(n_1151), .B(n_1152), .Y(n_1150) );
NAND3xp33_ASAP7_75t_L g1257 ( .A(n_1049), .B(n_1258), .C(n_1260), .Y(n_1257) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
XNOR2x1_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1177), .Y(n_1065) );
XNOR2x1_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1136), .Y(n_1066) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1068), .Y(n_1134) );
OAI211xp5_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .B(n_1086), .C(n_1096), .Y(n_1068) );
NAND4xp25_ASAP7_75t_SL g1182 ( .A(n_1077), .B(n_1183), .C(n_1186), .D(n_1189), .Y(n_1182) );
NAND4xp25_ASAP7_75t_SL g1243 ( .A(n_1077), .B(n_1244), .C(n_1247), .D(n_1254), .Y(n_1243) );
AND2x4_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1084), .Y(n_1082) );
AND2x4_ASAP7_75t_L g1595 ( .A(n_1083), .B(n_1084), .Y(n_1595) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
NOR2xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1118), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_1099), .A2(n_1100), .B1(n_1102), .B2(n_1103), .Y(n_1098) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
BUFx2_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1109), .Y(n_1537) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1116), .Y(n_1622) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
OAI22xp5_ASAP7_75t_L g1548 ( .A1(n_1123), .A2(n_1528), .B1(n_1529), .B2(n_1549), .Y(n_1548) );
OAI221xp5_ASAP7_75t_L g1608 ( .A1(n_1123), .A2(n_1609), .B1(n_1610), .B2(n_1612), .C(n_1613), .Y(n_1608) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
NAND4xp25_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1163), .C(n_1174), .D(n_1176), .Y(n_1137) );
OAI31xp33_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1160), .A3(n_1161), .B(n_1162), .Y(n_1138) );
OAI221xp5_ASAP7_75t_L g1139 ( .A1(n_1140), .A2(n_1144), .B1(n_1147), .B2(n_1150), .C(n_1153), .Y(n_1139) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1142), .Y(n_1201) );
INVx2_ASAP7_75t_SL g1259 ( .A(n_1142), .Y(n_1259) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
OA22x2_ASAP7_75t_L g1177 ( .A1(n_1178), .A2(n_1229), .B1(n_1230), .B2(n_1274), .Y(n_1177) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1178), .Y(n_1274) );
XNOR2xp5_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1180), .Y(n_1178) );
AOI211xp5_ASAP7_75t_L g1180 ( .A1(n_1181), .A2(n_1182), .B(n_1194), .C(n_1215), .Y(n_1180) );
OAI31xp33_ASAP7_75t_L g1590 ( .A1(n_1181), .A2(n_1591), .A3(n_1592), .B(n_1596), .Y(n_1590) );
NAND2xp5_ASAP7_75t_SL g1194 ( .A(n_1195), .B(n_1204), .Y(n_1194) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
AOI31xp33_ASAP7_75t_SL g1215 ( .A1(n_1216), .A2(n_1222), .A3(n_1225), .B(n_1228), .Y(n_1215) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1220), .Y(n_1240) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1231), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1236), .Y(n_1232) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
NAND4xp25_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1261), .C(n_1265), .D(n_1268), .Y(n_1256) );
OAI221xp5_ASAP7_75t_L g1277 ( .A1(n_1278), .A2(n_1517), .B1(n_1521), .B2(n_1566), .C(n_1571), .Y(n_1277) );
NOR2x1_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1457), .Y(n_1278) );
NAND4xp25_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1394), .C(n_1421), .D(n_1434), .Y(n_1279) );
A2O1A1Ixp33_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1306), .B(n_1336), .C(n_1382), .Y(n_1280) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1281), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1281), .B(n_1370), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1281), .B(n_1340), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1281), .B(n_1445), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1302), .Y(n_1281) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1282), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1282), .B(n_1303), .Y(n_1378) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1283), .B(n_1303), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1283), .B(n_1398), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1296), .Y(n_1283) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1291), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
OR2x2_ASAP7_75t_L g1332 ( .A(n_1287), .B(n_1292), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1290), .Y(n_1287) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1290), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1293 ( .A(n_1291), .B(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
OR2x2_ASAP7_75t_L g1335 ( .A(n_1292), .B(n_1295), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1636 ( .A(n_1294), .Y(n_1636) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1299), .Y(n_1297) );
AND2x4_ASAP7_75t_L g1301 ( .A(n_1298), .B(n_1300), .Y(n_1301) );
AND2x4_ASAP7_75t_L g1313 ( .A(n_1298), .B(n_1299), .Y(n_1313) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1301), .Y(n_1322) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1303), .Y(n_1339) );
INVxp67_ASAP7_75t_SL g1398 ( .A(n_1303), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1303), .B(n_1340), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1305), .Y(n_1303) );
NOR2xp33_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1324), .Y(n_1306) );
OAI221xp5_ASAP7_75t_L g1507 ( .A1(n_1307), .A2(n_1508), .B1(n_1513), .B2(n_1514), .C(n_1515), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1317), .Y(n_1307) );
INVx2_ASAP7_75t_L g1377 ( .A(n_1308), .Y(n_1377) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1308), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1314), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1309), .B(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1310), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1310), .B(n_1314), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1310), .B(n_1317), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1310), .B(n_1346), .Y(n_1410) );
BUFx6f_ASAP7_75t_L g1422 ( .A(n_1310), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1312), .Y(n_1310) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1313), .Y(n_1320) );
BUFx3_ASAP7_75t_L g1386 ( .A(n_1313), .Y(n_1386) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1314), .Y(n_1346) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1314), .Y(n_1360) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1314), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1314), .B(n_1349), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1314), .B(n_1326), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1316), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1317), .B(n_1345), .Y(n_1344) );
CKINVDCx6p67_ASAP7_75t_R g1349 ( .A(n_1317), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1317), .B(n_1355), .Y(n_1354) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1317), .B(n_1350), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1317), .B(n_1350), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1317), .B(n_1359), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_1317), .B(n_1384), .Y(n_1513) );
OR2x6_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_1318), .B(n_1319), .Y(n_1374) );
OAI22xp5_ASAP7_75t_SL g1319 ( .A1(n_1320), .A2(n_1321), .B1(n_1322), .B2(n_1323), .Y(n_1319) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1322), .Y(n_1328) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1322), .Y(n_1387) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1324), .B(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1325), .B(n_1369), .Y(n_1402) );
NOR2xp33_ASAP7_75t_L g1509 ( .A(n_1325), .B(n_1510), .Y(n_1509) );
BUFx3_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVx2_ASAP7_75t_SL g1356 ( .A(n_1326), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1326), .B(n_1366), .Y(n_1365) );
NOR2xp33_ASAP7_75t_L g1381 ( .A(n_1326), .B(n_1346), .Y(n_1381) );
BUFx2_ASAP7_75t_L g1430 ( .A(n_1326), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1326), .B(n_1340), .Y(n_1445) );
INVx2_ASAP7_75t_SL g1326 ( .A(n_1327), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1327), .B(n_1346), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1327), .B(n_1370), .Y(n_1399) );
OAI22xp33_ASAP7_75t_L g1329 ( .A1(n_1330), .A2(n_1331), .B1(n_1333), .B2(n_1334), .Y(n_1329) );
BUFx3_ASAP7_75t_L g1390 ( .A(n_1331), .Y(n_1390) );
BUFx6f_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
HB1xp67_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1335), .Y(n_1393) );
OAI211xp5_ASAP7_75t_L g1336 ( .A1(n_1337), .A2(n_1343), .B(n_1347), .C(n_1376), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1340), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1339), .B(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1339), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1339), .B(n_1340), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1340), .B(n_1352), .Y(n_1351) );
CKINVDCx5p33_ASAP7_75t_R g1370 ( .A(n_1340), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g1424 ( .A(n_1340), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1340), .B(n_1361), .Y(n_1436) );
NOR2xp33_ASAP7_75t_L g1452 ( .A(n_1340), .B(n_1362), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1340), .B(n_1397), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1340), .B(n_1362), .Y(n_1482) );
NOR2xp33_ASAP7_75t_L g1484 ( .A(n_1340), .B(n_1485), .Y(n_1484) );
AND2x4_ASAP7_75t_SL g1340 ( .A(n_1341), .B(n_1342), .Y(n_1340) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
AOI221xp5_ASAP7_75t_L g1470 ( .A1(n_1344), .A2(n_1397), .B1(n_1471), .B2(n_1472), .C(n_1473), .Y(n_1470) );
NAND3xp33_ASAP7_75t_L g1417 ( .A(n_1345), .B(n_1418), .C(n_1419), .Y(n_1417) );
AOI221xp5_ASAP7_75t_L g1498 ( .A1(n_1345), .A2(n_1360), .B1(n_1461), .B2(n_1499), .C(n_1502), .Y(n_1498) );
AOI211xp5_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1351), .B(n_1353), .C(n_1371), .Y(n_1347) );
AOI331xp33_ASAP7_75t_L g1421 ( .A1(n_1348), .A2(n_1382), .A3(n_1396), .B1(n_1422), .B2(n_1423), .B3(n_1428), .C1(n_1431), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1350), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1349), .B(n_1410), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1349), .B(n_1383), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1404 ( .A(n_1350), .B(n_1383), .Y(n_1404) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1350), .Y(n_1447) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1351), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1516 ( .A(n_1351), .B(n_1429), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1352), .B(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1352), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1380 ( .A(n_1352), .B(n_1381), .Y(n_1380) );
OAI321xp33_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1357), .A3(n_1361), .B1(n_1363), .B2(n_1364), .C(n_1367), .Y(n_1353) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1354), .Y(n_1418) );
INVxp67_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1356), .B(n_1436), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1464 ( .A(n_1356), .B(n_1465), .Y(n_1464) );
HB1xp67_ASAP7_75t_L g1468 ( .A(n_1356), .Y(n_1468) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1356), .B(n_1378), .Y(n_1501) );
O2A1O1Ixp33_ASAP7_75t_SL g1411 ( .A1(n_1357), .A2(n_1382), .B(n_1412), .C(n_1414), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1357), .B(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1358), .Y(n_1440) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1359), .B(n_1396), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1359), .B(n_1444), .Y(n_1443) );
INVx3_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1360), .B(n_1400), .Y(n_1438) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
AOI222xp33_ASAP7_75t_L g1508 ( .A1(n_1362), .A2(n_1368), .B1(n_1422), .B2(n_1509), .C1(n_1511), .C2(n_1512), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1366), .B(n_1463), .Y(n_1462) );
OAI221xp5_ASAP7_75t_SL g1493 ( .A1(n_1366), .A2(n_1494), .B1(n_1496), .B2(n_1497), .C(n_1498), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1369), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1368), .B(n_1430), .Y(n_1504) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1368), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1370), .B(n_1397), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1370), .B(n_1378), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1370), .B(n_1464), .Y(n_1463) );
OR2x2_ASAP7_75t_L g1500 ( .A(n_1370), .B(n_1501), .Y(n_1500) );
NOR2xp33_ASAP7_75t_L g1502 ( .A(n_1370), .B(n_1503), .Y(n_1502) );
NOR3xp33_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1374), .C(n_1375), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
A2O1A1Ixp33_ASAP7_75t_L g1376 ( .A1(n_1374), .A2(n_1377), .B(n_1378), .C(n_1379), .Y(n_1376) );
NOR2xp33_ASAP7_75t_L g1431 ( .A(n_1374), .B(n_1432), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1375), .B(n_1427), .Y(n_1426) );
OR2x2_ASAP7_75t_L g1476 ( .A(n_1375), .B(n_1477), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1378), .B(n_1399), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1378), .B(n_1445), .Y(n_1495) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1381), .B(n_1433), .Y(n_1432) );
INVx3_ASAP7_75t_L g1491 ( .A(n_1382), .Y(n_1491) );
A2O1A1Ixp33_ASAP7_75t_L g1515 ( .A1(n_1382), .A2(n_1440), .B(n_1446), .C(n_1516), .Y(n_1515) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
NOR2xp33_ASAP7_75t_L g1446 ( .A(n_1385), .B(n_1447), .Y(n_1446) );
OAI22xp33_ASAP7_75t_L g1388 ( .A1(n_1389), .A2(n_1390), .B1(n_1391), .B2(n_1392), .Y(n_1388) );
HB1xp67_ASAP7_75t_L g1520 ( .A(n_1392), .Y(n_1520) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
AOI221xp5_ASAP7_75t_L g1394 ( .A1(n_1395), .A2(n_1400), .B1(n_1401), .B2(n_1403), .C(n_1405), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1399), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1397), .B(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1397), .Y(n_1465) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1399), .Y(n_1477) );
AOI21xp5_ASAP7_75t_L g1479 ( .A1(n_1400), .A2(n_1480), .B(n_1486), .Y(n_1479) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
OAI221xp5_ASAP7_75t_L g1405 ( .A1(n_1406), .A2(n_1408), .B1(n_1411), .B2(n_1415), .C(n_1417), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1406), .B(n_1449), .Y(n_1471) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1410), .Y(n_1478) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1410), .B(n_1430), .Y(n_1496) );
CKINVDCx5p33_ASAP7_75t_R g1412 ( .A(n_1413), .Y(n_1412) );
AOI211xp5_ASAP7_75t_L g1458 ( .A1(n_1414), .A2(n_1459), .B(n_1462), .C(n_1466), .Y(n_1458) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
NOR2xp33_ASAP7_75t_L g1488 ( .A(n_1420), .B(n_1489), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_1422), .B(n_1488), .Y(n_1487) );
NOR2xp33_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1425), .Y(n_1423) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1429), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1429), .B(n_1484), .Y(n_1512) );
INVx2_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1430), .B(n_1447), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1483 ( .A(n_1430), .B(n_1484), .Y(n_1483) );
AOI221xp5_ASAP7_75t_L g1434 ( .A1(n_1435), .A2(n_1437), .B1(n_1439), .B2(n_1446), .C(n_1448), .Y(n_1434) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
OAI21xp33_ASAP7_75t_L g1439 ( .A1(n_1440), .A2(n_1441), .B(n_1443), .Y(n_1439) );
OAI21xp33_ASAP7_75t_L g1480 ( .A1(n_1440), .A2(n_1481), .B(n_1483), .Y(n_1480) );
AOI21xp33_ASAP7_75t_SL g1466 ( .A1(n_1441), .A2(n_1467), .B(n_1469), .Y(n_1466) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
AOI21xp5_ASAP7_75t_L g1448 ( .A1(n_1449), .A2(n_1450), .B(n_1453), .Y(n_1448) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
HB1xp67_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
A2O1A1Ixp33_ASAP7_75t_L g1457 ( .A1(n_1458), .A2(n_1470), .B(n_1490), .C(n_1492), .Y(n_1457) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1461), .B(n_1468), .Y(n_1467) );
A2O1A1Ixp33_ASAP7_75t_L g1473 ( .A1(n_1474), .A2(n_1476), .B(n_1478), .C(n_1479), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
NOR2xp33_ASAP7_75t_L g1494 ( .A(n_1475), .B(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
AOI21xp33_ASAP7_75t_SL g1492 ( .A1(n_1493), .A2(n_1505), .B(n_1507), .Y(n_1492) );
INVx2_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
INVxp67_ASAP7_75t_L g1514 ( .A(n_1512), .Y(n_1514) );
CKINVDCx5p33_ASAP7_75t_R g1517 ( .A(n_1518), .Y(n_1517) );
INVx1_ASAP7_75t_SL g1518 ( .A(n_1519), .Y(n_1518) );
BUFx2_ASAP7_75t_SL g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
AND4x1_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1543), .C(n_1545), .D(n_1563), .Y(n_1523) );
OAI21xp33_ASAP7_75t_SL g1550 ( .A1(n_1532), .A2(n_1551), .B(n_1552), .Y(n_1550) );
OAI22xp5_ASAP7_75t_L g1533 ( .A1(n_1534), .A2(n_1535), .B1(n_1536), .B2(n_1538), .Y(n_1533) );
INVx2_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
NOR2xp33_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1565), .Y(n_1563) );
CKINVDCx14_ASAP7_75t_R g1566 ( .A(n_1567), .Y(n_1566) );
INVx2_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
CKINVDCx5p33_ASAP7_75t_R g1568 ( .A(n_1569), .Y(n_1568) );
OAI21xp5_ASAP7_75t_L g1635 ( .A1(n_1570), .A2(n_1636), .B(n_1637), .Y(n_1635) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1580), .Y(n_1632) );
NAND3xp33_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1590), .C(n_1597), .Y(n_1580) );
HB1xp67_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
AOI22xp33_ASAP7_75t_L g1593 ( .A1(n_1587), .A2(n_1588), .B1(n_1594), .B2(n_1595), .Y(n_1593) );
NOR3xp33_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1607), .C(n_1623), .Y(n_1597) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
OAI21xp33_ASAP7_75t_SL g1625 ( .A1(n_1618), .A2(n_1626), .B(n_1627), .Y(n_1625) );
INVx2_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
INVx2_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
BUFx2_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
endmodule