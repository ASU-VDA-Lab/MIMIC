module fake_netlist_6_241_n_510 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_510);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_510;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_400;
wire n_284;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_491;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_493;
wire n_397;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_456;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_357;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_319;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_249;
wire n_201;
wire n_386;
wire n_487;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_404;
wire n_271;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVxp33_ASAP7_75t_L g167 ( 
.A(n_18),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_83),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_32),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_131),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_75),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_73),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_37),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_42),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_36),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_115),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_2),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_7),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_93),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_38),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_110),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_22),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_11),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_100),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_99),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_45),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_69),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_5),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_28),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_78),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_15),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_27),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_70),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_92),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_133),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_89),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_17),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_71),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_135),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_21),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_29),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_57),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g228 ( 
.A(n_41),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_126),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_68),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_77),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_122),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_91),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_112),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_72),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_76),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_132),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_87),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_26),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_141),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_31),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_59),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_123),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_43),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_23),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_60),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_46),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g250 ( 
.A(n_49),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_64),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_96),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_148),
.Y(n_253)
);

INVxp33_ASAP7_75t_SL g254 ( 
.A(n_62),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_66),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_162),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_48),
.Y(n_258)
);

INVxp33_ASAP7_75t_SL g259 ( 
.A(n_165),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_97),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_25),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_151),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_153),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_24),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_82),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_134),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_53),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_144),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_95),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_105),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_34),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_47),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_147),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_114),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_104),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_90),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_67),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_142),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_9),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_159),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_0),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_16),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_154),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_152),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_58),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_107),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_149),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_56),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_183),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_174),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_176),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_177),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_195),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_232),
.B(n_0),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_170),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_296)
);

CKINVDCx8_ASAP7_75t_R g297 ( 
.A(n_169),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_171),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_181),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_175),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_205),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_205),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g306 ( 
.A(n_229),
.B(n_12),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_206),
.A2(n_13),
.B1(n_19),
.B2(n_20),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_220),
.B(n_30),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_185),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_205),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_180),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_190),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_SL g313 ( 
.A(n_167),
.B(n_33),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_225),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_188),
.B(n_35),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_191),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_225),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_193),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_194),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_196),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_192),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_225),
.Y(n_322)
);

INVx3_ASAP7_75t_SL g323 ( 
.A(n_168),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_197),
.Y(n_324)
);

NAND2x1_ASAP7_75t_L g325 ( 
.A(n_229),
.B(n_39),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_201),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_244),
.B(n_40),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_202),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_203),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_204),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_247),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_207),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_222),
.B(n_44),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_230),
.B(n_245),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_208),
.B(n_50),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_209),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_210),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_218),
.B(n_51),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_211),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_248),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_250),
.B(n_52),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_212),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_254),
.B(n_54),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_217),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_221),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_226),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_333),
.A2(n_259),
.B1(n_263),
.B2(n_257),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_304),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_305),
.Y(n_352)
);

NAND2x1p5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_184),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_295),
.A2(n_255),
.B1(n_179),
.B2(n_187),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_328),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_300),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

NAND2x1p5_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_227),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_294),
.B(n_246),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_302),
.Y(n_364)
);

BUFx8_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_336),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_331),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g368 ( 
.A1(n_335),
.A2(n_287),
.B1(n_283),
.B2(n_282),
.Y(n_368)
);

AO22x2_ASAP7_75t_L g369 ( 
.A1(n_335),
.A2(n_251),
.B1(n_280),
.B2(n_279),
.Y(n_369)
);

AO22x2_ASAP7_75t_L g370 ( 
.A1(n_338),
.A2(n_243),
.B1(n_278),
.B2(n_277),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

OAI221xp5_ASAP7_75t_L g374 ( 
.A1(n_289),
.A2(n_249),
.B1(n_288),
.B2(n_216),
.C(n_233),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_299),
.B(n_189),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_313),
.A2(n_276),
.B1(n_262),
.B2(n_258),
.Y(n_376)
);

AO22x2_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_242),
.B1(n_275),
.B2(n_274),
.Y(n_377)
);

AO22x2_ASAP7_75t_L g378 ( 
.A1(n_343),
.A2(n_272),
.B1(n_269),
.B2(n_268),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_291),
.Y(n_379)
);

AO22x2_ASAP7_75t_L g380 ( 
.A1(n_298),
.A2(n_267),
.B1(n_266),
.B2(n_264),
.Y(n_380)
);

AO22x2_ASAP7_75t_L g381 ( 
.A1(n_329),
.A2(n_261),
.B1(n_253),
.B2(n_252),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_340),
.A2(n_241),
.B1(n_240),
.B2(n_239),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_292),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_323),
.B(n_231),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_293),
.Y(n_385)
);

BUFx8_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

BUFx12f_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_347),
.Y(n_388)
);

NAND2x1p5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_325),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_379),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_301),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_355),
.A2(n_334),
.B1(n_307),
.B2(n_303),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_383),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_309),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

BUFx8_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

BUFx12f_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_297),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_312),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_376),
.A2(n_327),
.B1(n_215),
.B2(n_199),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_346),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_374),
.A2(n_200),
.B1(n_228),
.B2(n_265),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_316),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_378),
.A2(n_182),
.B1(n_186),
.B2(n_198),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_384),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_358),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_392),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_394),
.A2(n_369),
.B1(n_368),
.B2(n_380),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_391),
.A2(n_306),
.B(n_359),
.Y(n_415)
);

AOI221x1_ASAP7_75t_SL g416 ( 
.A1(n_406),
.A2(n_289),
.B1(n_290),
.B2(n_296),
.C(n_337),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_403),
.A2(n_223),
.B(n_219),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_402),
.A2(n_235),
.B(n_234),
.C(n_236),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_407),
.A2(n_382),
.B1(n_381),
.B2(n_324),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_405),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_409),
.A2(n_381),
.B1(n_173),
.B2(n_178),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_390),
.Y(n_422)
);

INVx3_ASAP7_75t_SL g423 ( 
.A(n_412),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_357),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_321),
.Y(n_425)
);

BUFx4_ASAP7_75t_R g426 ( 
.A(n_387),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_396),
.A2(n_371),
.B(n_366),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_389),
.A2(n_397),
.B(n_393),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_361),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_350),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_238),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_352),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_399),
.B(n_356),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_285),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_L g436 ( 
.A1(n_431),
.A2(n_237),
.B(n_318),
.C(n_342),
.Y(n_436)
);

AOI221xp5_ASAP7_75t_L g437 ( 
.A1(n_416),
.A2(n_319),
.B1(n_320),
.B2(n_332),
.C(n_345),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_429),
.B(n_410),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_422),
.A2(n_344),
.B(n_351),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_410),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_270),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_415),
.A2(n_346),
.B(n_260),
.C(n_256),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_434),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_290),
.Y(n_444)
);

O2A1O1Ixp33_ASAP7_75t_SL g445 ( 
.A1(n_418),
.A2(n_284),
.B(n_271),
.C(n_224),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_416),
.A2(n_214),
.B(n_172),
.C(n_386),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_386),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_398),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_414),
.A2(n_55),
.B1(n_61),
.B2(n_63),
.Y(n_450)
);

AO32x2_ASAP7_75t_L g451 ( 
.A1(n_419),
.A2(n_421),
.A3(n_417),
.B1(n_430),
.B2(n_428),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_65),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_398),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_L g455 ( 
.A1(n_427),
.A2(n_74),
.B(n_80),
.C(n_81),
.Y(n_455)
);

AO22x2_ASAP7_75t_L g456 ( 
.A1(n_450),
.A2(n_446),
.B1(n_449),
.B2(n_448),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_439),
.A2(n_85),
.B(n_86),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_442),
.A2(n_88),
.B(n_101),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_444),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_106),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_438),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_452),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_454),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_108),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

AO21x1_ASAP7_75t_L g467 ( 
.A1(n_441),
.A2(n_451),
.B(n_453),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_451),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_451),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_457),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_462),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_462),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_464),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_463),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_465),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_461),
.Y(n_476)
);

AOI21xp33_ASAP7_75t_L g477 ( 
.A1(n_456),
.A2(n_436),
.B(n_437),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_455),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_467),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_480),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_459),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_468),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_469),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_485),
.B(n_470),
.Y(n_488)
);

NAND3x1_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_481),
.C(n_471),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_476),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_484),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_474),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_479),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_493),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_488),
.B(n_477),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_490),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_492),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_494),
.B(n_491),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g499 ( 
.A(n_497),
.B(n_478),
.Y(n_499)
);

CKINVDCx6p67_ASAP7_75t_R g500 ( 
.A(n_495),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_496),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_SL g502 ( 
.A(n_500),
.B(n_489),
.C(n_426),
.Y(n_502)
);

XNOR2x1_ASAP7_75t_L g503 ( 
.A(n_499),
.B(n_109),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_503),
.B(n_113),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_502),
.A2(n_501),
.B(n_445),
.Y(n_505)
);

XNOR2x1_ASAP7_75t_L g506 ( 
.A(n_504),
.B(n_116),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_505),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_507)
);

OAI322xp33_ASAP7_75t_L g508 ( 
.A1(n_507),
.A2(n_124),
.A3(n_127),
.B1(n_130),
.B2(n_136),
.C1(n_139),
.C2(n_146),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_508),
.Y(n_509)
);

AOI221xp5_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_506),
.B1(n_150),
.B2(n_155),
.C(n_161),
.Y(n_510)
);


endmodule