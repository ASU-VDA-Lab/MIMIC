module real_jpeg_14119_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_1),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_1),
.B(n_33),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_4),
.B(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_4),
.B(n_54),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_5),
.B(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_5),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_5),
.B(n_23),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_5),
.B(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_5),
.B(n_33),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_5),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_6),
.B(n_49),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_6),
.B(n_54),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_9),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_9),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_9),
.B(n_29),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_9),
.B(n_23),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_9),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_12),
.B(n_54),
.Y(n_61)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_94),
.CON(n_14),
.SN(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_80),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_17),
.B(n_80),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_55),
.B2(n_56),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_25),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_34),
.B(n_123),
.Y(n_122)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_46),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.C(n_42),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_40),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_41),
.B(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_50),
.B(n_123),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_70),
.B2(n_71),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_69),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_62),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.C(n_77),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.C(n_89),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_81),
.A2(n_82),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_97),
.C(n_102),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_134),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.CI(n_88),
.CON(n_85),
.SN(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_107),
.B(n_137),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_104),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_131),
.B(n_136),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_120),
.B(n_130),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_118),
.C(n_119),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_125),
.B(n_129),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);


endmodule