module fake_jpeg_10256_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_26),
.B1(n_35),
.B2(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_22),
.B1(n_27),
.B2(n_30),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_26),
.B1(n_35),
.B2(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_27),
.B1(n_22),
.B2(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_29),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_37),
.C(n_39),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_39),
.C(n_20),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_96),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_81),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_37),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_80),
.B(n_95),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_43),
.B1(n_35),
.B2(n_37),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_79),
.B1(n_88),
.B2(n_24),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_35),
.B1(n_19),
.B2(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_55),
.B(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_94),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_92),
.B(n_97),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_42),
.B1(n_30),
.B2(n_21),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_91),
.B(n_93),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_42),
.B(n_32),
.C(n_23),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_33),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_39),
.B(n_20),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_33),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_39),
.B1(n_41),
.B2(n_38),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_34),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_39),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_110),
.C(n_122),
.Y(n_133)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_118),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_0),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_120),
.B(n_31),
.Y(n_146)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_115),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_52),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_78),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_125),
.B1(n_73),
.B2(n_81),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_0),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_23),
.B(n_32),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_92),
.B(n_97),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_53),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_78),
.Y(n_123)
);

NOR4xp25_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_98),
.C(n_90),
.D(n_34),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_56),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_57),
.B1(n_65),
.B2(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_132),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_83),
.B(n_76),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_147),
.B(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_92),
.B1(n_77),
.B2(n_91),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_119),
.B1(n_102),
.B2(n_112),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_88),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_137),
.A2(n_143),
.B1(n_120),
.B2(n_123),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_140),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_125),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_87),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_145),
.C(n_155),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_146),
.B(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_149),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_98),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_99),
.B(n_111),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_154),
.B1(n_151),
.B2(n_128),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_97),
.B(n_54),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_90),
.B1(n_92),
.B2(n_97),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_92),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_159),
.B(n_174),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_165),
.B1(n_171),
.B2(n_175),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

AO22x1_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_108),
.B1(n_117),
.B2(n_110),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_169),
.B1(n_170),
.B2(n_178),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_105),
.B1(n_97),
.B2(n_103),
.Y(n_165)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_184),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_105),
.B1(n_48),
.B2(n_59),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_48),
.B1(n_59),
.B2(n_34),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_156),
.B1(n_147),
.B2(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_172),
.B(n_176),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_89),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_189),
.C(n_146),
.Y(n_193)
);

AOI32xp33_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_33),
.A3(n_32),
.B1(n_38),
.B2(n_28),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_24),
.B1(n_28),
.B2(n_86),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_139),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_24),
.B1(n_28),
.B2(n_86),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_182),
.B(n_183),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_141),
.B1(n_143),
.B2(n_155),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_86),
.B1(n_33),
.B2(n_32),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_188),
.B(n_25),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_133),
.B(n_38),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_216),
.Y(n_223)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_202),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_195),
.B(n_197),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_182),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_209),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_175),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_132),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_205),
.B(n_210),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_160),
.B(n_164),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_206),
.A2(n_207),
.B(n_211),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_135),
.B(n_145),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_38),
.C(n_25),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_170),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_38),
.B(n_25),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_213),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_25),
.C(n_31),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_31),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_221),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_198),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_225),
.B(n_227),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_158),
.B(n_164),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_244),
.C(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_242),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_159),
.B1(n_172),
.B2(n_163),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_243),
.B1(n_241),
.B2(n_232),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_165),
.B1(n_176),
.B2(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_1),
.B(n_2),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_212),
.B1(n_205),
.B2(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_218),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_199),
.C(n_193),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_258),
.C(n_259),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_228),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_250),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_227),
.Y(n_275)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_225),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_208),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_250),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_240),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_217),
.C(n_209),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_207),
.C(n_216),
.Y(n_259)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_190),
.C(n_192),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_263),
.C(n_251),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_190),
.C(n_192),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_234),
.A2(n_197),
.B1(n_202),
.B2(n_3),
.Y(n_265)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_257),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_265),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_249),
.Y(n_269)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_279),
.B(n_256),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_243),
.B(n_237),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_281),
.B(n_252),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_1),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_231),
.C(n_236),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_282),
.C(n_9),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_220),
.B(n_219),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_230),
.C(n_229),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_294),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_270),
.A2(n_255),
.B1(n_263),
.B2(n_261),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_293),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_259),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_295),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_222),
.B1(n_248),
.B2(n_258),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_273),
.B1(n_268),
.B2(n_277),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_296),
.C(n_276),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_9),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_278),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_274),
.C(n_272),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_271),
.B(n_285),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_300),
.A2(n_5),
.B(n_11),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_305),
.C(n_1),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_304),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_272),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_274),
.C(n_279),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_5),
.Y(n_314)
);

OAI221xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.C(n_4),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_10),
.B(n_12),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_288),
.B1(n_293),
.B2(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_16),
.B1(n_6),
.B2(n_4),
.Y(n_311)
);

OAI21x1_ASAP7_75t_SL g324 ( 
.A1(n_313),
.A2(n_317),
.B(n_12),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_297),
.B(n_301),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_298),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_305),
.B(n_317),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_297),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_323),
.B(n_324),
.Y(n_326)
);

OAI311xp33_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_327),
.A3(n_303),
.B1(n_321),
.C1(n_320),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_326),
.B1(n_12),
.B2(n_16),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_2),
.B(n_3),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_2),
.B(n_3),
.Y(n_332)
);


endmodule