module fake_ibex_291_n_361 (n_85, n_84, n_64, n_3, n_73, n_65, n_95, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_92, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_361);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_95;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_92;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_361;

wire n_151;
wire n_171;
wire n_103;
wire n_204;
wire n_274;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_124;
wire n_256;
wire n_193;
wire n_108;
wire n_350;
wire n_165;
wire n_255;
wire n_175;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_239;
wire n_134;
wire n_357;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_176;
wire n_216;
wire n_166;
wire n_163;
wire n_114;
wire n_236;
wire n_189;
wire n_280;
wire n_317;
wire n_340;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_113;
wire n_117;
wire n_265;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_210;
wire n_348;
wire n_220;
wire n_287;
wire n_243;
wire n_228;
wire n_147;
wire n_251;
wire n_244;
wire n_343;
wire n_310;
wire n_323;
wire n_143;
wire n_106;
wire n_224;
wire n_183;
wire n_333;
wire n_110;
wire n_306;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_109;
wire n_127;
wire n_121;
wire n_325;
wire n_301;
wire n_296;
wire n_120;
wire n_168;
wire n_155;
wire n_315;
wire n_122;
wire n_116;
wire n_289;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_235;
wire n_136;
wire n_261;
wire n_221;
wire n_355;
wire n_102;
wire n_99;
wire n_269;
wire n_156;
wire n_126;
wire n_356;
wire n_104;
wire n_141;
wire n_222;
wire n_186;
wire n_349;
wire n_295;
wire n_331;
wire n_230;
wire n_96;
wire n_185;
wire n_352;
wire n_290;
wire n_174;
wire n_157;
wire n_219;
wire n_246;
wire n_146;
wire n_207;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_139;
wire n_275;
wire n_129;
wire n_98;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_347;
wire n_335;
wire n_263;
wire n_353;
wire n_359;
wire n_262;
wire n_299;
wire n_137;
wire n_338;
wire n_173;
wire n_180;
wire n_201;
wire n_351;
wire n_257;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_179;
wire n_100;
wire n_354;
wire n_206;
wire n_329;
wire n_188;
wire n_200;
wire n_199;
wire n_308;
wire n_135;
wire n_283;
wire n_111;
wire n_322;
wire n_227;
wire n_115;
wire n_248;
wire n_101;
wire n_190;
wire n_138;
wire n_238;
wire n_214;
wire n_332;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_225;
wire n_360;
wire n_272;
wire n_223;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_148;
wire n_342;
wire n_233;
wire n_118;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_178;
wire n_303;
wire n_162;
wire n_240;
wire n_282;
wire n_266;
wire n_294;
wire n_112;
wire n_284;
wire n_172;
wire n_250;
wire n_313;
wire n_345;
wire n_119;
wire n_319;
wire n_195;
wire n_212;
wire n_311;
wire n_97;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_302;
wire n_344;
wire n_297;
wire n_252;
wire n_107;
wire n_149;
wire n_254;
wire n_213;
wire n_271;
wire n_241;
wire n_292;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_160;
wire n_184;
wire n_232;
wire n_281;

INVxp67_ASAP7_75t_SL g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_51),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_36),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_56),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_59),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_31),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_16),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_40),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_14),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_43),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_29),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_42),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_58),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_17),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_37),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_19),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_79),
.Y(n_138)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_70),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_60),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_0),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_77),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_68),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_38),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_32),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_49),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_22),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_83),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_2),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_18),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_13),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_55),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_1),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_46),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_23),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_6),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_9),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_87),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_7),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_41),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_0),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_54),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_2),
.Y(n_169)
);

BUFx2_ASAP7_75t_SL g170 ( 
.A(n_89),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_15),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_50),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_63),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_4),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_3),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_24),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_33),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

AO21x2_ASAP7_75t_L g184 ( 
.A1(n_101),
.A2(n_1),
.B(n_3),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

AND3x2_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_4),
.C(n_11),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_126),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_R g190 ( 
.A(n_156),
.B(n_28),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_30),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_107),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_109),
.B(n_135),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_128),
.B(n_103),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_62),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_109),
.B(n_73),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_109),
.B(n_76),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_135),
.B(n_85),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_135),
.B(n_90),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_130),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_133),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_110),
.B(n_129),
.Y(n_213)
);

NAND2xp33_ASAP7_75t_L g214 ( 
.A(n_151),
.B(n_94),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_136),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_145),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_146),
.B(n_179),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_147),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_152),
.B(n_159),
.C(n_171),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_170),
.B(n_162),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_153),
.B(n_154),
.Y(n_226)
);

NAND2xp33_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_178),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_150),
.A2(n_174),
.B1(n_168),
.B2(n_117),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_100),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_122),
.B(n_155),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_134),
.A2(n_96),
.B1(n_158),
.B2(n_140),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_98),
.B(n_99),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_139),
.B(n_175),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_102),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_105),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_120),
.B(n_123),
.C(n_127),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_215),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_113),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_148),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_149),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_144),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_185),
.B(n_161),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_131),
.B1(n_132),
.B2(n_138),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_164),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g254 ( 
.A(n_187),
.B(n_166),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_213),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_143),
.B1(n_172),
.B2(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_183),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

OR2x6_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_181),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

BUFx4f_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_196),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_191),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

BUFx4f_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_229),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_196),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_221),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_194),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_186),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_233),
.B(n_224),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_236),
.A2(n_233),
.B1(n_224),
.B2(n_227),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_226),
.B(n_203),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_195),
.A2(n_208),
.B1(n_217),
.B2(n_211),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_204),
.B(n_228),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_204),
.B(n_200),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_222),
.B(n_184),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_228),
.B(n_201),
.Y(n_289)
);

OA22x2_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_184),
.B1(n_206),
.B2(n_205),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_214),
.B(n_207),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_242),
.A2(n_209),
.B(n_201),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_222),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_288),
.A2(n_190),
.B(n_222),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

OAI22x1_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_255),
.B1(n_249),
.B2(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_264),
.B(n_272),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_280),
.B(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_281),
.A2(n_241),
.B(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_248),
.B(n_246),
.Y(n_304)
);

AO31x2_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_266),
.A3(n_263),
.B(n_268),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_244),
.A2(n_245),
.B(n_247),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_243),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_267),
.B(n_258),
.Y(n_309)
);

AO31x2_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_273),
.A3(n_283),
.B(n_257),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_262),
.A2(n_259),
.B(n_254),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_256),
.A2(n_250),
.B1(n_254),
.B2(n_251),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_277),
.B(n_285),
.C(n_279),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_240),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_240),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_240),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_303),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_292),
.A2(n_279),
.B(n_282),
.C(n_307),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_297),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_309),
.Y(n_322)
);

AOI221xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_279),
.B1(n_282),
.B2(n_300),
.C(n_306),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_290),
.A2(n_282),
.B1(n_304),
.B2(n_311),
.Y(n_324)
);

O2A1O1Ixp5_ASAP7_75t_L g325 ( 
.A1(n_293),
.A2(n_291),
.B(n_299),
.C(n_310),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_310),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_294),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_297),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_321),
.Y(n_333)
);

AO31x2_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_315),
.A3(n_320),
.B(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_327),
.B(n_325),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_330),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_329),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_SL g340 ( 
.A(n_323),
.B(n_326),
.C(n_325),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_332),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_335),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_337),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_314),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_339),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_331),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_343),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_342),
.B(n_333),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

NAND4xp25_ASAP7_75t_L g352 ( 
.A(n_350),
.B(n_341),
.C(n_340),
.D(n_324),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_351),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_352),
.A2(n_349),
.B(n_322),
.Y(n_354)
);

NOR2x1_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_348),
.Y(n_355)
);

NOR3xp33_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_347),
.C(n_346),
.Y(n_356)
);

AOI221xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_353),
.B1(n_341),
.B2(n_331),
.C(n_345),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_357),
.A2(n_346),
.B1(n_341),
.B2(n_345),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_345),
.B1(n_344),
.B2(n_346),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_359),
.A2(n_344),
.B(n_336),
.Y(n_360)
);

AOI221xp5_ASAP7_75t_L g361 ( 
.A1(n_360),
.A2(n_318),
.B1(n_316),
.B2(n_344),
.C(n_334),
.Y(n_361)
);


endmodule