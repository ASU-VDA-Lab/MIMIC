module real_jpeg_6687_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_286;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_297;
wire n_180;
wire n_58;
wire n_52;
wire n_209;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_295;
wire n_167;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_0),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_0),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_1),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_1),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_1),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_1),
.B(n_229),
.Y(n_228)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_3),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_3),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_3),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_3),
.B(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_4),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_5),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_5),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_5),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_5),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_5),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_5),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_5),
.B(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_7),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_8),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_8),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_8),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_8),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_8),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_9),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_9),
.B(n_28),
.Y(n_175)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_12),
.Y(n_91)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_13),
.Y(n_117)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_13),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_13),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_14),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_15),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_15),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_182),
.B1(n_183),
.B2(n_304),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_18),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_180),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_156),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_20),
.B(n_156),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_55),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_23),
.B(n_178),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_23),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_31),
.CI(n_35),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_31),
.C(n_35),
.Y(n_155)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_28),
.Y(n_240)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_29),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_37),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_38),
.Y(n_129)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_38),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_39),
.A2(n_55),
.B1(n_56),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_39),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_52),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_40),
.A2(n_52),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_40),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_70),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_41),
.B(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_44),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_45),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_45),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_46),
.B(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_52),
.Y(n_164)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_176)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_60),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_60),
.Y(n_259)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_84),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_72),
.Y(n_174)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_73),
.Y(n_218)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_76),
.A2(n_83),
.B1(n_125),
.B2(n_126),
.Y(n_223)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_93),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_86),
.B(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_92),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_97),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_97),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_97),
.B(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_140),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_120),
.C(n_122),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_103),
.A2(n_120),
.B1(n_121),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_119),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_109),
.C(n_115),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_107),
.Y(n_222)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_107),
.Y(n_233)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.C(n_136),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_123),
.A2(n_124),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_130),
.A2(n_131),
.B1(n_136),
.B2(n_137),
.Y(n_296)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_155),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.C(n_177),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_157),
.A2(n_158),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_161),
.B(n_177),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_176),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_162),
.B(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_166),
.B(n_176),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.C(n_175),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_298),
.B(n_303),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_283),
.B(n_297),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_235),
.B(n_282),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_224),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_187),
.B(n_224),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_209),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_205),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_189),
.B(n_205),
.C(n_209),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_196),
.C(n_201),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_219),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_210),
.B(n_292),
.C(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.C(n_234),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_225),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_234),
.B1(n_274),
.B2(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_276),
.B(n_281),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_261),
.B(n_275),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_245),
.B(n_260),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_256),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_256),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_251),
.B(n_255),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_251),
.Y(n_255)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_263),
.B1(n_269),
.B2(n_270),
.Y(n_262)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_271),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_271),
.Y(n_275)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_264),
.A2(n_266),
.B(n_269),
.Y(n_277)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_285),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_291),
.C(n_294),
.Y(n_299)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);


endmodule