module fake_jpeg_28473_n_376 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_376);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_376;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_50),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_10),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_51),
.B(n_53),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_10),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_11),
.C(n_9),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_45),
.C(n_29),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_64),
.Y(n_107)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_24),
.B(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_70),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g106 ( 
.A(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_39),
.B(n_11),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_72),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_74),
.Y(n_147)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_9),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_80),
.Y(n_114)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_9),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_82),
.Y(n_139)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_86),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_88),
.Y(n_120)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_90),
.Y(n_121)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_92),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_45),
.B(n_3),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_97),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_29),
.B1(n_42),
.B2(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_18),
.B(n_4),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_32),
.Y(n_141)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_105),
.A2(n_123),
.B1(n_130),
.B2(n_142),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_122),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_112),
.A2(n_106),
.B1(n_102),
.B2(n_117),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_42),
.B(n_5),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_32),
.B1(n_44),
.B2(n_40),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_50),
.A2(n_37),
.B1(n_31),
.B2(n_27),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_52),
.A2(n_60),
.B1(n_56),
.B2(n_86),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_64),
.A2(n_85),
.B1(n_42),
.B2(n_87),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_61),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_107),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_85),
.A2(n_42),
.B1(n_27),
.B2(n_23),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_59),
.A2(n_35),
.B1(n_44),
.B2(n_40),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_150),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_63),
.A2(n_35),
.B1(n_38),
.B2(n_46),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_51),
.A2(n_38),
.B1(n_46),
.B2(n_6),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_148),
.B1(n_142),
.B2(n_123),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_53),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_72),
.B(n_8),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_110),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_89),
.A2(n_8),
.B1(n_91),
.B2(n_92),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_8),
.B1(n_134),
.B2(n_141),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_8),
.B1(n_139),
.B2(n_114),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_164),
.B1(n_178),
.B2(n_183),
.Y(n_196)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_118),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_158),
.B(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_118),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_163),
.Y(n_215)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_171),
.Y(n_199)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_175),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_191),
.B(n_147),
.Y(n_212)
);

BUFx2_ASAP7_75t_SL g174 ( 
.A(n_106),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_179),
.Y(n_224)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_104),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_176),
.B(n_177),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_111),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_109),
.A2(n_113),
.B1(n_139),
.B2(n_114),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_103),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_180),
.B(n_181),
.Y(n_222)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_113),
.A2(n_154),
.B1(n_127),
.B2(n_115),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_106),
.B1(n_133),
.B2(n_125),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_109),
.A2(n_139),
.B1(n_114),
.B2(n_143),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_185),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_121),
.B1(n_107),
.B2(n_120),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_192),
.B1(n_151),
.B2(n_101),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_187),
.A2(n_133),
.B1(n_102),
.B2(n_117),
.Y(n_195)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_147),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_190),
.B(n_128),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_107),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_124),
.A2(n_101),
.B1(n_127),
.B2(n_125),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_194),
.Y(n_213)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_207),
.B1(n_211),
.B2(n_223),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_170),
.B(n_128),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_170),
.B(n_150),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_131),
.C(n_116),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_210),
.C(n_221),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_131),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_165),
.A2(n_115),
.B1(n_144),
.B2(n_146),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_159),
.B(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_160),
.B(n_146),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_158),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_168),
.A2(n_144),
.B1(n_147),
.B2(n_186),
.Y(n_223)
);

AOI32xp33_ASAP7_75t_L g225 ( 
.A1(n_160),
.A2(n_157),
.A3(n_165),
.B1(n_192),
.B2(n_161),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_194),
.Y(n_235)
);

NAND2xp33_ASAP7_75t_SL g270 ( 
.A(n_227),
.B(n_198),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_228),
.A2(n_224),
.B(n_223),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_233),
.Y(n_261)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_225),
.A2(n_171),
.B1(n_181),
.B2(n_162),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_196),
.A2(n_167),
.B1(n_169),
.B2(n_188),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_203),
.B1(n_204),
.B2(n_219),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_199),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_175),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_238),
.Y(n_251)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_179),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_214),
.C(n_221),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_210),
.C(n_196),
.Y(n_262)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_166),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_245),
.B(n_199),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

BUFx12f_ASAP7_75t_SL g247 ( 
.A(n_212),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_212),
.B(n_203),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_252),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_199),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_255),
.B(n_258),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_236),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_263),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_266),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_270),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_238),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_222),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_205),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_231),
.B(n_229),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_249),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_247),
.B(n_227),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_241),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_258),
.C(n_268),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_226),
.B1(n_235),
.B2(n_248),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_285),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_241),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_257),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_243),
.B(n_226),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_289),
.Y(n_293)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_281),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_200),
.A3(n_244),
.B1(n_231),
.B2(n_243),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_242),
.B1(n_234),
.B2(n_246),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_263),
.B1(n_256),
.B2(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_215),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_252),
.A2(n_224),
.B(n_216),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_264),
.Y(n_294)
);

OAI32xp33_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_207),
.A3(n_220),
.B1(n_216),
.B2(n_215),
.Y(n_292)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_304),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_269),
.B1(n_277),
.B2(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_251),
.C(n_259),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_301),
.B(n_305),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_283),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_286),
.A2(n_252),
.B1(n_264),
.B2(n_250),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_273),
.B(n_251),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_283),
.A2(n_252),
.B(n_260),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_309),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_260),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_282),
.Y(n_315)
);

XOR2x1_ASAP7_75t_SL g313 ( 
.A(n_295),
.B(n_274),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_323),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_321),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_282),
.C(n_278),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_324),
.C(n_303),
.Y(n_334)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_307),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_284),
.Y(n_323)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_276),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_336),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_293),
.B(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_302),
.B1(n_299),
.B2(n_306),
.Y(n_329)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_313),
.A2(n_264),
.B1(n_291),
.B2(n_288),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_335),
.B(n_304),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_302),
.Y(n_331)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_318),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_264),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_299),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_322),
.B(n_287),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_337),
.B(n_326),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_340),
.A2(n_290),
.B(n_335),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_341),
.A2(n_254),
.B1(n_267),
.B2(n_307),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_318),
.C(n_333),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_348),
.C(n_346),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_338),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_323),
.C(n_316),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_SL g349 ( 
.A(n_340),
.B(n_330),
.Y(n_349)
);

NAND5xp2_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_270),
.C(n_253),
.D(n_265),
.E(n_230),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_350),
.A2(n_354),
.B1(n_253),
.B2(n_265),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_351),
.B(n_353),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_347),
.A2(n_291),
.B(n_287),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_352),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_343),
.A2(n_324),
.B1(n_292),
.B2(n_254),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_355),
.B(n_342),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_357),
.B(n_358),
.Y(n_366)
);

AOI322xp5_ASAP7_75t_L g358 ( 
.A1(n_352),
.A2(n_344),
.A3(n_345),
.B1(n_348),
.B2(n_339),
.C1(n_281),
.C2(n_321),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_356),
.A2(n_267),
.B1(n_315),
.B2(n_338),
.Y(n_359)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_359),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_363),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_362),
.A2(n_355),
.B(n_350),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_364),
.A2(n_237),
.B(n_253),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_351),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_368),
.B(n_358),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_369),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_370),
.A2(n_371),
.B(n_367),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_218),
.C(n_219),
.Y(n_371)
);

AOI311xp33_ASAP7_75t_L g374 ( 
.A1(n_372),
.A2(n_365),
.A3(n_367),
.B(n_218),
.C(n_163),
.Y(n_374)
);

OAI21x1_ASAP7_75t_L g375 ( 
.A1(n_374),
.A2(n_373),
.B(n_156),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_375),
.B(n_187),
.Y(n_376)
);


endmodule