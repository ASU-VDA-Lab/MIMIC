module fake_jpeg_1027_n_501 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_501);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_501;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g56 ( 
.A(n_13),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_58),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_18),
.C(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_61),
.B(n_68),
.Y(n_124)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_56),
.Y(n_63)
);

CKINVDCx6p67_ASAP7_75t_R g182 ( 
.A(n_63),
.Y(n_182)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_64),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_15),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_71),
.Y(n_168)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_73),
.B(n_80),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_74),
.B(n_106),
.Y(n_129)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_75),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_76),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_1),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_38),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_84),
.B(n_95),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_86),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_89),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_92),
.B(n_99),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_107),
.B1(n_119),
.B2(n_50),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_26),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_2),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_96),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx12f_ASAP7_75t_SL g158 ( 
.A(n_97),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_3),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_3),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_112),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_101),
.B(n_103),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_105),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_109),
.Y(n_128)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_115),
.Y(n_136)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_47),
.B(n_13),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_117),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_SL g152 ( 
.A(n_116),
.Y(n_152)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_22),
.B(n_4),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_122),
.Y(n_146)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_121),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_39),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_51),
.B1(n_50),
.B2(n_55),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_127),
.A2(n_134),
.B1(n_156),
.B2(n_179),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_132),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_58),
.A2(n_51),
.B1(n_27),
.B2(n_49),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_107),
.A2(n_24),
.B1(n_54),
.B2(n_42),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_137),
.A2(n_142),
.B1(n_144),
.B2(n_159),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_94),
.A2(n_24),
.B1(n_54),
.B2(n_42),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_61),
.A2(n_55),
.B1(n_36),
.B2(n_28),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_148),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_73),
.B(n_36),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_87),
.A2(n_28),
.B1(n_48),
.B2(n_44),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_154),
.A2(n_166),
.B1(n_170),
.B2(n_197),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_90),
.A2(n_19),
.B1(n_48),
.B2(n_44),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_68),
.A2(n_49),
.B1(n_41),
.B2(n_39),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_163),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_80),
.B(n_41),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_165),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_84),
.B(n_23),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_91),
.A2(n_20),
.B1(n_19),
.B2(n_23),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_95),
.B(n_20),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_167),
.B(n_177),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_75),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_172),
.A2(n_192),
.B1(n_201),
.B2(n_205),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_98),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_174),
.A2(n_185),
.B1(n_194),
.B2(n_134),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_100),
.B(n_5),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_105),
.A2(n_13),
.B1(n_9),
.B2(n_11),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_12),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_110),
.B(n_8),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_196),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_65),
.B(n_8),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_184),
.B(n_186),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_93),
.A2(n_8),
.B1(n_9),
.B2(n_66),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_72),
.B(n_79),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_77),
.B(n_123),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_188),
.B(n_200),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_115),
.A2(n_120),
.B1(n_121),
.B2(n_78),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_70),
.A2(n_62),
.B1(n_57),
.B2(n_59),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_76),
.B(n_74),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_82),
.A2(n_102),
.B1(n_105),
.B2(n_121),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_74),
.B(n_112),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_107),
.A2(n_56),
.B1(n_43),
.B2(n_119),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_107),
.A2(n_56),
.B1(n_43),
.B2(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_209),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g210 ( 
.A(n_139),
.B(n_151),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_210),
.B(n_222),
.Y(n_312)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_212),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_157),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_214),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_183),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_216),
.B(n_220),
.Y(n_286)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_218),
.B(n_219),
.Y(n_282)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_129),
.B(n_130),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_171),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_221),
.B(n_245),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_130),
.B(n_187),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_223),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_124),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_168),
.C(n_203),
.Y(n_277)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_136),
.A2(n_145),
.B1(n_197),
.B2(n_170),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_227),
.A2(n_238),
.B1(n_241),
.B2(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_229),
.Y(n_290)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_154),
.A2(n_166),
.B1(n_185),
.B2(n_125),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_230),
.A2(n_257),
.B(n_217),
.C(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_231),
.Y(n_293)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_133),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_234),
.B(n_257),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_182),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_236),
.B(n_239),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_237),
.B(n_255),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_124),
.B1(n_125),
.B2(n_136),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_182),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_133),
.A2(n_178),
.B1(n_194),
.B2(n_180),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_240),
.A2(n_255),
.B1(n_254),
.B2(n_243),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_145),
.A2(n_131),
.B1(n_135),
.B2(n_175),
.Y(n_241)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_242),
.Y(n_300)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_135),
.A2(n_175),
.B1(n_199),
.B2(n_190),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_150),
.Y(n_248)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_178),
.A2(n_157),
.B1(n_138),
.B2(n_128),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_249),
.B(n_265),
.Y(n_303)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_199),
.A2(n_190),
.B1(n_157),
.B2(n_204),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_251),
.A2(n_153),
.B1(n_169),
.B2(n_198),
.Y(n_294)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_158),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_182),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_256),
.B(n_259),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_148),
.B(n_156),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_127),
.A2(n_169),
.B1(n_191),
.B2(n_150),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_153),
.B1(n_143),
.B2(n_160),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_178),
.B(n_140),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_148),
.B(n_189),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_261),
.B(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_152),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_171),
.A2(n_158),
.B(n_155),
.C(n_180),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_264),
.A2(n_243),
.B(n_242),
.Y(n_310)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_171),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_269),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_147),
.B(n_189),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_147),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_274),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_149),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_271),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_143),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_272),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_SL g273 ( 
.A(n_140),
.B(n_168),
.C(n_198),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_155),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_277),
.B(n_248),
.Y(n_340)
);

XOR2x2_ASAP7_75t_L g278 ( 
.A(n_211),
.B(n_155),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_314),
.C(n_267),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_216),
.B(n_160),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_280),
.B(n_252),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_291),
.B1(n_294),
.B2(n_308),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_237),
.A2(n_211),
.B1(n_215),
.B2(n_214),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_155),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_296),
.B(n_299),
.Y(n_319)
);

OAI32xp33_ASAP7_75t_L g297 ( 
.A1(n_220),
.A2(n_149),
.A3(n_173),
.B1(n_214),
.B2(n_234),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_310),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_208),
.B(n_173),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_226),
.B(n_246),
.Y(n_333)
);

NOR2x1p5_ASAP7_75t_SL g306 ( 
.A(n_249),
.B(n_209),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_230),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_227),
.A2(n_230),
.B1(n_206),
.B2(n_207),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_213),
.B(n_210),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_313),
.B(n_316),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_224),
.B(n_207),
.C(n_268),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_235),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_230),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_322),
.B(n_338),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_325),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_206),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_332),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_254),
.B1(n_241),
.B2(n_251),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_327),
.A2(n_344),
.B1(n_348),
.B2(n_349),
.Y(n_387)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_288),
.Y(n_330)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_330),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_295),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g369 ( 
.A1(n_333),
.A2(n_310),
.B(n_298),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_292),
.A2(n_212),
.B1(n_228),
.B2(n_229),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_337),
.Y(n_383)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_307),
.Y(n_336)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_292),
.A2(n_231),
.B1(n_272),
.B2(n_253),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_295),
.A2(n_264),
.B(n_265),
.C(n_260),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_290),
.Y(n_339)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_340),
.B(n_277),
.Y(n_373)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_341),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_342),
.B(n_343),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_280),
.B(n_232),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_291),
.A2(n_247),
.B1(n_225),
.B2(n_223),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_248),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_345),
.B(n_352),
.Y(n_366)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_346),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_233),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_285),
.C(n_284),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_263),
.B1(n_271),
.B2(n_270),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_302),
.A2(n_250),
.B1(n_274),
.B2(n_298),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_304),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_350),
.Y(n_381)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_279),
.B(n_316),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_353),
.B(n_354),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_279),
.B(n_299),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_303),
.A2(n_297),
.B(n_306),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_355),
.A2(n_357),
.B(n_303),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_356),
.Y(n_376)
);

AOI32xp33_ASAP7_75t_L g357 ( 
.A1(n_306),
.A2(n_303),
.A3(n_313),
.B1(n_305),
.B2(n_298),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_344),
.B(n_327),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_369),
.A2(n_379),
.B(n_330),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_326),
.A2(n_276),
.B1(n_278),
.B2(n_309),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_371),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_321),
.A2(n_276),
.B1(n_278),
.B2(n_309),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_373),
.B(n_374),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_312),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_321),
.A2(n_294),
.B1(n_318),
.B2(n_275),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_375),
.A2(n_348),
.B1(n_329),
.B2(n_328),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_318),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_378),
.B(n_349),
.Y(n_398)
);

AO21x1_ASAP7_75t_L g379 ( 
.A1(n_335),
.A2(n_311),
.B(n_285),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_356),
.C(n_284),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_345),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_385),
.B(n_388),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_334),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_322),
.A2(n_275),
.B1(n_296),
.B2(n_315),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_338),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_369),
.A2(n_323),
.B(n_355),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_390),
.A2(n_396),
.B(n_399),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_347),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_401),
.C(n_414),
.Y(n_431)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_367),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_400),
.Y(n_421)
);

OAI322xp33_ASAP7_75t_L g394 ( 
.A1(n_385),
.A2(n_324),
.A3(n_335),
.B1(n_331),
.B2(n_319),
.C1(n_343),
.C2(n_340),
.Y(n_394)
);

AOI322xp5_ASAP7_75t_SL g429 ( 
.A1(n_394),
.A2(n_282),
.A3(n_360),
.B1(n_377),
.B2(n_381),
.C1(n_384),
.C2(n_372),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_369),
.A2(n_335),
.B(n_323),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_363),
.Y(n_397)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_397),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_379),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_379),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_366),
.B(n_320),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_405),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_386),
.B(n_333),
.C(n_339),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_361),
.C(n_380),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_404),
.A2(n_415),
.B(n_381),
.Y(n_434)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_366),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_407),
.Y(n_426)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_378),
.B(n_352),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_409),
.Y(n_433)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_410),
.A2(n_388),
.B1(n_387),
.B2(n_383),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_358),
.A2(n_351),
.B(n_336),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_413),
.A2(n_289),
.B(n_376),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_386),
.B(n_337),
.Y(n_414)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_416),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_423),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_400),
.A2(n_365),
.B1(n_383),
.B2(n_376),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_418),
.A2(n_428),
.B1(n_399),
.B2(n_406),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_391),
.B(n_374),
.C(n_370),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_422),
.C(n_432),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_365),
.C(n_371),
.Y(n_422)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_424),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_390),
.A2(n_389),
.B(n_375),
.Y(n_427)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_427),
.A2(n_434),
.B(n_437),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_410),
.A2(n_362),
.B1(n_367),
.B2(n_360),
.Y(n_428)
);

OAI322xp33_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_399),
.A3(n_426),
.B1(n_412),
.B2(n_425),
.C1(n_421),
.C2(n_433),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_395),
.B(n_414),
.C(n_403),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_384),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_415),
.C(n_401),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_415),
.A2(n_377),
.B(n_372),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_440),
.Y(n_456)
);

NOR3xp33_ASAP7_75t_SL g440 ( 
.A(n_421),
.B(n_411),
.C(n_412),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_420),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_429),
.B(n_428),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_411),
.C(n_408),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_448),
.C(n_422),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_418),
.A2(n_396),
.B1(n_402),
.B2(n_394),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_446),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_416),
.A2(n_413),
.B1(n_409),
.B2(n_407),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_431),
.B(n_282),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_449),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_431),
.C(n_417),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_437),
.A2(n_405),
.B1(n_397),
.B2(n_392),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_426),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_453),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_425),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_432),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_SL g468 ( 
.A(n_455),
.B(n_458),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_457),
.A2(n_445),
.B(n_439),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_417),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_448),
.B(n_422),
.C(n_436),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_460),
.B(n_467),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_463),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_423),
.C(n_420),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_466),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_424),
.C(n_434),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_382),
.C(n_359),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_456),
.A2(n_452),
.B1(n_464),
.B2(n_450),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_469),
.A2(n_472),
.B1(n_476),
.B2(n_350),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_462),
.A2(n_451),
.B(n_450),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_470),
.A2(n_478),
.B(n_350),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_471),
.B(n_472),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_459),
.A2(n_451),
.B1(n_442),
.B2(n_427),
.Y(n_472)
);

OAI221xp5_ASAP7_75t_L g475 ( 
.A1(n_461),
.A2(n_433),
.B1(n_441),
.B2(n_440),
.C(n_442),
.Y(n_475)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_475),
.Y(n_481)
);

AOI221xp5_ASAP7_75t_L g476 ( 
.A1(n_462),
.A2(n_449),
.B1(n_446),
.B2(n_430),
.C(n_435),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_466),
.A2(n_442),
.B(n_435),
.Y(n_478)
);

NOR2x1_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_463),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_479),
.A2(n_484),
.B(n_485),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_477),
.A2(n_458),
.B1(n_430),
.B2(n_359),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_470),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_368),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_486),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_483),
.Y(n_491)
);

AOI221xp5_ASAP7_75t_L g484 ( 
.A1(n_478),
.A2(n_341),
.B1(n_346),
.B2(n_455),
.C(n_315),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_473),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_492),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_488),
.B(n_483),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_468),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_493),
.B(n_495),
.C(n_491),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_490),
.B(n_479),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_283),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_491),
.B(n_300),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_498),
.B(n_317),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_497),
.A2(n_494),
.B(n_493),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_499),
.B(n_500),
.Y(n_501)
);


endmodule