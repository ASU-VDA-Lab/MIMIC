module real_aes_4398_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_1106, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_1106;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_1067;
wire n_518;
wire n_792;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_1034;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_626;
wire n_539;
wire n_400;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_1078;
wire n_495;
wire n_994;
wire n_892;
wire n_370;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_1053;
wire n_466;
wire n_636;
wire n_559;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_1086;
wire n_343;
wire n_369;
wire n_1070;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_298;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_733;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_1041;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1028;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_1043;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_1090;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_756;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_1045;
wire n_465;
wire n_473;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_1055;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_652;
wire n_703;
wire n_393;
wire n_500;
wire n_307;
wire n_1101;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_802;
wire n_877;
wire n_868;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_1104;
wire n_842;
wire n_1061;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_0), .A2(n_122), .B1(n_359), .B2(n_636), .Y(n_667) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_1), .Y(n_308) );
AND2x4_ASAP7_75t_L g810 ( .A(n_1), .B(n_811), .Y(n_810) );
AND2x4_ASAP7_75t_L g819 ( .A(n_1), .B(n_288), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_2), .A2(n_244), .B1(n_375), .B2(n_633), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_3), .A2(n_135), .B1(n_822), .B2(n_836), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_4), .A2(n_178), .B1(n_790), .B2(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g598 ( .A(n_5), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_6), .A2(n_226), .B1(n_851), .B2(n_853), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_7), .A2(n_66), .B1(n_405), .B2(n_612), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_8), .A2(n_294), .B1(n_433), .B2(n_434), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_9), .A2(n_41), .B1(n_620), .B2(n_621), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_10), .A2(n_22), .B1(n_457), .B2(n_458), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g1052 ( .A1(n_11), .A2(n_243), .B1(n_453), .B2(n_455), .Y(n_1052) );
AOI21xp33_ASAP7_75t_SL g404 ( .A1(n_12), .A2(n_405), .B(n_407), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_13), .A2(n_120), .B1(n_476), .B2(n_477), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_14), .A2(n_438), .B(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_15), .A2(n_198), .B1(n_488), .B2(n_494), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_16), .A2(n_128), .B1(n_424), .B2(n_425), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_17), .A2(n_463), .B(n_464), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_18), .A2(n_257), .B1(n_379), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_19), .A2(n_292), .B1(n_490), .B2(n_491), .Y(n_489) );
XOR2xp5_ASAP7_75t_L g592 ( .A(n_20), .B(n_593), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_21), .A2(n_148), .B1(n_477), .B2(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_23), .A2(n_152), .B1(n_626), .B2(n_628), .Y(n_625) );
AO22x1_ASAP7_75t_L g731 ( .A1(n_24), .A2(n_31), .B1(n_732), .B2(n_733), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_25), .Y(n_820) );
INVxp33_ASAP7_75t_SL g846 ( .A(n_26), .Y(n_846) );
AO22x2_ASAP7_75t_L g871 ( .A1(n_27), .A2(n_79), .B1(n_822), .B2(n_836), .Y(n_871) );
AO22x1_ASAP7_75t_L g872 ( .A1(n_28), .A2(n_296), .B1(n_851), .B2(n_857), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_29), .A2(n_146), .B1(n_422), .B2(n_424), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_30), .B(n_536), .Y(n_1041) );
INVx1_ASAP7_75t_L g743 ( .A(n_32), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_33), .A2(n_227), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_34), .A2(n_57), .B1(n_540), .B2(n_670), .C(n_671), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_35), .A2(n_86), .B1(n_579), .B2(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g759 ( .A(n_36), .Y(n_759) );
INVx1_ASAP7_75t_L g509 ( .A(n_37), .Y(n_509) );
INVx1_ASAP7_75t_L g672 ( .A(n_38), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_39), .A2(n_129), .B1(n_818), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_40), .A2(n_49), .B1(n_740), .B2(n_741), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_42), .A2(n_284), .B1(n_457), .B2(n_566), .Y(n_1051) );
INVx1_ASAP7_75t_SL g1095 ( .A(n_43), .Y(n_1095) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_44), .B(n_222), .Y(n_306) );
INVx1_ASAP7_75t_L g337 ( .A(n_44), .Y(n_337) );
INVxp67_ASAP7_75t_L g390 ( .A(n_44), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_45), .A2(n_224), .B1(n_381), .B2(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_46), .A2(n_137), .B1(n_463), .B2(n_612), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_47), .A2(n_62), .B1(n_452), .B2(n_453), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_48), .A2(n_231), .B1(n_812), .B2(n_822), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_50), .A2(n_133), .B1(n_851), .B2(n_853), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_51), .A2(n_150), .B1(n_430), .B2(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_52), .B(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_53), .A2(n_64), .B1(n_496), .B2(n_497), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g1050 ( .A1(n_54), .A2(n_78), .B1(n_317), .B2(n_450), .Y(n_1050) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_55), .B(n_322), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_56), .A2(n_116), .B1(n_576), .B2(n_578), .Y(n_575) );
INVx1_ASAP7_75t_SL g1088 ( .A(n_58), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_59), .A2(n_287), .B1(n_379), .B2(n_630), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_60), .A2(n_250), .B1(n_375), .B2(n_424), .Y(n_634) );
INVx1_ASAP7_75t_L g408 ( .A(n_61), .Y(n_408) );
INVx1_ASAP7_75t_L g757 ( .A(n_63), .Y(n_757) );
INVx1_ASAP7_75t_L g783 ( .A(n_65), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_67), .A2(n_276), .B1(n_352), .B2(n_359), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_68), .A2(n_147), .B1(n_457), .B2(n_458), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_69), .A2(n_251), .B1(n_836), .B2(n_864), .Y(n_863) );
INVx1_ASAP7_75t_SL g1093 ( .A(n_70), .Y(n_1093) );
INVx2_ASAP7_75t_L g303 ( .A(n_71), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_72), .A2(n_111), .B1(n_340), .B2(n_449), .Y(n_795) );
INVx1_ASAP7_75t_L g779 ( .A(n_73), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_74), .A2(n_126), .B1(n_365), .B2(n_369), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_75), .A2(n_142), .B1(n_434), .B2(n_449), .Y(n_596) );
INVx1_ASAP7_75t_L g809 ( .A(n_76), .Y(n_809) );
AND2x4_ASAP7_75t_L g815 ( .A(n_76), .B(n_303), .Y(n_815) );
INVx1_ASAP7_75t_SL g852 ( .A(n_76), .Y(n_852) );
INVxp33_ASAP7_75t_SL g823 ( .A(n_77), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g1069 ( .A1(n_80), .A2(n_91), .B1(n_1070), .B2(n_1073), .Y(n_1069) );
INVx1_ASAP7_75t_SL g1091 ( .A(n_81), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_82), .A2(n_103), .B1(n_427), .B2(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g1037 ( .A1(n_83), .A2(n_1038), .B(n_1039), .Y(n_1037) );
INVx1_ASAP7_75t_L g762 ( .A(n_84), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_85), .A2(n_186), .B1(n_519), .B2(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g616 ( .A(n_87), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_88), .A2(n_264), .B1(n_352), .B2(n_359), .Y(n_442) );
INVx1_ASAP7_75t_L g718 ( .A(n_89), .Y(n_718) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_90), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_92), .A2(n_207), .B1(n_359), .B2(n_636), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_93), .A2(n_291), .B1(n_434), .B2(n_525), .Y(n_720) );
INVx1_ASAP7_75t_L g753 ( .A(n_94), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_95), .A2(n_114), .B1(n_1045), .B2(n_1046), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_96), .A2(n_182), .B1(n_317), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_97), .A2(n_254), .B1(n_397), .B2(n_401), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_98), .A2(n_124), .B1(n_493), .B2(n_494), .Y(n_492) );
INVx1_ASAP7_75t_L g323 ( .A(n_99), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_99), .B(n_221), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_100), .A2(n_195), .B1(n_539), .B2(n_541), .Y(n_538) );
OAI22x1_ASAP7_75t_L g446 ( .A1(n_101), .A2(n_447), .B1(n_459), .B2(n_478), .Y(n_446) );
NAND5xp2_ASAP7_75t_SL g447 ( .A(n_101), .B(n_448), .C(n_451), .D(n_454), .E(n_456), .Y(n_447) );
INVx1_ASAP7_75t_L g603 ( .A(n_102), .Y(n_603) );
XNOR2x1_ASAP7_75t_L g645 ( .A(n_104), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_104), .A2(n_161), .B1(n_822), .B2(n_836), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_105), .A2(n_168), .B1(n_397), .B2(n_436), .C(n_439), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_106), .A2(n_160), .B1(n_429), .B2(n_430), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_107), .A2(n_582), .B(n_584), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_108), .B(n_540), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_109), .A2(n_237), .B1(n_352), .B2(n_359), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_110), .A2(n_214), .B1(n_449), .B2(n_450), .Y(n_563) );
INVx2_ASAP7_75t_R g774 ( .A(n_112), .Y(n_774) );
AO221x2_ASAP7_75t_L g804 ( .A1(n_112), .A2(n_113), .B1(n_805), .B2(n_812), .C(n_816), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_115), .B(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_117), .A2(n_169), .B1(n_420), .B2(n_422), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_118), .A2(n_140), .B1(n_544), .B2(n_692), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_119), .A2(n_293), .B1(n_807), .B2(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_121), .A2(n_202), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_123), .A2(n_255), .B1(n_491), .B2(n_493), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g716 ( .A1(n_125), .A2(n_500), .B(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_127), .A2(n_164), .B1(n_612), .B2(n_1098), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_130), .A2(n_201), .B1(n_379), .B2(n_381), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_131), .B(n_574), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_132), .A2(n_196), .B1(n_589), .B2(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_134), .A2(n_158), .B1(n_352), .B2(n_514), .Y(n_513) );
NAND2xp33_ASAP7_75t_L g687 ( .A(n_136), .B(n_434), .Y(n_687) );
INVx1_ASAP7_75t_L g653 ( .A(n_138), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_139), .A2(n_261), .B1(n_449), .B2(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g587 ( .A(n_141), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_143), .A2(n_245), .B1(n_317), .B2(n_455), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_144), .A2(n_159), .B1(n_373), .B2(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_145), .A2(n_211), .B1(n_628), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_149), .A2(n_184), .B1(n_544), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_151), .A2(n_275), .B1(n_429), .B2(n_490), .Y(n_655) );
INVx1_ASAP7_75t_L g465 ( .A(n_153), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_154), .A2(n_191), .B1(n_420), .B2(n_521), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_155), .A2(n_234), .B1(n_427), .B2(n_430), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_156), .A2(n_229), .B1(n_702), .B2(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g751 ( .A(n_157), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g794 ( .A1(n_162), .A2(n_212), .B1(n_455), .B2(n_525), .Y(n_794) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_163), .A2(n_200), .B1(n_543), .B2(n_545), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_165), .A2(n_283), .B1(n_352), .B2(n_702), .Y(n_723) );
INVx1_ASAP7_75t_L g1087 ( .A(n_166), .Y(n_1087) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_167), .A2(n_265), .B1(n_424), .B2(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g778 ( .A(n_170), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_171), .A2(n_282), .B1(n_373), .B2(n_375), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_172), .A2(n_192), .B1(n_630), .B2(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_173), .A2(n_295), .B1(n_477), .B2(n_1043), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_174), .A2(n_258), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g1066 ( .A1(n_175), .A2(n_252), .B1(n_453), .B2(n_1067), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_176), .A2(n_285), .B1(n_373), .B2(n_433), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_177), .A2(n_213), .B1(n_516), .B2(n_517), .Y(n_515) );
XNOR2x1_ASAP7_75t_L g710 ( .A(n_179), .B(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_180), .Y(n_415) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_181), .Y(n_559) );
INVx1_ASAP7_75t_L g784 ( .A(n_183), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_185), .A2(n_233), .B1(n_317), .B2(n_340), .Y(n_316) );
XOR2x2_ASAP7_75t_L g728 ( .A(n_187), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_188), .B(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_189), .A2(n_215), .B1(n_807), .B2(n_818), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_189), .A2(n_1035), .B1(n_1053), .B2(n_1054), .Y(n_1034) );
INVx1_ASAP7_75t_L g1053 ( .A(n_189), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_189), .A2(n_1061), .B1(n_1099), .B2(n_1101), .Y(n_1060) );
INVx1_ASAP7_75t_L g1040 ( .A(n_190), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_193), .A2(n_274), .B1(n_317), .B2(n_455), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_194), .A2(n_236), .B1(n_487), .B2(n_502), .Y(n_648) );
OA22x2_ASAP7_75t_L g327 ( .A1(n_197), .A2(n_222), .B1(n_322), .B2(n_326), .Y(n_327) );
INVx1_ASAP7_75t_L g347 ( .A(n_197), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_199), .A2(n_219), .B1(n_702), .B2(n_703), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_203), .A2(n_240), .B1(n_379), .B2(n_401), .Y(n_613) );
INVx1_ASAP7_75t_L g505 ( .A(n_204), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_205), .A2(n_528), .B(n_531), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_206), .A2(n_267), .B1(n_317), .B2(n_365), .Y(n_665) );
INVx1_ASAP7_75t_L g537 ( .A(n_208), .Y(n_537) );
AOI221x1_ASAP7_75t_L g688 ( .A1(n_209), .A2(n_263), .B1(n_352), .B2(n_433), .C(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g534 ( .A(n_210), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_216), .A2(n_260), .B1(n_457), .B2(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g841 ( .A(n_217), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_218), .A2(n_272), .B1(n_449), .B2(n_740), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_220), .A2(n_230), .B1(n_807), .B2(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g339 ( .A(n_221), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_221), .B(n_345), .Y(n_414) );
OAI21xp33_ASAP7_75t_L g348 ( .A1(n_222), .A2(n_238), .B(n_349), .Y(n_348) );
AO22x2_ASAP7_75t_L g510 ( .A1(n_223), .A2(n_511), .B1(n_547), .B2(n_548), .Y(n_510) );
INVx1_ASAP7_75t_L g548 ( .A(n_223), .Y(n_548) );
AND2x2_ASAP7_75t_L g689 ( .A(n_225), .B(n_421), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_228), .A2(n_262), .B1(n_452), .B2(n_453), .Y(n_798) );
INVx1_ASAP7_75t_SL g1083 ( .A(n_232), .Y(n_1083) );
INVx1_ASAP7_75t_SL g842 ( .A(n_235), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_238), .B(n_278), .Y(n_307) );
INVx1_ASAP7_75t_L g325 ( .A(n_238), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_239), .A2(n_273), .B1(n_496), .B2(n_497), .Y(n_495) );
AOI21xp33_ASAP7_75t_L g601 ( .A1(n_241), .A2(n_574), .B(n_602), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g1080 ( .A(n_242), .Y(n_1080) );
INVx1_ASAP7_75t_L g440 ( .A(n_246), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_247), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_248), .B(n_694), .Y(n_693) );
XNOR2x1_ASAP7_75t_L g416 ( .A(n_249), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g786 ( .A(n_253), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_256), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_259), .A2(n_266), .B1(n_523), .B2(n_524), .Y(n_522) );
XOR2xp5_ASAP7_75t_L g1061 ( .A(n_268), .B(n_1062), .Y(n_1061) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_269), .A2(n_281), .B1(n_365), .B2(n_639), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_270), .B(n_686), .C(n_690), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_270), .A2(n_690), .B1(n_696), .B2(n_1106), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_270), .A2(n_686), .B(n_700), .Y(n_707) );
INVx1_ASAP7_75t_SL g1077 ( .A(n_271), .Y(n_1077) );
INVx1_ASAP7_75t_L g746 ( .A(n_277), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_278), .B(n_332), .Y(n_331) );
AOI21xp33_ASAP7_75t_L g503 ( .A1(n_279), .A2(n_429), .B(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_280), .A2(n_289), .B1(n_365), .B2(n_525), .Y(n_595) );
INVx1_ASAP7_75t_SL g1078 ( .A(n_286), .Y(n_1078) );
INVx1_ASAP7_75t_L g811 ( .A(n_288), .Y(n_811) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_288), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_290), .B(n_472), .Y(n_471) );
XNOR2x1_ASAP7_75t_L g661 ( .A(n_293), .B(n_662), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_309), .B(n_799), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx4_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND3xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .C(n_308), .Y(n_300) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_301), .B(n_1058), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_301), .B(n_1059), .Y(n_1100) );
AOI21xp5_ASAP7_75t_L g1104 ( .A1(n_301), .A2(n_308), .B(n_852), .Y(n_1104) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AO21x1_ASAP7_75t_L g1102 ( .A1(n_302), .A2(n_1103), .B(n_1104), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g808 ( .A(n_303), .B(n_809), .Y(n_808) );
AND3x4_ASAP7_75t_L g851 ( .A(n_303), .B(n_810), .C(n_852), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g1058 ( .A(n_304), .B(n_1059), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AO21x2_ASAP7_75t_L g411 ( .A1(n_305), .A2(n_412), .B(n_413), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g1059 ( .A(n_308), .Y(n_1059) );
XOR2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_554), .Y(n_309) );
OA22x2_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_443), .B1(n_550), .B2(n_551), .Y(n_310) );
INVx1_ASAP7_75t_L g550 ( .A(n_311), .Y(n_550) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
XNOR2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_416), .Y(n_312) );
XNOR2x1_ASAP7_75t_L g313 ( .A(n_314), .B(n_415), .Y(n_313) );
NOR4xp75_ASAP7_75t_L g314 ( .A(n_315), .B(n_363), .C(n_377), .D(n_395), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_351), .Y(n_315) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_318), .Y(n_422) );
BUFx12f_ASAP7_75t_L g525 ( .A(n_318), .Y(n_525) );
BUFx3_ASAP7_75t_L g748 ( .A(n_318), .Y(n_748) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_328), .Y(n_318) );
AND2x2_ASAP7_75t_L g366 ( .A(n_319), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g380 ( .A(n_319), .B(n_357), .Y(n_380) );
AND2x2_ASAP7_75t_L g394 ( .A(n_319), .B(n_361), .Y(n_394) );
AND2x2_ASAP7_75t_L g421 ( .A(n_319), .B(n_367), .Y(n_421) );
AND2x4_ASAP7_75t_L g427 ( .A(n_319), .B(n_357), .Y(n_427) );
AND2x2_ASAP7_75t_L g438 ( .A(n_319), .B(n_361), .Y(n_438) );
AND2x4_ASAP7_75t_L g490 ( .A(n_319), .B(n_367), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_319), .B(n_350), .Y(n_491) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_327), .Y(n_319) );
INVx1_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
NAND2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g326 ( .A(n_322), .Y(n_326) );
INVx3_ASAP7_75t_L g332 ( .A(n_322), .Y(n_332) );
NAND2xp33_ASAP7_75t_L g338 ( .A(n_322), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_322), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_323), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_325), .A2(n_349), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g356 ( .A(n_327), .Y(n_356) );
AND2x2_ASAP7_75t_L g388 ( .A(n_327), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g400 ( .A(n_327), .B(n_355), .Y(n_400) );
AND2x4_ASAP7_75t_L g487 ( .A(n_328), .B(n_354), .Y(n_487) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g350 ( .A(n_329), .Y(n_350) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_334), .Y(n_329) );
AND2x4_ASAP7_75t_L g357 ( .A(n_330), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g362 ( .A(n_330), .Y(n_362) );
AND2x4_ASAP7_75t_L g367 ( .A(n_330), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g384 ( .A(n_330), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_332), .B(n_337), .Y(n_336) );
INVxp67_ASAP7_75t_L g345 ( .A(n_332), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_333), .B(n_344), .C(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g358 ( .A(n_335), .Y(n_358) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx5_ASAP7_75t_L g434 ( .A(n_341), .Y(n_434) );
INVx3_ASAP7_75t_L g633 ( .A(n_341), .Y(n_633) );
INVx2_ASAP7_75t_L g734 ( .A(n_341), .Y(n_734) );
INVx6_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx12f_ASAP7_75t_L g450 ( .A(n_342), .Y(n_450) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_350), .Y(n_342) );
AND2x4_ASAP7_75t_L g371 ( .A(n_343), .B(n_367), .Y(n_371) );
AND2x4_ASAP7_75t_L g403 ( .A(n_343), .B(n_361), .Y(n_403) );
AND2x4_ASAP7_75t_L g430 ( .A(n_343), .B(n_361), .Y(n_430) );
AND2x4_ASAP7_75t_L g488 ( .A(n_343), .B(n_350), .Y(n_488) );
AND2x4_ASAP7_75t_L g494 ( .A(n_343), .B(n_367), .Y(n_494) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_348), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AND2x4_ASAP7_75t_L g376 ( .A(n_350), .B(n_354), .Y(n_376) );
HB1xp67_ASAP7_75t_L g1082 ( .A(n_352), .Y(n_1082) );
BUFx12f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_353), .Y(n_457) );
INVx3_ASAP7_75t_L g637 ( .A(n_353), .Y(n_637) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
AND2x2_ASAP7_75t_L g360 ( .A(n_354), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g374 ( .A(n_354), .B(n_367), .Y(n_374) );
AND2x4_ASAP7_75t_L g493 ( .A(n_354), .B(n_367), .Y(n_493) );
AND2x4_ASAP7_75t_L g496 ( .A(n_354), .B(n_357), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_354), .B(n_361), .Y(n_497) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x4_ASAP7_75t_L g406 ( .A(n_357), .B(n_400), .Y(n_406) );
AND2x4_ASAP7_75t_L g429 ( .A(n_357), .B(n_400), .Y(n_429) );
AND2x4_ASAP7_75t_L g361 ( .A(n_358), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g1084 ( .A(n_359), .Y(n_1084) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx5_ASAP7_75t_L g458 ( .A(n_360), .Y(n_458) );
INVx1_ASAP7_75t_L g568 ( .A(n_360), .Y(n_568) );
BUFx3_ASAP7_75t_L g702 ( .A(n_360), .Y(n_702) );
AND2x4_ASAP7_75t_L g399 ( .A(n_361), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g508 ( .A(n_361), .B(n_400), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_372), .Y(n_363) );
BUFx3_ASAP7_75t_L g523 ( .A(n_365), .Y(n_523) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx8_ASAP7_75t_L g455 ( .A(n_366), .Y(n_455) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_SL g425 ( .A(n_370), .Y(n_425) );
INVx4_ASAP7_75t_L g453 ( .A(n_370), .Y(n_453) );
INVx2_ASAP7_75t_L g521 ( .A(n_370), .Y(n_521) );
INVx4_ASAP7_75t_L g609 ( .A(n_370), .Y(n_609) );
INVx2_ASAP7_75t_L g639 ( .A(n_370), .Y(n_639) );
INVx4_ASAP7_75t_L g703 ( .A(n_370), .Y(n_703) );
INVx1_ASAP7_75t_L g741 ( .A(n_370), .Y(n_741) );
INVx8_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_SL g519 ( .A(n_373), .Y(n_519) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx12f_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_374), .Y(n_452) );
BUFx3_ASAP7_75t_L g516 ( .A(n_375), .Y(n_516) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_376), .Y(n_433) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_376), .Y(n_449) );
BUFx6f_ASAP7_75t_L g1072 ( .A(n_376), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_391), .Y(n_377) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g469 ( .A(n_380), .Y(n_469) );
INVx2_ASAP7_75t_L g580 ( .A(n_380), .Y(n_580) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g470 ( .A(n_382), .Y(n_470) );
INVx2_ASAP7_75t_L g533 ( .A(n_382), .Y(n_533) );
INVx4_ASAP7_75t_L g612 ( .A(n_382), .Y(n_612) );
OAI21xp33_ASAP7_75t_L g1039 ( .A1(n_382), .A2(n_1040), .B(n_1041), .Y(n_1039) );
INVx5_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g586 ( .A(n_383), .Y(n_586) );
BUFx2_ASAP7_75t_L g630 ( .A(n_383), .Y(n_630) );
BUFx4f_ASAP7_75t_L g790 ( .A(n_383), .Y(n_790) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
AND2x2_ASAP7_75t_L g502 ( .A(n_384), .B(n_388), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx1_ASAP7_75t_L g412 ( .A(n_386), .Y(n_412) );
INVx1_ASAP7_75t_L g763 ( .A(n_392), .Y(n_763) );
INVx3_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g620 ( .A(n_393), .Y(n_620) );
INVx2_ASAP7_75t_L g670 ( .A(n_393), .Y(n_670) );
INVx2_ASAP7_75t_L g788 ( .A(n_393), .Y(n_788) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g474 ( .A(n_394), .Y(n_474) );
BUFx3_ASAP7_75t_L g500 ( .A(n_394), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_396), .B(n_404), .Y(n_395) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_SL g476 ( .A(n_398), .Y(n_476) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx8_ASAP7_75t_SL g540 ( .A(n_399), .Y(n_540) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_399), .Y(n_574) );
INVx2_ASAP7_75t_L g624 ( .A(n_399), .Y(n_624) );
BUFx3_ASAP7_75t_L g694 ( .A(n_399), .Y(n_694) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g628 ( .A(n_402), .Y(n_628) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_403), .Y(n_477) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_403), .Y(n_692) );
INVx4_ASAP7_75t_L g752 ( .A(n_405), .Y(n_752) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g463 ( .A(n_406), .Y(n_463) );
BUFx3_ASAP7_75t_L g544 ( .A(n_406), .Y(n_544) );
INVx1_ASAP7_75t_L g627 ( .A(n_406), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx2_ASAP7_75t_L g589 ( .A(n_409), .Y(n_589) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_410), .Y(n_441) );
INVx2_ASAP7_75t_L g605 ( .A(n_410), .Y(n_605) );
INVx1_ASAP7_75t_L g621 ( .A(n_410), .Y(n_621) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_410), .Y(n_1098) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g467 ( .A(n_411), .Y(n_467) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_418), .B(n_431), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_419), .B(n_423), .C(n_426), .D(n_428), .Y(n_418) );
BUFx4f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_421), .Y(n_745) );
BUFx12f_ASAP7_75t_L g740 ( .A(n_424), .Y(n_740) );
INVx1_ASAP7_75t_L g1068 ( .A(n_424), .Y(n_1068) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .C(n_442), .Y(n_431) );
BUFx3_ASAP7_75t_L g732 ( .A(n_433), .Y(n_732) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_441), .B(n_718), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_510), .B2(n_549), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_444), .A2(n_549), .B1(n_552), .B2(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_444), .Y(n_552) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
XNOR2x1_ASAP7_75t_L g445 ( .A(n_446), .B(n_482), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g479 ( .A(n_448), .B(n_451), .C(n_456), .D(n_471), .Y(n_479) );
BUFx3_ASAP7_75t_L g517 ( .A(n_450), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_454), .B(n_475), .Y(n_481) );
BUFx3_ASAP7_75t_L g514 ( .A(n_458), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .C(n_475), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g480 ( .A(n_461), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_468), .Y(n_461) );
INVx2_ASAP7_75t_L g577 ( .A(n_463), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_466), .B(n_653), .Y(n_652) );
INVx4_ASAP7_75t_L g765 ( .A(n_466), .Y(n_765) );
INVx1_ASAP7_75t_L g791 ( .A(n_466), .Y(n_791) );
INVx4_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx3_ASAP7_75t_L g506 ( .A(n_467), .Y(n_506) );
INVx2_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
INVx1_ASAP7_75t_L g1096 ( .A(n_472), .Y(n_1096) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g530 ( .A(n_473), .Y(n_530) );
INVx2_ASAP7_75t_L g600 ( .A(n_473), .Y(n_600) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g699 ( .A(n_474), .Y(n_699) );
INVx2_ASAP7_75t_L g1092 ( .A(n_476), .Y(n_1092) );
BUFx3_ASAP7_75t_L g541 ( .A(n_477), .Y(n_541) );
INVx4_ASAP7_75t_L g760 ( .A(n_477), .Y(n_760) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
XOR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_509), .Y(n_483) );
NOR2xp67_ASAP7_75t_L g484 ( .A(n_485), .B(n_498), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_489), .C(n_492), .D(n_495), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .C(n_503), .D(n_507), .Y(n_498) );
INVx1_ASAP7_75t_L g583 ( .A(n_500), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx4_ASAP7_75t_L g536 ( .A(n_506), .Y(n_536) );
INVx4_ASAP7_75t_L g549 ( .A(n_510), .Y(n_549) );
INVx1_ASAP7_75t_L g547 ( .A(n_511), .Y(n_547) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_512), .B(n_526), .Y(n_511) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .C(n_518), .D(n_522), .Y(n_512) );
BUFx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g1076 ( .A(n_523), .Y(n_1076) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .C(n_542), .Y(n_526) );
INVx2_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_534), .B1(n_535), .B2(n_537), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g553 ( .A(n_549), .Y(n_553) );
XOR2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_680), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_642), .B2(n_643), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OA22x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_591), .B1(n_640), .B2(n_641), .Y(n_557) );
INVx2_ASAP7_75t_L g641 ( .A(n_558), .Y(n_641) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B(n_590), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_559), .B(n_562), .C(n_571), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_570), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND4xp25_ASAP7_75t_SL g562 ( .A(n_563), .B(n_564), .C(n_565), .D(n_569), .Y(n_562) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .C(n_581), .Y(n_571) );
INVx1_ASAP7_75t_L g758 ( .A(n_573), .Y(n_758) );
BUFx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g1045 ( .A(n_577), .Y(n_1045) );
BUFx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g1047 ( .A(n_579), .Y(n_1047) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_580), .Y(n_676) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_587), .B(n_588), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g640 ( .A(n_591), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_614), .Y(n_591) );
NAND4xp75_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .C(n_606), .D(n_610), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
OA21x2_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_601), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_604), .B(n_672), .Y(n_671) );
INVx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
XNOR2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_616), .Y(n_615) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_618), .B(n_631), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .C(n_625), .D(n_629), .Y(n_618) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_624), .A2(n_760), .B1(n_783), .B2(n_784), .Y(n_782) );
INVx2_ASAP7_75t_L g1043 ( .A(n_624), .Y(n_1043) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .C(n_635), .D(n_638), .Y(n_631) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g738 ( .A(n_637), .Y(n_738) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AO22x1_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_659), .B1(n_677), .B2(n_678), .Y(n_643) );
INVx1_ASAP7_75t_L g677 ( .A(n_644), .Y(n_677) );
AO22x2_ASAP7_75t_L g769 ( .A1(n_644), .A2(n_770), .B1(n_772), .B2(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g771 ( .A(n_645), .Y(n_771) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_654), .Y(n_646) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .C(n_650), .D(n_651), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .C(n_657), .D(n_658), .Y(n_654) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g679 ( .A(n_660), .Y(n_679) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_668), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .C(n_666), .D(n_667), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_673), .C(n_674), .Y(n_668) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g755 ( .A(n_676), .Y(n_755) );
INVx2_ASAP7_75t_L g781 ( .A(n_676), .Y(n_781) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_768), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_727), .B1(n_766), .B2(n_767), .Y(n_681) );
INVx1_ASAP7_75t_L g766 ( .A(n_682), .Y(n_766) );
OA22x2_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_708), .B1(n_724), .B2(n_725), .Y(n_682) );
INVx1_ASAP7_75t_L g724 ( .A(n_683), .Y(n_724) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AO21x2_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_695), .B(n_705), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_691), .B(n_693), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_700), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_699), .Y(n_1038) );
NAND2x1_ASAP7_75t_SL g700 ( .A(n_701), .B(n_704), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
BUFx4_ASAP7_75t_SL g726 ( .A(n_710), .Y(n_726) );
NOR2x1_ASAP7_75t_L g711 ( .A(n_712), .B(n_719), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .C(n_715), .D(n_716), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .C(n_722), .D(n_723), .Y(n_719) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g767 ( .A(n_727), .Y(n_767) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_749), .Y(n_729) );
NOR3xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_735), .C(n_742), .Y(n_730) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g1074 ( .A(n_734), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .Y(n_735) );
BUFx4f_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_746), .B2(n_747), .Y(n_742) );
INVxp67_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_747), .A2(n_1076), .B1(n_1077), .B2(n_1078), .Y(n_1075) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NOR3xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_756), .C(n_761), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_752), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_752), .A2(n_1087), .B1(n_1088), .B2(n_1089), .Y(n_1086) );
INVxp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g1090 ( .A1(n_760), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
OAI21xp33_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B(n_764), .Y(n_761) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
XNOR2x1_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
AND2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_792), .Y(n_775) );
NOR3xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_782), .C(n_785), .Y(n_776) );
INVxp67_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g1089 ( .A(n_781), .Y(n_1089) );
OAI21xp33_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B(n_789), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_796), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NAND2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_1032), .B1(n_1034), .B2(n_1055), .C(n_1060), .Y(n_799) );
NOR3xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_954), .C(n_994), .Y(n_800) );
OAI211xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_827), .B(n_894), .C(n_928), .Y(n_801) );
INVxp67_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_824), .Y(n_803) );
INVx2_ASAP7_75t_L g899 ( .A(n_804), .Y(n_899) );
HB1xp67_ASAP7_75t_SL g900 ( .A(n_804), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_804), .B(n_903), .Y(n_947) );
AOI31xp33_ASAP7_75t_L g954 ( .A1(n_804), .A2(n_955), .A3(n_960), .B(n_987), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_804), .B(n_881), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_805), .Y(n_1033) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_806), .A2(n_844), .B1(n_845), .B2(n_846), .Y(n_843) );
INVx3_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AND2x4_ASAP7_75t_L g807 ( .A(n_808), .B(n_810), .Y(n_807) );
AND2x4_ASAP7_75t_L g818 ( .A(n_808), .B(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g853 ( .A(n_808), .B(n_819), .Y(n_853) );
AND2x2_ASAP7_75t_L g857 ( .A(n_808), .B(n_819), .Y(n_857) );
AND2x4_ASAP7_75t_L g814 ( .A(n_810), .B(n_815), .Y(n_814) );
AND2x4_ASAP7_75t_L g836 ( .A(n_810), .B(n_815), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_810), .B(n_815), .Y(n_845) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
AND2x4_ASAP7_75t_L g822 ( .A(n_815), .B(n_819), .Y(n_822) );
AND2x2_ASAP7_75t_L g834 ( .A(n_815), .B(n_819), .Y(n_834) );
AND2x2_ASAP7_75t_L g864 ( .A(n_815), .B(n_819), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_820), .B1(n_821), .B2(n_823), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_817), .A2(n_821), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx3_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx3_ASAP7_75t_L g904 ( .A(n_824), .Y(n_904) );
OR2x2_ASAP7_75t_L g927 ( .A(n_824), .B(n_869), .Y(n_927) );
AND2x2_ASAP7_75t_L g969 ( .A(n_824), .B(n_944), .Y(n_969) );
OR2x2_ASAP7_75t_L g999 ( .A(n_824), .B(n_1000), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
AOI221xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_859), .B1(n_866), .B2(n_873), .C(n_874), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_837), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_830), .B(n_848), .Y(n_873) );
AND2x2_ASAP7_75t_L g892 ( .A(n_830), .B(n_893), .Y(n_892) );
AND2x2_ASAP7_75t_L g908 ( .A(n_830), .B(n_848), .Y(n_908) );
AND2x2_ASAP7_75t_L g921 ( .A(n_830), .B(n_898), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_830), .B(n_855), .Y(n_978) );
NOR3xp33_ASAP7_75t_L g1030 ( .A(n_830), .B(n_931), .C(n_1007), .Y(n_1030) );
INVx3_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx3_ASAP7_75t_L g877 ( .A(n_832), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_832), .B(n_867), .Y(n_890) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_832), .B(n_855), .Y(n_1027) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_847), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g880 ( .A(n_838), .B(n_881), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_838), .B(n_897), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_838), .B(n_903), .Y(n_911) );
INVx1_ASAP7_75t_L g922 ( .A(n_838), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_838), .B(n_942), .Y(n_976) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx3_ASAP7_75t_L g867 ( .A(n_839), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_839), .B(n_862), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_839), .B(n_877), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_839), .B(n_870), .Y(n_964) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_839), .Y(n_1002) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_839), .B(n_862), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_839), .B(n_861), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_839), .B(n_905), .Y(n_1028) );
OR2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .Y(n_839) );
INVx1_ASAP7_75t_L g888 ( .A(n_847), .Y(n_888) );
OAI221xp5_ASAP7_75t_SL g901 ( .A1(n_847), .A2(n_902), .B1(n_906), .B2(n_907), .C(n_909), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_847), .B(n_918), .Y(n_1003) );
OR2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_855), .Y(n_847) );
AND2x2_ASAP7_75t_L g893 ( .A(n_848), .B(n_855), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_848), .B(n_877), .Y(n_943) );
OR2x2_ASAP7_75t_L g986 ( .A(n_848), .B(n_877), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_848), .B(n_1011), .Y(n_1010) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_849), .Y(n_848) );
OR2x2_ASAP7_75t_L g876 ( .A(n_849), .B(n_855), .Y(n_876) );
AND2x2_ASAP7_75t_L g898 ( .A(n_849), .B(n_855), .Y(n_898) );
AND2x2_ASAP7_75t_L g849 ( .A(n_850), .B(n_854), .Y(n_849) );
AOI322xp5_ASAP7_75t_L g909 ( .A1(n_855), .A2(n_882), .A3(n_903), .B1(n_910), .B2(n_912), .C1(n_913), .C2(n_916), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_855), .B(n_877), .Y(n_932) );
INVx1_ASAP7_75t_L g937 ( .A(n_855), .Y(n_937) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_858), .Y(n_855) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g912 ( .A(n_860), .Y(n_912) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AND2x2_ASAP7_75t_L g879 ( .A(n_861), .B(n_870), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
OR2x2_ASAP7_75t_L g869 ( .A(n_862), .B(n_870), .Y(n_869) );
BUFx2_ASAP7_75t_L g883 ( .A(n_862), .Y(n_883) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_862), .Y(n_885) );
AND2x2_ASAP7_75t_L g905 ( .A(n_862), .B(n_870), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_862), .B(n_934), .Y(n_933) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_862), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_862), .B(n_867), .Y(n_984) );
AND2x4_ASAP7_75t_L g862 ( .A(n_863), .B(n_865), .Y(n_862) );
AND2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx1_ASAP7_75t_SL g931 ( .A(n_867), .Y(n_931) );
AND2x2_ASAP7_75t_L g959 ( .A(n_867), .B(n_893), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_868), .A2(n_920), .B1(n_924), .B2(n_927), .Y(n_919) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_868), .A2(n_956), .B(n_957), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g979 ( .A(n_868), .B(n_892), .Y(n_979) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
CKINVDCx6p67_ASAP7_75t_R g882 ( .A(n_870), .Y(n_882) );
AOI321xp33_ASAP7_75t_L g894 ( .A1(n_870), .A2(n_895), .A3(n_899), .B1(n_900), .B2(n_901), .C(n_919), .Y(n_894) );
OR2x2_ASAP7_75t_L g934 ( .A(n_870), .B(n_904), .Y(n_934) );
INVx1_ASAP7_75t_L g945 ( .A(n_870), .Y(n_945) );
OR2x6_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
OAI221xp5_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_877), .B1(n_878), .B2(n_880), .C(n_884), .Y(n_874) );
INVx1_ASAP7_75t_L g972 ( .A(n_875), .Y(n_972) );
OR2x2_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_876), .B(n_890), .Y(n_939) );
INVx1_ASAP7_75t_L g951 ( .A(n_876), .Y(n_951) );
NOR2xp33_ASAP7_75t_L g1001 ( .A(n_876), .B(n_1002), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_876), .B(n_914), .Y(n_1031) );
AND2x2_ASAP7_75t_L g897 ( .A(n_877), .B(n_898), .Y(n_897) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_877), .Y(n_926) );
AND2x2_ASAP7_75t_L g950 ( .A(n_877), .B(n_951), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_877), .B(n_959), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_877), .B(n_888), .Y(n_989) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_879), .B(n_903), .Y(n_906) );
AOI32xp33_ASAP7_75t_L g1029 ( .A1(n_879), .A2(n_910), .A3(n_985), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_881), .B(n_931), .Y(n_936) );
INVx1_ASAP7_75t_L g940 ( .A(n_881), .Y(n_940) );
AND2x2_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_882), .B(n_904), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_883), .B(n_958), .Y(n_957) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_883), .B(n_904), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_891), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
AND2x2_ASAP7_75t_L g996 ( .A(n_892), .B(n_983), .Y(n_996) );
AND2x2_ASAP7_75t_L g916 ( .A(n_893), .B(n_917), .Y(n_916) );
AND2x2_ASAP7_75t_L g925 ( .A(n_893), .B(n_926), .Y(n_925) );
AOI211xp5_ASAP7_75t_L g960 ( .A1(n_893), .A2(n_961), .B(n_962), .C(n_973), .Y(n_960) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g1022 ( .A(n_897), .Y(n_1022) );
INVx1_ASAP7_75t_L g914 ( .A(n_898), .Y(n_914) );
AND2x2_ASAP7_75t_L g956 ( .A(n_898), .B(n_917), .Y(n_956) );
INVx1_ASAP7_75t_L g923 ( .A(n_899), .Y(n_923) );
INVxp67_ASAP7_75t_L g1015 ( .A(n_900), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
INVx5_ASAP7_75t_L g953 ( .A(n_903), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_903), .B(n_971), .Y(n_993) );
NOR3xp33_ASAP7_75t_L g1013 ( .A(n_903), .B(n_914), .C(n_1014), .Y(n_1013) );
INVx3_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_904), .B(n_944), .Y(n_1008) );
INVx2_ASAP7_75t_L g1000 ( .A(n_905), .Y(n_1000) );
INVx1_ASAP7_75t_L g961 ( .A(n_906), .Y(n_961) );
CKINVDCx16_ASAP7_75t_R g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
A2O1A1Ixp33_ASAP7_75t_SL g995 ( .A1(n_912), .A2(n_944), .B(n_988), .C(n_996), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
INVx1_ASAP7_75t_L g952 ( .A(n_915), .Y(n_952) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_916), .B(n_971), .Y(n_1025) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
NAND3xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .C(n_923), .Y(n_920) );
INVx1_ASAP7_75t_L g967 ( .A(n_921), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_922), .B(n_972), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_924), .B(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
AOI221xp5_ASAP7_75t_L g928 ( .A1(n_929), .A2(n_933), .B1(n_935), .B2(n_946), .C(n_948), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_931), .B(n_942), .Y(n_941) );
OAI211xp5_ASAP7_75t_L g973 ( .A1(n_934), .A2(n_974), .B(n_979), .C(n_980), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_934), .A2(n_941), .B1(n_999), .B2(n_1024), .Y(n_1023) );
OAI222xp33_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_938), .B2(n_940), .C1(n_941), .C2(n_944), .Y(n_935) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_944), .B(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVxp67_ASAP7_75t_SL g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_952), .C(n_953), .Y(n_949) );
OAI22xp33_ASAP7_75t_L g962 ( .A1(n_963), .A2(n_965), .B1(n_968), .B2(n_970), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
OAI221xp5_ASAP7_75t_L g1006 ( .A1(n_967), .A2(n_1007), .B1(n_1009), .B2(n_1010), .C(n_1012), .Y(n_1006) );
A2O1A1Ixp33_ASAP7_75t_L g1026 ( .A1(n_967), .A2(n_1027), .B(n_1028), .C(n_1029), .Y(n_1026) );
A2O1A1Ixp33_ASAP7_75t_L g1017 ( .A1(n_968), .A2(n_993), .B(n_1018), .C(n_1019), .Y(n_1017) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_972), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_971), .B(n_978), .Y(n_977) );
NOR2xp33_ASAP7_75t_L g974 ( .A(n_975), .B(n_977), .Y(n_974) );
INVxp33_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVxp67_ASAP7_75t_SL g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_983), .B(n_985), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
OAI21xp33_ASAP7_75t_L g987 ( .A1(n_988), .A2(n_990), .B(n_992), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
A2O1A1Ixp33_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_997), .B(n_1015), .C(n_1016), .Y(n_994) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_1001), .B1(n_1003), .B2(n_1004), .C(n_1006), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1003), .Y(n_1018) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
NOR3xp33_ASAP7_75t_SL g1016 ( .A(n_1017), .B(n_1023), .C(n_1026), .Y(n_1016) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
NOR2xp33_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1022), .Y(n_1020) );
INVxp67_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g1032 ( .A(n_1033), .Y(n_1032) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1035), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1048), .Y(n_1035) );
NAND3xp33_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1042), .C(n_1044), .Y(n_1036) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
NAND4xp25_ASAP7_75t_SL g1048 ( .A(n_1049), .B(n_1050), .C(n_1051), .D(n_1052), .Y(n_1048) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
NAND2xp5_ASAP7_75t_SL g1063 ( .A(n_1064), .B(n_1085), .Y(n_1063) );
NOR3xp33_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1075), .C(n_1079), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1069), .Y(n_1065) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
OAI22x1_ASAP7_75t_SL g1079 ( .A1(n_1080), .A2(n_1081), .B1(n_1083), .B2(n_1084), .Y(n_1079) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
NOR3xp33_ASAP7_75t_SL g1085 ( .A(n_1086), .B(n_1090), .C(n_1094), .Y(n_1085) );
OAI21xp33_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1096), .B(n_1097), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
endmodule