module fake_jpeg_12306_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_23),
.B(n_9),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_19),
.B(n_0),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_66),
.B(n_35),
.C(n_38),
.Y(n_118)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_23),
.B(n_9),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_39),
.B1(n_36),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_83),
.B1(n_90),
.B2(n_110),
.Y(n_127)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_30),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_81),
.B(n_82),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_30),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_43),
.B1(n_27),
.B2(n_22),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_85),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_47),
.B(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_92),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_43),
.B1(n_27),
.B2(n_22),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_31),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_26),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_37),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

CKINVDCx12_ASAP7_75t_R g102 ( 
.A(n_65),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_22),
.B1(n_27),
.B2(n_36),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_103),
.A2(n_107),
.B1(n_93),
.B2(n_99),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_18),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_118),
.C(n_41),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_42),
.B1(n_25),
.B2(n_31),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_52),
.B1(n_50),
.B2(n_49),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_119),
.A2(n_122),
.B1(n_125),
.B2(n_136),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_38),
.B1(n_17),
.B2(n_25),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_17),
.B1(n_42),
.B2(n_36),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_114),
.B1(n_88),
.B2(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_33),
.B1(n_19),
.B2(n_37),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_46),
.B1(n_33),
.B2(n_19),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_76),
.A2(n_34),
.B1(n_111),
.B2(n_74),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_152),
.B1(n_109),
.B2(n_113),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_77),
.A2(n_41),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_41),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_8),
.B1(n_14),
.B2(n_15),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_144),
.Y(n_164)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_145),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_1),
.Y(n_144)
);

AO22x2_ASAP7_75t_L g146 ( 
.A1(n_80),
.A2(n_2),
.B1(n_3),
.B2(n_16),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_146),
.B(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_2),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_106),
.B1(n_115),
.B2(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_153),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_3),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_87),
.B(n_5),
.C(n_7),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_7),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_112),
.B(n_78),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_160),
.A2(n_183),
.B(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_169),
.B1(n_189),
.B2(n_191),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_179),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_166),
.A2(n_176),
.B1(n_177),
.B2(n_175),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_91),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_168),
.B(n_173),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_115),
.B1(n_106),
.B2(n_91),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_113),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_119),
.A2(n_113),
.B1(n_112),
.B2(n_13),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_7),
.B1(n_8),
.B2(n_13),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_14),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_184),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_129),
.B(n_16),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_127),
.A2(n_136),
.B1(n_147),
.B2(n_145),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_193),
.B1(n_178),
.B2(n_169),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_146),
.B(n_133),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_142),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_156),
.B(n_148),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_193),
.B(n_191),
.C(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_146),
.B(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_174),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_138),
.A2(n_152),
.B1(n_154),
.B2(n_135),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_123),
.B1(n_131),
.B2(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_123),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_196),
.B(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_132),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_181),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_188),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_204),
.B(n_208),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_184),
.B1(n_183),
.B2(n_174),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_212),
.B1(n_192),
.B2(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_171),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_209),
.B(n_213),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_164),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_211),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_164),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_183),
.A2(n_163),
.B1(n_159),
.B2(n_194),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_185),
.C(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_217),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_218),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

INVx2_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_220),
.Y(n_247)
);

AND2x4_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_223),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_200),
.B1(n_222),
.B2(n_217),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_199),
.B(n_201),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_161),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_245),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_234),
.B1(n_235),
.B2(n_238),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_213),
.B(n_209),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_230),
.A2(n_240),
.B(n_250),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_220),
.B1(n_221),
.B2(n_207),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_207),
.A2(n_198),
.B(n_215),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_236),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_211),
.B1(n_210),
.B2(n_203),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_218),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_241),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_199),
.A2(n_195),
.B1(n_208),
.B2(n_226),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_196),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_240),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_195),
.B(n_214),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_200),
.A2(n_212),
.B1(n_205),
.B2(n_209),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_247),
.B(n_252),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_219),
.C(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_254),
.C(n_255),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_237),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_235),
.A2(n_251),
.B1(n_229),
.B2(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_269),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_261),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_239),
.C(n_246),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_266),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_242),
.C(n_250),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_267),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_239),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_248),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_233),
.Y(n_281)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_241),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_228),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_234),
.B1(n_251),
.B2(n_231),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_234),
.B1(n_247),
.B2(n_232),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_254),
.B(n_244),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_265),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_233),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_288),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_256),
.A2(n_232),
.B1(n_228),
.B2(n_227),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_260),
.B1(n_258),
.B2(n_256),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_263),
.C(n_255),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_284),
.C(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_257),
.B1(n_270),
.B2(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_298),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_270),
.B1(n_267),
.B2(n_274),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_253),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_293),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_273),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_305),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_287),
.B1(n_289),
.B2(n_228),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_258),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_310),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_296),
.A2(n_275),
.B(n_282),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_282),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_297),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_277),
.B1(n_284),
.B2(n_283),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_297),
.C(n_303),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_228),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_323),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_307),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_316),
.B(n_298),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_308),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_299),
.B1(n_304),
.B2(n_272),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_295),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_326),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_317),
.A2(n_299),
.B1(n_313),
.B2(n_310),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_320),
.C(n_322),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_330),
.B1(n_320),
.B2(n_315),
.Y(n_334)
);

NOR2x1_ASAP7_75t_SL g330 ( 
.A(n_321),
.B(n_311),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_327),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_290),
.B(n_326),
.C(n_227),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_331),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_336),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_290),
.C(n_325),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_307),
.Y(n_341)
);


endmodule