module fake_jpeg_18254_n_225 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_225);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_14;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_29),
.Y(n_32)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_27),
.B1(n_26),
.B2(n_28),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_39),
.A2(n_40),
.B1(n_52),
.B2(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_27),
.B1(n_26),
.B2(n_13),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_13),
.B1(n_28),
.B2(n_16),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_29),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_27),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_26),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_28),
.B1(n_22),
.B2(n_30),
.Y(n_52)
);

OA21x2_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_22),
.B(n_33),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_56),
.B(n_48),
.C(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_33),
.B(n_36),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_31),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_67),
.Y(n_73)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_74),
.Y(n_84)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_61),
.B(n_53),
.Y(n_95)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_79),
.Y(n_85)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_67),
.B1(n_54),
.B2(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_88),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_77),
.B1(n_72),
.B2(n_70),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_64),
.C(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_60),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_61),
.B1(n_63),
.B2(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_47),
.B(n_52),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_66),
.B(n_60),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_23),
.B(n_41),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_64),
.B1(n_42),
.B2(n_44),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_105),
.B1(n_115),
.B2(n_106),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_58),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_107),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_39),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_113),
.B(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_16),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_111),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_87),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_71),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_40),
.C(n_12),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_12),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_31),
.A3(n_28),
.B1(n_38),
.B2(n_23),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_69),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_89),
.B1(n_99),
.B2(n_86),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_141),
.B1(n_135),
.B2(n_136),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_89),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_102),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_99),
.C(n_65),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_31),
.C(n_34),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_89),
.B1(n_62),
.B2(n_38),
.Y(n_128)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_112),
.B(n_19),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_138),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_113),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_62),
.B1(n_38),
.B2(n_36),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_51),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_120),
.B(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_51),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_30),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_134),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_129),
.B1(n_130),
.B2(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_148),
.C(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_31),
.C(n_34),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_109),
.B(n_11),
.C(n_14),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_154),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_122),
.B1(n_139),
.B2(n_157),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_11),
.C(n_14),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_155),
.C(n_6),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_30),
.C(n_24),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_30),
.C(n_24),
.Y(n_154)
);

XOR2x1_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_19),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_9),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_24),
.C(n_20),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_163),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_140),
.B1(n_123),
.B2(n_128),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_167),
.B(n_173),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_140),
.B1(n_123),
.B2(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_129),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_11),
.B1(n_14),
.B2(n_18),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_147),
.C(n_148),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_25),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_25),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_146),
.B1(n_131),
.B2(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_171),
.B1(n_18),
.B2(n_2),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_154),
.B(n_152),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_173),
.C(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_161),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_192),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_169),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_190),
.B1(n_184),
.B2(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_24),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_180),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_195),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_18),
.B(n_25),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_182),
.B(n_183),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_19),
.C(n_1),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_177),
.B1(n_175),
.B2(n_3),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_202),
.B1(n_6),
.B2(n_2),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_204),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_17),
.C(n_15),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_191),
.B(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_206),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_17),
.C(n_15),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_25),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_17),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_3),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_200),
.A3(n_17),
.B1(n_15),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_15),
.C(n_2),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_216),
.B(n_208),
.Y(n_217)
);

AOI31xp33_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_212),
.A3(n_214),
.B(n_215),
.Y(n_219)
);

OAI321xp33_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_220),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_3),
.C(n_4),
.Y(n_220)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_8),
.B(n_9),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_8),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_8),
.B(n_0),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_0),
.B(n_221),
.Y(n_225)
);


endmodule