module fake_jpeg_25820_n_75 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_75);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_38;
wire n_36;
wire n_74;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_32),
.Y(n_45)
);

CKINVDCx12_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_4),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_12),
.B(n_27),
.C(n_26),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_42),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_41),
.B1(n_34),
.B2(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_30),
.B(n_3),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_48),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_32),
.B1(n_30),
.B2(n_34),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_61)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_17),
.B1(n_28),
.B2(n_23),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_5),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_34),
.B1(n_8),
.B2(n_7),
.Y(n_57)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.C(n_61),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_16),
.A3(n_21),
.B1(n_9),
.B2(n_10),
.Y(n_60)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_64),
.C(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_64),
.B1(n_61),
.B2(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_70),
.B1(n_51),
.B2(n_65),
.Y(n_71)
);

AOI322xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_63),
.A3(n_51),
.B1(n_59),
.B2(n_49),
.C1(n_58),
.C2(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_51),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_68),
.C(n_55),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_43),
.C(n_20),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_22),
.Y(n_75)
);


endmodule