module fake_jpeg_11431_n_178 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_85),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_91),
.Y(n_102)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_0),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_1),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_0),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_63),
.B1(n_88),
.B2(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_71),
.B1(n_80),
.B2(n_75),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_66),
.B1(n_63),
.B2(n_73),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_96),
.B1(n_65),
.B2(n_64),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_66),
.B1(n_76),
.B2(n_59),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_106),
.Y(n_125)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_105),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_58),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_113),
.B1(n_8),
.B2(n_9),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_6),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_80),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_118),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_61),
.B1(n_57),
.B2(n_60),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_69),
.B1(n_74),
.B2(n_72),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_7),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_54),
.B1(n_70),
.B2(n_67),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_123),
.B1(n_126),
.B2(n_23),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_79),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_122),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_24),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_21),
.B1(n_50),
.B2(n_47),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_19),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_8),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_20),
.C(n_46),
.Y(n_128)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_132),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_145),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_15),
.B(n_45),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_140),
.B(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_52),
.C(n_44),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_125),
.B1(n_12),
.B2(n_13),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_146),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_139),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_11),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_160),
.B1(n_134),
.B2(n_138),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_156),
.Y(n_167)
);

AO22x1_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_42),
.B1(n_25),
.B2(n_30),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_158),
.A2(n_131),
.B1(n_132),
.B2(n_128),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_11),
.B(n_12),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_14),
.A3(n_40),
.B1(n_135),
.B2(n_138),
.C1(n_156),
.C2(n_154),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_13),
.B1(n_14),
.B2(n_31),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_157),
.A2(n_137),
.B1(n_141),
.B2(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_162),
.B(n_164),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_166),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_155),
.C(n_165),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_172),
.B1(n_165),
.B2(n_153),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_167),
.B(n_152),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_153),
.B(n_161),
.C(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_151),
.B(n_170),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_163),
.Y(n_178)
);


endmodule