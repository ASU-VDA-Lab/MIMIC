module fake_ibex_2016_n_1007 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1007);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1007;

wire n_599;
wire n_822;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_375;
wire n_317;
wire n_340;
wire n_280;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_470;
wire n_276;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_999;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_472;
wire n_209;
wire n_229;
wire n_589;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_562;
wire n_564;
wire n_506;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_285;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_912;
wire n_890;
wire n_921;
wire n_874;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_503;
wire n_241;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_298;
wire n_202;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

BUFx10_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_33),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_64),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_54),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_71),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_68),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_109),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_43),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_38),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_85),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_17),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_29),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_112),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_22),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_100),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_105),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_15),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_51),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_31),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_80),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_36),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_69),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_110),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_20),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_157),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_89),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_158),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_161),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_145),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_159),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_76),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_25),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_179),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_104),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_41),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_98),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_24),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_L g241 ( 
.A(n_155),
.B(n_139),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_94),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_133),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_46),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_18),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_63),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_174),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_5),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_101),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_90),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_102),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_34),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_52),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_26),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_35),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_21),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_27),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_140),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_82),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_13),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_26),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_97),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_25),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_24),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_138),
.B(n_37),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_11),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_153),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_66),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_31),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_70),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_180),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_72),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_121),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_125),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_150),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_81),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_107),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_154),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_143),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_108),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_6),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_23),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_165),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_47),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_135),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_113),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_166),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_78),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_137),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_33),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_127),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_84),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_144),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_141),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_115),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_6),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_146),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_3),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_168),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_40),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_200),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_200),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_210),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_210),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_200),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_224),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_192),
.B(n_0),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g311 ( 
.A1(n_224),
.A2(n_83),
.B(n_182),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g312 ( 
.A(n_184),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_206),
.B(n_0),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_192),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_272),
.A2(n_77),
.B(n_178),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_208),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_219),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_263),
.B(n_1),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_219),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_273),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_263),
.B(n_1),
.Y(n_324)
);

CKINVDCx6p67_ASAP7_75t_R g325 ( 
.A(n_207),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_215),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_2),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_184),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_219),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_219),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_208),
.B(n_2),
.Y(n_332)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_209),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_217),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_265),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_248),
.B(n_4),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_256),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_236),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_209),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_282),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_186),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

OAI21x1_ASAP7_75t_L g343 ( 
.A1(n_287),
.A2(n_86),
.B(n_175),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_232),
.B(n_7),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_249),
.B(n_8),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_217),
.B(n_9),
.Y(n_346)
);

AOI22x1_ASAP7_75t_SL g347 ( 
.A1(n_239),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_269),
.B(n_10),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_216),
.Y(n_349)
);

BUFx12f_ASAP7_75t_L g350 ( 
.A(n_277),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_R g351 ( 
.A1(n_204),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_234),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_287),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_245),
.Y(n_354)
);

OAI21x1_ASAP7_75t_L g355 ( 
.A1(n_299),
.A2(n_87),
.B(n_173),
.Y(n_355)
);

BUFx8_ASAP7_75t_SL g356 ( 
.A(n_258),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_236),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_252),
.B(n_12),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_264),
.B(n_14),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_236),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_270),
.Y(n_361)
);

BUFx12f_ASAP7_75t_L g362 ( 
.A(n_187),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_292),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_214),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_269),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_295),
.B(n_15),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_295),
.B(n_16),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_185),
.A2(n_88),
.B(n_167),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_189),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_190),
.B(n_16),
.Y(n_371)
);

BUFx8_ASAP7_75t_SL g372 ( 
.A(n_191),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_196),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_197),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_198),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_199),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_188),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_201),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_236),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_238),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_305),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_326),
.B(n_205),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_307),
.Y(n_384)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_305),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_306),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_314),
.B(n_278),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_339),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_307),
.Y(n_390)
);

AND3x2_ASAP7_75t_L g391 ( 
.A(n_322),
.B(n_212),
.C(n_211),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_307),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_307),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_278),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_266),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_306),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_309),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

CKINVDCx6p67_ASAP7_75t_R g401 ( 
.A(n_325),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_225),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_222),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_318),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_310),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_240),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_323),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_310),
.B(n_254),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_310),
.A2(n_250),
.B1(n_213),
.B2(n_242),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_344),
.B(n_193),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_332),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

AO21x2_ASAP7_75t_L g426 ( 
.A1(n_343),
.A2(n_228),
.B(n_223),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_334),
.Y(n_427)
);

NOR2x1p5_ASAP7_75t_L g428 ( 
.A(n_312),
.B(n_262),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_328),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_364),
.B(n_267),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_303),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_328),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_341),
.B(n_283),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_349),
.B(n_284),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_342),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_346),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_376),
.B(n_300),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_304),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_304),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_346),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_312),
.B(n_230),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_304),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_308),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_345),
.B(n_194),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_376),
.B(n_244),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_308),
.Y(n_452)
);

AND3x2_ASAP7_75t_L g453 ( 
.A(n_351),
.B(n_253),
.C(n_246),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_319),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_358),
.B(n_302),
.C(n_257),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_319),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_321),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_366),
.B(n_370),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_321),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_320),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_352),
.B(n_298),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_357),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_345),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_345),
.B(n_195),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_357),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_348),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_362),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_365),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_348),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_357),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_367),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_372),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_366),
.B(n_202),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_360),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_360),
.Y(n_479)
);

CKINVDCx6p67_ASAP7_75t_R g480 ( 
.A(n_329),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_371),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_371),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_333),
.B(n_259),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_354),
.B(n_203),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_360),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_368),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_438),
.B(n_221),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_333),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_388),
.B(n_324),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

INVx8_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_412),
.Y(n_492)
);

OAI22x1_ASAP7_75t_SL g493 ( 
.A1(n_475),
.A2(n_356),
.B1(n_351),
.B2(n_347),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_486),
.A2(n_368),
.B1(n_336),
.B2(n_327),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_350),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_416),
.B(n_350),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_412),
.B(n_336),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_480),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_427),
.Y(n_499)
);

A2O1A1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_476),
.A2(n_482),
.B(n_481),
.C(n_486),
.Y(n_500)
);

NOR2x1p5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_401),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_361),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_389),
.B(n_313),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_420),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_389),
.B(n_370),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_373),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_420),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_470),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_470),
.Y(n_509)
);

OR2x4_ASAP7_75t_L g510 ( 
.A(n_444),
.B(n_337),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_471),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_383),
.B(n_373),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_438),
.B(n_336),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_405),
.B(n_440),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g515 ( 
.A(n_404),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_435),
.B(n_374),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_424),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_463),
.B(n_359),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_405),
.B(n_374),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_316),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_436),
.B(n_316),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_381),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_436),
.B(n_316),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_418),
.B(n_218),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_432),
.B(n_340),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_382),
.Y(n_526)
);

OR2x6_ASAP7_75t_L g527 ( 
.A(n_410),
.B(n_343),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_418),
.B(n_220),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_394),
.B(n_226),
.Y(n_529)
);

NOR3xp33_ASAP7_75t_L g530 ( 
.A(n_419),
.B(n_289),
.C(n_274),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_382),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_410),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_381),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_447),
.B(n_17),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_421),
.B(n_233),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_451),
.B(n_227),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_465),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_472),
.B(n_229),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_451),
.B(n_231),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_481),
.B(n_311),
.C(n_315),
.Y(n_541)
);

NOR2x1p5_ASAP7_75t_L g542 ( 
.A(n_401),
.B(n_475),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_469),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_395),
.B(n_235),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_386),
.Y(n_546)
);

NOR2xp67_ASAP7_75t_L g547 ( 
.A(n_457),
.B(n_18),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_386),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_387),
.Y(n_550)
);

NAND3xp33_ASAP7_75t_L g551 ( 
.A(n_457),
.B(n_311),
.C(n_315),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_387),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_472),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_397),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_397),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_450),
.B(n_294),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_398),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_469),
.B(n_356),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_399),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_466),
.B(n_301),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_431),
.B(n_355),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_391),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_431),
.B(n_237),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_399),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_402),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_402),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_443),
.B(n_243),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_483),
.B(n_247),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_403),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_419),
.B(n_19),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_443),
.B(n_445),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_443),
.B(n_445),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_445),
.B(n_251),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_428),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_395),
.B(n_255),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_468),
.B(n_260),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_408),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_409),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_562),
.A2(n_474),
.B(n_426),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_541),
.A2(n_551),
.B(n_562),
.Y(n_581)
);

NOR3xp33_ASAP7_75t_L g582 ( 
.A(n_495),
.B(n_408),
.C(n_477),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_578),
.B(n_460),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_518),
.B(n_409),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_490),
.B(n_492),
.Y(n_585)
);

O2A1O1Ixp33_ASAP7_75t_L g586 ( 
.A1(n_543),
.A2(n_439),
.B(n_437),
.C(n_434),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_525),
.A2(n_453),
.B1(n_417),
.B2(n_449),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_489),
.B(n_514),
.Y(n_588)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_500),
.A2(n_572),
.B(n_573),
.C(n_503),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_501),
.B(n_456),
.Y(n_590)
);

O2A1O1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_519),
.A2(n_439),
.B(n_455),
.C(n_417),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_516),
.B(n_422),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_516),
.B(n_422),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_491),
.B(n_430),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_515),
.B(n_385),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_498),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_491),
.B(n_430),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_487),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_541),
.A2(n_426),
.B(n_369),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_491),
.B(n_434),
.Y(n_600)
);

OA22x2_ASAP7_75t_L g601 ( 
.A1(n_544),
.A2(n_437),
.B1(n_449),
.B2(n_455),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_551),
.A2(n_369),
.B(n_433),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_544),
.B(n_20),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_532),
.B(n_21),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_559),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_530),
.A2(n_385),
.B1(n_288),
.B2(n_268),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_572),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_573),
.A2(n_497),
.B(n_564),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_502),
.B(n_385),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_490),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_506),
.B(n_385),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_558),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_492),
.B(n_271),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_512),
.B(n_276),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_SL g615 ( 
.A1(n_568),
.A2(n_577),
.B(n_574),
.C(n_529),
.Y(n_615)
);

O2A1O1Ixp5_ASAP7_75t_L g616 ( 
.A1(n_513),
.A2(n_406),
.B(n_384),
.C(n_390),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_487),
.A2(n_291),
.B1(n_293),
.B2(n_280),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_488),
.B(n_281),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_494),
.B(n_286),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_492),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_571),
.A2(n_296),
.B1(n_297),
.B2(n_241),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_504),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_522),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_496),
.B(n_22),
.Y(n_624)
);

BUFx4f_ASAP7_75t_L g625 ( 
.A(n_563),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_527),
.A2(n_485),
.B(n_479),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_527),
.A2(n_478),
.B(n_473),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_507),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_575),
.B(n_23),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_536),
.B(n_27),
.Y(n_630)
);

OAI21xp33_ASAP7_75t_L g631 ( 
.A1(n_524),
.A2(n_528),
.B(n_545),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_517),
.A2(n_441),
.B(n_464),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_540),
.B(n_520),
.Y(n_633)
);

OAI21xp33_ASAP7_75t_L g634 ( 
.A1(n_576),
.A2(n_569),
.B(n_523),
.Y(n_634)
);

OR2x2_ASAP7_75t_SL g635 ( 
.A(n_493),
.B(n_238),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_553),
.B(n_238),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_508),
.Y(n_637)
);

O2A1O1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_521),
.A2(n_550),
.B(n_555),
.C(n_579),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_L g639 ( 
.A(n_547),
.B(n_285),
.C(n_290),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_510),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_549),
.A2(n_285),
.B(n_290),
.C(n_360),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_526),
.B(n_28),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_510),
.B(n_29),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_542),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_535),
.B(n_30),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_534),
.B(n_30),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_531),
.B(n_32),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_556),
.A2(n_290),
.B1(n_380),
.B2(n_379),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_533),
.A2(n_360),
.B1(n_380),
.B2(n_379),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_546),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_560),
.B(n_32),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_552),
.A2(n_557),
.B(n_554),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_509),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

AO21x1_ASAP7_75t_L g655 ( 
.A1(n_505),
.A2(n_393),
.B(n_396),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_565),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_561),
.B(n_34),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_567),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_539),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_537),
.A2(n_379),
.B1(n_380),
.B2(n_393),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_511),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_499),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_538),
.A2(n_392),
.B(n_396),
.C(n_400),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_598),
.B(n_610),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_610),
.B(n_548),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_607),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_637),
.Y(n_668)
);

BUFx4f_ASAP7_75t_SL g669 ( 
.A(n_640),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_590),
.B(n_407),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_653),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_588),
.B(n_39),
.Y(n_672)
);

O2A1O1Ixp5_ASAP7_75t_L g673 ( 
.A1(n_655),
.A2(n_448),
.B(n_461),
.C(n_446),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_601),
.A2(n_411),
.B1(n_413),
.B2(n_415),
.Y(n_674)
);

INVx3_ASAP7_75t_SL g675 ( 
.A(n_590),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_601),
.Y(n_676)
);

AO21x2_ASAP7_75t_L g677 ( 
.A1(n_581),
.A2(n_448),
.B(n_461),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_584),
.B(n_582),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_605),
.B(n_42),
.Y(n_679)
);

AOI211xp5_ASAP7_75t_L g680 ( 
.A1(n_643),
.A2(n_415),
.B(n_423),
.C(n_425),
.Y(n_680)
);

AO21x1_ASAP7_75t_L g681 ( 
.A1(n_626),
.A2(n_423),
.B(n_425),
.Y(n_681)
);

OAI21x1_ASAP7_75t_SL g682 ( 
.A1(n_652),
.A2(n_44),
.B(n_45),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_585),
.B(n_654),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_583),
.B(n_48),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_633),
.B(n_50),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_625),
.Y(n_686)
);

AO31x2_ASAP7_75t_L g687 ( 
.A1(n_627),
.A2(n_454),
.A3(n_452),
.B(n_458),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_612),
.B(n_53),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_592),
.A2(n_429),
.B1(n_459),
.B2(n_442),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_603),
.Y(n_690)
);

OAI21x1_ASAP7_75t_SL g691 ( 
.A1(n_652),
.A2(n_55),
.B(n_56),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_602),
.A2(n_57),
.B(n_58),
.Y(n_692)
);

NAND2x1p5_ASAP7_75t_L g693 ( 
.A(n_620),
.B(n_467),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_585),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_590),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_650),
.B(n_59),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_587),
.A2(n_459),
.B1(n_442),
.B2(n_467),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_631),
.B(n_60),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_604),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_591),
.A2(n_61),
.B(n_62),
.Y(n_700)
);

NOR2x1_ASAP7_75t_L g701 ( 
.A(n_620),
.B(n_442),
.Y(n_701)
);

AOI21xp33_ASAP7_75t_L g702 ( 
.A1(n_586),
.A2(n_65),
.B(n_67),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_594),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_659),
.B(n_183),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_656),
.B(n_73),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_662),
.Y(n_706)
);

OAI21xp5_ASAP7_75t_L g707 ( 
.A1(n_634),
.A2(n_74),
.B(n_75),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_616),
.A2(n_91),
.B(n_92),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_645),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

BUFx12f_ASAP7_75t_L g711 ( 
.A(n_635),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_658),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_624),
.A2(n_103),
.B1(n_106),
.B2(n_116),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_657),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_714)
);

NOR2x1_ASAP7_75t_L g715 ( 
.A(n_630),
.B(n_120),
.Y(n_715)
);

AOI21xp33_ASAP7_75t_L g716 ( 
.A1(n_618),
.A2(n_595),
.B(n_619),
.Y(n_716)
);

AOI221x1_ASAP7_75t_L g717 ( 
.A1(n_639),
.A2(n_641),
.B1(n_647),
.B2(n_642),
.C(n_651),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_632),
.A2(n_122),
.B(n_124),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_SL g719 ( 
.A1(n_636),
.A2(n_130),
.B(n_131),
.C(n_134),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_660),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_609),
.A2(n_148),
.B(n_149),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_593),
.B(n_151),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_597),
.B(n_156),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_611),
.A2(n_160),
.B(n_162),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_600),
.B(n_164),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_606),
.B(n_614),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_596),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_617),
.B(n_654),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_623),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_621),
.B(n_646),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_622),
.A2(n_628),
.B(n_664),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_663),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_663),
.B(n_629),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_644),
.B(n_613),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_648),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_661),
.B(n_649),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_615),
.A2(n_562),
.B(n_580),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_638),
.A2(n_631),
.B(n_634),
.C(n_608),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_625),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_638),
.A2(n_631),
.B(n_634),
.C(n_608),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_588),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_588),
.B(n_578),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_610),
.B(n_588),
.Y(n_743)
);

BUFx4f_ASAP7_75t_L g744 ( 
.A(n_590),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_615),
.A2(n_562),
.B(n_580),
.Y(n_745)
);

AND3x4_ASAP7_75t_L g746 ( 
.A(n_635),
.B(n_571),
.C(n_530),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_638),
.A2(n_631),
.B(n_634),
.C(n_608),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_580),
.A2(n_608),
.B(n_551),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_588),
.B(n_578),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_588),
.B(n_578),
.Y(n_750)
);

OAI21x1_ASAP7_75t_SL g751 ( 
.A1(n_652),
.A2(n_610),
.B(n_638),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_580),
.A2(n_608),
.B(n_551),
.Y(n_752)
);

AOI221xp5_ASAP7_75t_SL g753 ( 
.A1(n_631),
.A2(n_395),
.B1(n_634),
.B2(n_586),
.C(n_589),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_601),
.Y(n_754)
);

CKINVDCx6p67_ASAP7_75t_R g755 ( 
.A(n_590),
.Y(n_755)
);

OA21x2_ASAP7_75t_L g756 ( 
.A1(n_599),
.A2(n_581),
.B(n_602),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_588),
.B(n_578),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_741),
.A2(n_711),
.B1(n_744),
.B2(n_742),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_749),
.B(n_750),
.Y(n_759)
);

AOI21xp33_ASAP7_75t_L g760 ( 
.A1(n_753),
.A2(n_678),
.B(n_726),
.Y(n_760)
);

INVx6_ASAP7_75t_SL g761 ( 
.A(n_670),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_670),
.B(n_686),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_738),
.B(n_747),
.C(n_740),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_667),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_667),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_712),
.Y(n_766)
);

INVx3_ASAP7_75t_SL g767 ( 
.A(n_755),
.Y(n_767)
);

OA21x2_ASAP7_75t_L g768 ( 
.A1(n_673),
.A2(n_717),
.B(n_692),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_757),
.B(n_743),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_720),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_699),
.B(n_743),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_668),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_671),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_703),
.B(n_690),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_730),
.B(n_676),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_744),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_706),
.Y(n_777)
);

NAND2x1_ASAP7_75t_L g778 ( 
.A(n_694),
.B(n_672),
.Y(n_778)
);

CKINVDCx6p67_ASAP7_75t_R g779 ( 
.A(n_675),
.Y(n_779)
);

OA21x2_ASAP7_75t_L g780 ( 
.A1(n_707),
.A2(n_708),
.B(n_681),
.Y(n_780)
);

BUFx12f_ASAP7_75t_L g781 ( 
.A(n_739),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_672),
.B(n_665),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_716),
.B(n_688),
.Y(n_783)
);

AO21x1_ASAP7_75t_L g784 ( 
.A1(n_702),
.A2(n_698),
.B(n_697),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_695),
.B(n_666),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_727),
.B(n_704),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_746),
.A2(n_704),
.B1(n_679),
.B2(n_723),
.Y(n_787)
);

OAI21x1_ASAP7_75t_SL g788 ( 
.A1(n_682),
.A2(n_691),
.B(n_731),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_669),
.B(n_734),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_694),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_732),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_732),
.B(n_723),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_710),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_728),
.B(n_733),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_693),
.B(n_710),
.Y(n_795)
);

AO21x2_ASAP7_75t_L g796 ( 
.A1(n_677),
.A2(n_697),
.B(n_735),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_685),
.A2(n_735),
.B(n_684),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_722),
.A2(n_756),
.B(n_736),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_705),
.Y(n_799)
);

OAI221xp5_ASAP7_75t_L g800 ( 
.A1(n_680),
.A2(n_713),
.B1(n_709),
.B2(n_714),
.C(n_715),
.Y(n_800)
);

INVx3_ASAP7_75t_SL g801 ( 
.A(n_729),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_696),
.B(n_725),
.Y(n_802)
);

AO31x2_ASAP7_75t_L g803 ( 
.A1(n_674),
.A2(n_718),
.A3(n_689),
.B(n_721),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_729),
.B(n_687),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_701),
.Y(n_805)
);

OA21x2_ASAP7_75t_L g806 ( 
.A1(n_724),
.A2(n_687),
.B(n_719),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_701),
.A2(n_683),
.B(n_687),
.Y(n_807)
);

BUFx6f_ASAP7_75t_SL g808 ( 
.A(n_686),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_741),
.A2(n_598),
.B1(n_754),
.B2(n_601),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_737),
.A2(n_580),
.B(n_745),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_667),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_743),
.Y(n_812)
);

BUFx8_ASAP7_75t_L g813 ( 
.A(n_711),
.Y(n_813)
);

NAND2x1p5_ASAP7_75t_L g814 ( 
.A(n_744),
.B(n_610),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_741),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_755),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_667),
.Y(n_817)
);

OAI21x1_ASAP7_75t_SL g818 ( 
.A1(n_751),
.A2(n_700),
.B(n_691),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_743),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_741),
.B(n_515),
.Y(n_820)
);

OAI21x1_ASAP7_75t_SL g821 ( 
.A1(n_751),
.A2(n_700),
.B(n_691),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_667),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_755),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_741),
.A2(n_598),
.B1(n_754),
.B2(n_601),
.Y(n_824)
);

BUFx2_ASAP7_75t_R g825 ( 
.A(n_675),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_743),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_667),
.Y(n_827)
);

AO21x2_ASAP7_75t_L g828 ( 
.A1(n_748),
.A2(n_752),
.B(n_745),
.Y(n_828)
);

BUFx12f_ASAP7_75t_L g829 ( 
.A(n_711),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_667),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_742),
.Y(n_831)
);

INVx2_ASAP7_75t_R g832 ( 
.A(n_667),
.Y(n_832)
);

AO21x2_ASAP7_75t_L g833 ( 
.A1(n_748),
.A2(n_752),
.B(n_745),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_764),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_765),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_819),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_820),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_804),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_809),
.A2(n_824),
.B1(n_786),
.B2(n_782),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_814),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_831),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_811),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_766),
.B(n_773),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_817),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_817),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_826),
.Y(n_846)
);

AO21x1_ASAP7_75t_SL g847 ( 
.A1(n_807),
.A2(n_787),
.B(n_827),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_822),
.Y(n_848)
);

AOI21xp33_ASAP7_75t_L g849 ( 
.A1(n_783),
.A2(n_760),
.B(n_800),
.Y(n_849)
);

AO21x1_ASAP7_75t_SL g850 ( 
.A1(n_807),
.A2(n_830),
.B(n_827),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_784),
.A2(n_763),
.B(n_818),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_830),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_816),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_774),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_812),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_828),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_778),
.B(n_792),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_769),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_759),
.A2(n_782),
.B1(n_794),
.B2(n_775),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_791),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_770),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_815),
.B(n_771),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_767),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_785),
.B(n_758),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_833),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_832),
.Y(n_866)
);

INVx8_ASAP7_75t_L g867 ( 
.A(n_812),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_772),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_777),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_785),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_801),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_776),
.A2(n_762),
.B1(n_761),
.B2(n_779),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_794),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_776),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_761),
.A2(n_792),
.B1(n_762),
.B2(n_802),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_805),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_790),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_793),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_763),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_789),
.B(n_781),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_796),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_790),
.B(n_799),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_821),
.B(n_788),
.Y(n_883)
);

AOI211xp5_ASAP7_75t_L g884 ( 
.A1(n_799),
.A2(n_798),
.B(n_797),
.C(n_810),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_834),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_841),
.B(n_795),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_858),
.B(n_823),
.Y(n_887)
);

INVx11_ASAP7_75t_L g888 ( 
.A(n_853),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_854),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_838),
.B(n_798),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_834),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_838),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_839),
.A2(n_829),
.B1(n_813),
.B2(n_797),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_843),
.B(n_813),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_879),
.B(n_768),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_879),
.B(n_780),
.Y(n_896)
);

NOR2x1_ASAP7_75t_L g897 ( 
.A(n_872),
.B(n_806),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_849),
.A2(n_847),
.B1(n_859),
.B2(n_864),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_856),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_883),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_842),
.B(n_845),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_878),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_835),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_853),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_844),
.B(n_806),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_844),
.B(n_803),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_837),
.B(n_825),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_848),
.B(n_852),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_852),
.B(n_808),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_866),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_857),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_900),
.B(n_883),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_906),
.B(n_850),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_893),
.A2(n_847),
.B1(n_873),
.B2(n_875),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_892),
.B(n_865),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_906),
.B(n_850),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_892),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_885),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_902),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_889),
.B(n_860),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_891),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_901),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_899),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_909),
.Y(n_924)
);

AND2x4_ASAP7_75t_SL g925 ( 
.A(n_911),
.B(n_857),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_898),
.A2(n_870),
.B1(n_876),
.B2(n_862),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_905),
.B(n_881),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_905),
.B(n_910),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_909),
.A2(n_840),
.B1(n_882),
.B2(n_884),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_908),
.B(n_851),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_920),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_930),
.B(n_895),
.Y(n_932)
);

INVx5_ASAP7_75t_L g933 ( 
.A(n_912),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_930),
.B(n_895),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_928),
.B(n_896),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_922),
.B(n_928),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_913),
.B(n_896),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_918),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_923),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_922),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_917),
.B(n_871),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_919),
.B(n_890),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_916),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_924),
.B(n_903),
.Y(n_944)
);

NAND2x1p5_ASAP7_75t_L g945 ( 
.A(n_912),
.B(n_911),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_912),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_931),
.B(n_921),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_936),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_938),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_939),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_935),
.B(n_921),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_932),
.B(n_934),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_943),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_943),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_940),
.B(n_915),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_944),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_942),
.B(n_927),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_956),
.B(n_935),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_957),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_957),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_947),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_949),
.Y(n_962)
);

AOI32xp33_ASAP7_75t_L g963 ( 
.A1(n_953),
.A2(n_937),
.A3(n_925),
.B1(n_946),
.B2(n_934),
.Y(n_963)
);

XNOR2xp5_ASAP7_75t_L g964 ( 
.A(n_954),
.B(n_904),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_952),
.A2(n_933),
.B1(n_945),
.B2(n_929),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_950),
.A2(n_941),
.B(n_897),
.Y(n_966)
);

INVxp33_ASAP7_75t_L g967 ( 
.A(n_955),
.Y(n_967)
);

OAI31xp33_ASAP7_75t_L g968 ( 
.A1(n_952),
.A2(n_907),
.A3(n_945),
.B(n_914),
.Y(n_968)
);

XNOR2x1_ASAP7_75t_L g969 ( 
.A(n_964),
.B(n_863),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_966),
.A2(n_897),
.B(n_894),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_968),
.A2(n_946),
.B1(n_912),
.B2(n_948),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_962),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_959),
.Y(n_973)
);

AOI211xp5_ASAP7_75t_L g974 ( 
.A1(n_970),
.A2(n_965),
.B(n_966),
.C(n_967),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_969),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_973),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_975),
.A2(n_971),
.B1(n_970),
.B2(n_961),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_976),
.B(n_972),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_978),
.Y(n_979)
);

AO22x2_ASAP7_75t_L g980 ( 
.A1(n_977),
.A2(n_887),
.B1(n_974),
.B2(n_960),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_979),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_980),
.B(n_888),
.Y(n_982)
);

XNOR2xp5_ASAP7_75t_L g983 ( 
.A(n_981),
.B(n_980),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_982),
.Y(n_984)
);

AND3x1_ASAP7_75t_L g985 ( 
.A(n_984),
.B(n_880),
.C(n_888),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_984),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_983),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_L g988 ( 
.A1(n_986),
.A2(n_874),
.B1(n_963),
.B2(n_926),
.C(n_840),
.Y(n_988)
);

OAI22x1_ASAP7_75t_SL g989 ( 
.A1(n_987),
.A2(n_840),
.B1(n_933),
.B2(n_911),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_985),
.A2(n_958),
.B1(n_871),
.B2(n_929),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_987),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_985),
.A2(n_945),
.B1(n_933),
.B2(n_911),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_991),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_989),
.Y(n_994)
);

OAI331xp33_ASAP7_75t_L g995 ( 
.A1(n_988),
.A2(n_886),
.A3(n_861),
.B1(n_877),
.B2(n_868),
.B3(n_869),
.C1(n_951),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_990),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_992),
.A2(n_933),
.B1(n_942),
.B2(n_871),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_991),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_991),
.A2(n_871),
.B(n_846),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_993),
.A2(n_871),
.B(n_836),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_998),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_SL g1002 ( 
.A1(n_994),
.A2(n_925),
.B(n_946),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_SL g1003 ( 
.A1(n_1001),
.A2(n_999),
.B(n_996),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_1003),
.A2(n_1000),
.B(n_1002),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_1004),
.B(n_997),
.Y(n_1005)
);

AOI221xp5_ASAP7_75t_L g1006 ( 
.A1(n_1005),
.A2(n_995),
.B1(n_836),
.B2(n_846),
.C(n_867),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_1006),
.A2(n_933),
.B1(n_867),
.B2(n_855),
.Y(n_1007)
);


endmodule