module fake_netlist_5_1376_n_1213 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1213);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1213;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_1194;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_1166;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_1141;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_1178;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_1161;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_1150;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_1139;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_1055;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_547;
wire n_1191;
wire n_1198;
wire n_721;
wire n_998;
wire n_1157;
wire n_1099;
wire n_841;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_983;
wire n_725;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_1203;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_1179;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_212;
wire n_933;
wire n_788;
wire n_507;
wire n_1152;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_1195;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_936;
wire n_947;
wire n_373;
wire n_820;
wire n_1090;
wire n_757;
wire n_1200;
wire n_307;
wire n_633;
wire n_1192;
wire n_439;
wire n_530;
wire n_1024;
wire n_1107;
wire n_1063;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1185;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1143;
wire n_513;
wire n_804;
wire n_867;
wire n_186;
wire n_1124;
wire n_537;
wire n_1158;
wire n_902;
wire n_191;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_1104;
wire n_792;
wire n_563;
wire n_171;
wire n_1182;
wire n_756;
wire n_1145;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_992;
wire n_1049;
wire n_1153;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_1068;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_1154;
wire n_286;
wire n_883;
wire n_1135;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_1163;
wire n_406;
wire n_1108;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_519;
wire n_325;
wire n_449;
wire n_1100;
wire n_1207;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_1147;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_940;
wire n_618;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_1169;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1172;
wire n_167;
wire n_976;
wire n_1096;
wire n_1095;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_1208;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_1168;
wire n_192;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_1142;
wire n_660;
wire n_223;
wire n_1201;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_1148;
wire n_264;
wire n_750;
wire n_472;
wire n_742;
wire n_669;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_1176;
wire n_374;
wire n_276;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_1149;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1073;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_181;
wire n_962;
wire n_436;
wire n_1204;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_1171;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1188;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1071;
wire n_1043;
wire n_496;
wire n_1165;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_1177;
wire n_680;
wire n_168;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_1159;
wire n_1210;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_328;
wire n_214;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_1167;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_829;
wire n_928;
wire n_749;
wire n_1064;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_1151;
wire n_1134;
wire n_881;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_1173;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_236;
wire n_1075;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_1193;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_1197;
wire n_1211;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1187;
wire n_1015;
wire n_1000;
wire n_891;
wire n_1140;
wire n_239;
wire n_466;
wire n_1164;
wire n_420;
wire n_630;
wire n_1202;
wire n_632;
wire n_699;
wire n_489;
wire n_1174;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_846;
wire n_586;
wire n_1058;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_170;
wire n_1101;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_1190;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_1212;
wire n_767;
wire n_206;
wire n_172;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_1175;
wire n_861;
wire n_534;
wire n_948;
wire n_1183;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_1131;
wire n_176;
wire n_1133;
wire n_970;
wire n_911;
wire n_557;
wire n_182;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_679;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_857;
wire n_795;
wire n_695;
wire n_832;
wire n_180;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_207;
wire n_561;
wire n_1044;
wire n_1205;
wire n_346;
wire n_937;
wire n_1209;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_1130;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_1156;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_1136;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_1037;
wire n_1160;
wire n_202;
wire n_1080;
wire n_266;
wire n_1162;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_1199;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_808;
wire n_1038;
wire n_520;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_1181;
wire n_1196;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_1138;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_1186;
wire n_242;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_222;
wire n_1155;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_1184;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_1189;
wire n_348;
wire n_1029;
wire n_166;
wire n_626;
wire n_925;
wire n_1180;
wire n_1206;
wire n_424;
wire n_1003;
wire n_1144;
wire n_1137;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_1170;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_9),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_75),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_83),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_122),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_34),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_95),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_49),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_33),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_48),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_82),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_39),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_45),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_68),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_110),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_38),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_89),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_33),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_18),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_88),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_43),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_3),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_137),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_134),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_36),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_61),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_30),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_47),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_91),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_144),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_56),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_162),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_90),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_142),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_30),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_15),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_151),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_25),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_19),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_174),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_176),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_178),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_179),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_180),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_181),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_182),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_183),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_188),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_196),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_175),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_191),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_199),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_165),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_200),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_201),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_203),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_204),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_239),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_227),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_233),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_235),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_244),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_245),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_249),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_250),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_252),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_240),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_228),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_224),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_243),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_224),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_256),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_262),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_262),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_266),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_266),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_273),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_273),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_253),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_261),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_277),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_277),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_271),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_278),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_278),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_299),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_268),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_271),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_303),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_280),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_254),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_258),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_281),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_211),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_294),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_287),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_287),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_296),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_290),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_298),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_327),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_307),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_327),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_332),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_341),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_326),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_332),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_354),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_319),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_326),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_305),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_269),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_306),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_308),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_323),
.B(n_301),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_318),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_317),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_345),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_320),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_321),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_345),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_322),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_331),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_324),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_325),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_315),
.B(n_301),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_329),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_276),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_354),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_347),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_350),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_352),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_336),
.B(n_334),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_363),
.A2(n_295),
.B1(n_297),
.B2(n_304),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_346),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_393),
.A2(n_304),
.B1(n_351),
.B2(n_348),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_316),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_380),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_380),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g411 ( 
.A1(n_369),
.A2(n_388),
.B(n_385),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_349),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_350),
.Y(n_414)
);

NOR2x1_ASAP7_75t_L g415 ( 
.A(n_357),
.B(n_215),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_397),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_395),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_396),
.B(n_284),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_365),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_372),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_366),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_378),
.B(n_311),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_221),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_394),
.A2(n_335),
.B1(n_313),
.B2(n_311),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_359),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_376),
.B(n_313),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

INVx6_ASAP7_75t_L g435 ( 
.A(n_400),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_284),
.Y(n_436)
);

BUFx12f_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_377),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_381),
.B(n_354),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_L g443 ( 
.A(n_384),
.B(n_387),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_390),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_390),
.B(n_255),
.Y(n_446)
);

CKINVDCx6p67_ASAP7_75t_R g447 ( 
.A(n_383),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_391),
.B(n_302),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_370),
.B(n_270),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_391),
.B(n_302),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_399),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_361),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_399),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

CKINVDCx6p67_ASAP7_75t_R g456 ( 
.A(n_386),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_361),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_367),
.Y(n_459)
);

CKINVDCx8_ASAP7_75t_R g460 ( 
.A(n_371),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_396),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_369),
.A2(n_279),
.B(n_274),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_363),
.A2(n_335),
.B1(n_220),
.B2(n_222),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_364),
.B(n_260),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_363),
.A2(n_166),
.B1(n_218),
.B2(n_217),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_363),
.B(n_309),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_363),
.B(n_309),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_363),
.A2(n_186),
.B1(n_197),
.B2(n_205),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_364),
.B(n_260),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_395),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

INVx6_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_392),
.B(n_221),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_362),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_379),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_364),
.B(n_259),
.Y(n_484)
);

AND2x2_ASAP7_75t_SL g485 ( 
.A(n_400),
.B(n_173),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_363),
.B(n_192),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_363),
.B(n_202),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_392),
.B(n_272),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_362),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_379),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_363),
.B(n_166),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_363),
.B(n_196),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_364),
.B(n_275),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_432),
.B(n_184),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_418),
.B(n_283),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_416),
.B(n_207),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_464),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_477),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_425),
.B(n_279),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_480),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_490),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_411),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_408),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_407),
.A2(n_209),
.B1(n_210),
.B2(n_213),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_425),
.B(n_264),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_463),
.B(n_265),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_421),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_408),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_416),
.B(n_214),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_419),
.B(n_264),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_419),
.B(n_267),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_413),
.B(n_267),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_406),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_468),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_463),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_432),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_412),
.A2(n_189),
.B(n_185),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_407),
.B(n_265),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_410),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_483),
.B(n_190),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_467),
.B(n_169),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_467),
.Y(n_534)
);

INVx6_ASAP7_75t_L g535 ( 
.A(n_410),
.Y(n_535)
);

INVxp33_ASAP7_75t_SL g536 ( 
.A(n_423),
.Y(n_536)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_491),
.B(n_472),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_461),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_475),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_461),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_475),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_414),
.B(n_194),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_470),
.B(n_198),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_474),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_488),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_458),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_488),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_462),
.B(n_35),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_484),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_484),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_492),
.B(n_169),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_427),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_412),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_536),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_526),
.Y(n_558)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_555),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_555),
.B(n_453),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_505),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_549),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g563 ( 
.A(n_538),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_535),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_536),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_549),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_505),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_524),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_506),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_552),
.B(n_494),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_538),
.B(n_491),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_500),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_542),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_501),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_506),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_556),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_506),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_496),
.B(n_427),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_551),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_506),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_512),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_512),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_512),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_512),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_515),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_R g587 ( 
.A(n_551),
.B(n_457),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_526),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_515),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_535),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_504),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_515),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_535),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_507),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_502),
.B(n_433),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_571),
.B(n_534),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_572),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_558),
.Y(n_598)
);

AO21x2_ASAP7_75t_L g599 ( 
.A1(n_561),
.A2(n_499),
.B(n_495),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_558),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_561),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_563),
.B(n_459),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g603 ( 
.A(n_595),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_567),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_558),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_576),
.B(n_496),
.Y(n_606)
);

INVxp33_ASAP7_75t_SL g607 ( 
.A(n_560),
.Y(n_607)
);

CKINVDCx6p67_ASAP7_75t_R g608 ( 
.A(n_559),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_588),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_567),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_557),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_594),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_570),
.B(n_540),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_568),
.B(n_544),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_574),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_594),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_588),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_588),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_566),
.A2(n_429),
.B1(n_433),
.B2(n_441),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_579),
.B(n_510),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_579),
.B(n_528),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_579),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_573),
.B(n_472),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_580),
.B(n_440),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_591),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_592),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_592),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_592),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_592),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_562),
.B(n_486),
.Y(n_630)
);

AOI21x1_ASAP7_75t_L g631 ( 
.A1(n_578),
.A2(n_527),
.B(n_499),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_569),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_569),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_569),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_564),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_584),
.B(n_440),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_584),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_564),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_587),
.A2(n_471),
.B1(n_485),
.B2(n_443),
.Y(n_639)
);

NOR2x1p5_ASAP7_75t_L g640 ( 
.A(n_565),
.B(n_447),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_575),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_577),
.B(n_526),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_581),
.Y(n_643)
);

CKINVDCx16_ASAP7_75t_R g644 ( 
.A(n_590),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_582),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_583),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_590),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_585),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_586),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_589),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_578),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_593),
.A2(n_487),
.B1(n_486),
.B2(n_452),
.Y(n_652)
);

CKINVDCx6p67_ASAP7_75t_R g653 ( 
.A(n_593),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_566),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_563),
.A2(n_403),
.B1(n_452),
.B2(n_428),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_595),
.B(n_487),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_564),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_561),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_571),
.B(n_545),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_595),
.B(n_497),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_561),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_572),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_571),
.B(n_511),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_595),
.B(n_554),
.Y(n_664)
);

INVx6_ASAP7_75t_L g665 ( 
.A(n_559),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_558),
.B(n_495),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_595),
.A2(n_545),
.B1(n_466),
.B2(n_415),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_595),
.B(n_554),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_564),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_558),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_561),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_595),
.B(n_508),
.C(n_466),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_561),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_595),
.B(n_439),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_561),
.Y(n_675)
);

AND3x2_ASAP7_75t_L g676 ( 
.A(n_595),
.B(n_444),
.C(n_442),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_656),
.B(n_533),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_611),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_607),
.B(n_427),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_625),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_599),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_672),
.B(n_469),
.C(n_455),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_599),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_597),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_663),
.B(n_530),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_660),
.B(n_523),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_611),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_615),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_628),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_628),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_617),
.B(n_523),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_603),
.B(n_430),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_599),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_622),
.B(n_514),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_662),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_601),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_663),
.B(n_530),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_601),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_665),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_604),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_604),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_603),
.B(n_430),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_610),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_659),
.B(n_498),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_665),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_610),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_612),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_639),
.A2(n_445),
.B1(n_438),
.B2(n_430),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_655),
.B(n_438),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_628),
.Y(n_710)
);

INVx4_ASAP7_75t_SL g711 ( 
.A(n_666),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_616),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_616),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_658),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_665),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_667),
.A2(n_530),
.B1(n_217),
.B2(n_218),
.Y(n_716)
);

BUFx8_ASAP7_75t_SL g717 ( 
.A(n_647),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_596),
.B(n_511),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_596),
.B(n_525),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_661),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_628),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_671),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_673),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_617),
.B(n_525),
.Y(n_725)
);

INVx4_ASAP7_75t_SL g726 ( 
.A(n_666),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_646),
.B(n_515),
.Y(n_727)
);

NAND3x1_ASAP7_75t_L g728 ( 
.A(n_674),
.B(n_473),
.C(n_448),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_598),
.B(n_518),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_R g730 ( 
.A(n_644),
.B(n_438),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_664),
.B(n_446),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_668),
.B(n_451),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_673),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_675),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_675),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_624),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_641),
.B(n_446),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_652),
.B(n_451),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_624),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_613),
.B(n_522),
.Y(n_740)
);

BUFx4f_ASAP7_75t_L g741 ( 
.A(n_608),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_646),
.Y(n_742)
);

OR2x2_ASAP7_75t_SL g743 ( 
.A(n_602),
.B(n_435),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_641),
.B(n_448),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_659),
.B(n_498),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_598),
.B(n_518),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_646),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_630),
.A2(n_216),
.B1(n_532),
.B2(n_531),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_666),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_648),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_614),
.B(n_509),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_607),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_628),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_666),
.Y(n_754)
);

AO22x2_ASAP7_75t_L g755 ( 
.A1(n_709),
.A2(n_636),
.B1(n_619),
.B2(n_621),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_699),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_678),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_741),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_684),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_716),
.A2(n_623),
.B1(n_653),
.B2(n_645),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_699),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_688),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_695),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_SL g764 ( 
.A1(n_715),
.A2(n_637),
.B1(n_650),
.B2(n_643),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_754),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_731),
.B(n_636),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_750),
.B(n_653),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_682),
.A2(n_608),
.B1(n_606),
.B2(n_620),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_741),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_728),
.A2(n_606),
.B1(n_676),
.B2(n_654),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_737),
.B(n_648),
.Y(n_771)
);

NAND2x1p5_ASAP7_75t_L g772 ( 
.A(n_715),
.B(n_622),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_680),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_751),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_738),
.A2(n_620),
.B1(n_621),
.B2(n_426),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_742),
.Y(n_776)
);

NAND3x1_ASAP7_75t_L g777 ( 
.A(n_744),
.B(n_638),
.C(n_651),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_742),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_747),
.B(n_649),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_736),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_739),
.Y(n_781)
);

AND2x6_ASAP7_75t_L g782 ( 
.A(n_689),
.B(n_649),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_747),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_700),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_704),
.B(n_642),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_730),
.Y(n_786)
);

AO22x2_ASAP7_75t_L g787 ( 
.A1(n_709),
.A2(n_642),
.B1(n_633),
.B2(n_634),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_692),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_749),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_711),
.B(n_635),
.Y(n_790)
);

BUFx4_ASAP7_75t_L g791 ( 
.A(n_730),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_685),
.B(n_626),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_717),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_SL g794 ( 
.A(n_687),
.B(n_460),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_711),
.B(n_635),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_SL g796 ( 
.A1(n_743),
.A2(n_454),
.B1(n_451),
.B2(n_437),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_703),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_727),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_706),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_711),
.B(n_657),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_692),
.Y(n_801)
);

NAND2x1p5_ASAP7_75t_L g802 ( 
.A(n_702),
.B(n_622),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_696),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_752),
.B(n_409),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_697),
.B(n_626),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_713),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_704),
.B(n_598),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_696),
.Y(n_808)
);

CKINVDCx16_ASAP7_75t_R g809 ( 
.A(n_679),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_708),
.B(n_454),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_689),
.B(n_632),
.Y(n_811)
);

INVx8_ASAP7_75t_L g812 ( 
.A(n_717),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_714),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_698),
.Y(n_814)
);

NAND2x1p5_ASAP7_75t_L g815 ( 
.A(n_702),
.B(n_622),
.Y(n_815)
);

NOR2x1p5_ASAP7_75t_L g816 ( 
.A(n_677),
.B(n_456),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_719),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_738),
.A2(n_478),
.B1(n_435),
.B2(n_449),
.Y(n_818)
);

AO22x2_ASAP7_75t_L g819 ( 
.A1(n_732),
.A2(n_629),
.B1(n_669),
.B2(n_657),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_705),
.Y(n_820)
);

AO22x2_ASAP7_75t_L g821 ( 
.A1(n_732),
.A2(n_669),
.B1(n_627),
.B2(n_605),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_718),
.B(n_627),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_727),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_812),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_759),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_774),
.B(n_745),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_807),
.B(n_745),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_770),
.B(n_454),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_785),
.B(n_723),
.Y(n_829)
);

CKINVDCx11_ASAP7_75t_R g830 ( 
.A(n_812),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_788),
.B(n_720),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_766),
.B(n_734),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_762),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_771),
.B(n_749),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_763),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_809),
.A2(n_716),
.B1(n_748),
.B2(n_740),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_780),
.B(n_686),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_781),
.B(n_698),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_801),
.B(n_701),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_773),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_764),
.B(n_729),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_784),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_797),
.B(n_701),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_768),
.B(n_748),
.C(n_516),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_767),
.B(n_707),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_779),
.B(n_729),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_803),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_779),
.B(n_622),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_799),
.B(n_707),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_756),
.B(n_729),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_808),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_806),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_765),
.B(n_681),
.Y(n_853)
);

O2A1O1Ixp5_ASAP7_75t_L g854 ( 
.A1(n_810),
.A2(n_631),
.B(n_753),
.C(n_710),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_813),
.B(n_712),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_814),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_761),
.B(n_712),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_760),
.B(n_746),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_796),
.B(n_726),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_817),
.B(n_721),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_L g861 ( 
.A(n_775),
.B(n_516),
.C(n_450),
.Y(n_861)
);

OAI22xp33_ASAP7_75t_L g862 ( 
.A1(n_818),
.A2(n_689),
.B1(n_722),
.B2(n_690),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_822),
.B(n_724),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_821),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_755),
.B(n_733),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_821),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_804),
.B(n_431),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_755),
.B(n_733),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_792),
.B(n_735),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_805),
.B(n_783),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_787),
.B(n_735),
.Y(n_871)
);

CKINVDCx11_ASAP7_75t_R g872 ( 
.A(n_793),
.Y(n_872)
);

NAND2xp33_ASAP7_75t_SL g873 ( 
.A(n_758),
.B(n_640),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_819),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_787),
.B(n_691),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_776),
.B(n_691),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_776),
.B(n_691),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_776),
.B(n_726),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_778),
.B(n_725),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_778),
.B(n_725),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_758),
.B(n_469),
.C(n_450),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_816),
.A2(n_216),
.B1(n_212),
.B2(n_172),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_802),
.B(n_746),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_778),
.B(n_726),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_819),
.B(n_725),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_786),
.A2(n_527),
.B1(n_690),
.B2(n_689),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_769),
.A2(n_690),
.B1(n_722),
.B2(n_694),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_789),
.B(n_683),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_791),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_823),
.B(n_693),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_777),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_757),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_820),
.Y(n_893)
);

BUFx12f_ASAP7_75t_L g894 ( 
.A(n_769),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_815),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_866),
.B(n_693),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_830),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_871),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_827),
.B(n_782),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_864),
.B(n_798),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_825),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_894),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_891),
.B(n_826),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_864),
.B(n_798),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_889),
.B(n_798),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_833),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_893),
.B(n_794),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_874),
.B(n_782),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_842),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_835),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_852),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_870),
.B(n_790),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_865),
.B(n_782),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_853),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_868),
.B(n_840),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_824),
.B(n_417),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_847),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_851),
.B(n_811),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_856),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_838),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_857),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_888),
.Y(n_922)
);

AND2x2_ASAP7_75t_SL g923 ( 
.A(n_841),
.B(n_795),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_831),
.B(n_795),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_844),
.A2(n_772),
.B(n_800),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_843),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_841),
.B(n_887),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_885),
.B(n_800),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_832),
.B(n_829),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_875),
.B(n_694),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_849),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_855),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_831),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_839),
.B(n_811),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_837),
.B(n_811),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_863),
.B(n_527),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_895),
.B(n_746),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_860),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_848),
.B(n_710),
.Y(n_939)
);

NAND2xp33_ASAP7_75t_SL g940 ( 
.A(n_859),
.B(n_791),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_890),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_845),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_869),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_834),
.B(n_753),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_897),
.B(n_887),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_933),
.B(n_846),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_929),
.B(n_846),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_897),
.B(n_862),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_927),
.A2(n_873),
.B(n_836),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_929),
.B(n_883),
.Y(n_950)
);

AOI21x1_ASAP7_75t_L g951 ( 
.A1(n_903),
.A2(n_904),
.B(n_900),
.Y(n_951)
);

BUFx4f_ASAP7_75t_L g952 ( 
.A(n_897),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_908),
.B(n_883),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_940),
.A2(n_828),
.B(n_862),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_923),
.B(n_850),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_897),
.B(n_892),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_900),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_925),
.A2(n_884),
.B(n_878),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_897),
.B(n_886),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_909),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_923),
.A2(n_886),
.B1(n_858),
.B2(n_882),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_925),
.A2(n_861),
.B(n_882),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_923),
.A2(n_881),
.B(n_854),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_897),
.B(n_858),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_898),
.A2(n_915),
.B(n_913),
.C(n_881),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_902),
.B(n_850),
.Y(n_966)
);

O2A1O1Ixp5_ASAP7_75t_L g967 ( 
.A1(n_913),
.A2(n_854),
.B(n_879),
.C(n_877),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_935),
.B(n_876),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_935),
.B(n_880),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_915),
.A2(n_902),
.B(n_899),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_908),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_904),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_920),
.B(n_867),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_902),
.B(n_690),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_L g975 ( 
.A(n_924),
.B(n_872),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_902),
.A2(n_722),
.B(n_449),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_920),
.B(n_600),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_930),
.A2(n_212),
.B(n_172),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_934),
.B(n_722),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_SL g980 ( 
.A(n_907),
.B(n_435),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_934),
.A2(n_489),
.B(n_481),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_918),
.A2(n_632),
.B(n_434),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_928),
.B(n_476),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_938),
.B(n_670),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_938),
.B(n_943),
.Y(n_985)
);

AOI22x1_ASAP7_75t_L g986 ( 
.A1(n_908),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_930),
.B(n_926),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_918),
.A2(n_632),
.B(n_605),
.Y(n_988)
);

INVxp67_ASAP7_75t_SL g989 ( 
.A(n_896),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_908),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_939),
.B(n_600),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_896),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_928),
.B(n_478),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_916),
.A2(n_167),
.B(n_168),
.C(n_170),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_905),
.A2(n_546),
.B(n_605),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_936),
.A2(n_618),
.B(n_609),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_936),
.A2(n_618),
.B(n_609),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_939),
.A2(n_546),
.B1(n_426),
.B2(n_478),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_901),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_950),
.B(n_922),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_956),
.B(n_912),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_963),
.A2(n_941),
.B(n_922),
.C(n_939),
.Y(n_1002)
);

NAND2x1p5_ASAP7_75t_L g1003 ( 
.A(n_945),
.B(n_914),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_952),
.B(n_975),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_948),
.A2(n_917),
.B(n_911),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_952),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_999),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_993),
.B(n_912),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_949),
.A2(n_941),
.B(n_922),
.C(n_921),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_962),
.A2(n_941),
.B(n_906),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_955),
.B(n_953),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_959),
.A2(n_906),
.B(n_901),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_999),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_954),
.B(n_944),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_961),
.A2(n_910),
.B(n_931),
.Y(n_1015)
);

OR2x2_ASAP7_75t_SL g1016 ( 
.A(n_973),
.B(n_942),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_965),
.B(n_932),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_981),
.B(n_921),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_953),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_967),
.A2(n_910),
.B(n_919),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1007),
.B(n_992),
.Y(n_1021)
);

NAND2x1p5_ASAP7_75t_L g1022 ( 
.A(n_1006),
.B(n_974),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_1004),
.B(n_983),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_1003),
.A2(n_964),
.B(n_978),
.C(n_967),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_1017),
.B(n_987),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_1003),
.B(n_970),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_1000),
.B(n_947),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1016),
.A2(n_958),
.B1(n_951),
.B2(n_957),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1011),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1019),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1006),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1008),
.B(n_971),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_1006),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_1012),
.A2(n_982),
.B(n_976),
.C(n_989),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1015),
.A2(n_966),
.B(n_979),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_1005),
.A2(n_990),
.B(n_971),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_1013),
.Y(n_1037)
);

INVxp67_ASAP7_75t_SL g1038 ( 
.A(n_1014),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_1002),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_1010),
.B(n_985),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_1018),
.A2(n_990),
.B1(n_986),
.B2(n_972),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1020),
.B(n_992),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1009),
.A2(n_946),
.B1(n_969),
.B2(n_968),
.Y(n_1043)
);

AO22x1_ASAP7_75t_L g1044 ( 
.A1(n_1001),
.A2(n_989),
.B1(n_995),
.B2(n_960),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_1006),
.B(n_988),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1031),
.B(n_991),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1037),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_1026),
.A2(n_998),
.B1(n_980),
.B2(n_937),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_1033),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1030),
.B(n_977),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1039),
.A2(n_996),
.B1(n_997),
.B2(n_984),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1038),
.B(n_932),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1049),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_1047),
.A2(n_1036),
.B(n_1028),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_1053),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_SL g1056 ( 
.A(n_1053),
.B(n_1039),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1054),
.B(n_1029),
.Y(n_1057)
);

AO21x2_ASAP7_75t_L g1058 ( 
.A1(n_1057),
.A2(n_1028),
.B(n_1042),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1056),
.B(n_1046),
.Y(n_1059)
);

AOI221xp5_ASAP7_75t_L g1060 ( 
.A1(n_1055),
.A2(n_1024),
.B1(n_1042),
.B2(n_1051),
.C(n_1044),
.Y(n_1060)
);

OA21x2_ASAP7_75t_L g1061 ( 
.A1(n_1060),
.A2(n_1051),
.B(n_1021),
.Y(n_1061)
);

CKINVDCx16_ASAP7_75t_R g1062 ( 
.A(n_1059),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1061),
.A2(n_1058),
.B(n_1034),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1062),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1064),
.Y(n_1065)
);

INVx3_ASAP7_75t_SL g1066 ( 
.A(n_1063),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1065),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1066),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1067),
.B(n_1061),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_1032),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_1070),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1069),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_1071),
.B(n_1052),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1072),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1071),
.B(n_1023),
.Y(n_1075)
);

INVxp33_ASAP7_75t_L g1076 ( 
.A(n_1075),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1074),
.B(n_1050),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1073),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_1078),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1077),
.A2(n_1045),
.B1(n_1021),
.B2(n_1041),
.Y(n_1080)
);

NAND2x1p5_ASAP7_75t_L g1081 ( 
.A(n_1079),
.B(n_1076),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1080),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1082),
.B(n_1045),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1083),
.B(n_1025),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1084),
.B(n_1040),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1086),
.B(n_1085),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1086),
.B(n_1048),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1087),
.B(n_1045),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1088),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1089),
.A2(n_1043),
.B1(n_1022),
.B2(n_1035),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1090),
.B(n_0),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_1089),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1093),
.A2(n_219),
.B(n_494),
.C(n_994),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1092),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1091),
.B(n_1022),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1096),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1095),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1098),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1097),
.A2(n_1094),
.B1(n_1043),
.B2(n_219),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1100),
.A2(n_1027),
.B1(n_551),
.B2(n_2),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1101),
.Y(n_1103)
);

AOI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_1102),
.A2(n_0),
.B(n_1),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1103),
.B(n_1),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1104),
.B(n_3),
.Y(n_1106)
);

AOI221xp5_ASAP7_75t_L g1107 ( 
.A1(n_1106),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_1105),
.B(n_4),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1108),
.B(n_5),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1107),
.B(n_6),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1108),
.B(n_7),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1109),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1110),
.A2(n_8),
.B(n_9),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_SL g1114 ( 
.A1(n_1111),
.A2(n_8),
.B(n_10),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1113),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1112),
.B(n_11),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1115),
.Y(n_1117)
);

NAND2x1_ASAP7_75t_L g1118 ( 
.A(n_1116),
.B(n_1114),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1117),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_1119)
);

AOI211xp5_ASAP7_75t_SL g1120 ( 
.A1(n_1118),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1120),
.B(n_16),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_16),
.C(n_17),
.Y(n_1122)
);

NAND4xp25_ASAP7_75t_SL g1123 ( 
.A(n_1121),
.B(n_17),
.C(n_18),
.D(n_19),
.Y(n_1123)
);

OAI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.C(n_23),
.Y(n_1124)
);

NAND3xp33_ASAP7_75t_SL g1125 ( 
.A(n_1124),
.B(n_20),
.C(n_21),
.Y(n_1125)
);

NAND4xp25_ASAP7_75t_SL g1126 ( 
.A(n_1123),
.B(n_22),
.C(n_23),
.D(n_24),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_L g1127 ( 
.A(n_1125),
.B(n_24),
.C(n_25),
.Y(n_1127)
);

NOR3xp33_ASAP7_75t_L g1128 ( 
.A(n_1126),
.B(n_26),
.C(n_27),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_SL g1129 ( 
.A(n_1125),
.B(n_26),
.C(n_27),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1129),
.B(n_28),
.Y(n_1130)
);

NAND4xp25_ASAP7_75t_SL g1131 ( 
.A(n_1127),
.B(n_28),
.C(n_29),
.D(n_31),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1128),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1132),
.B(n_29),
.Y(n_1133)
);

AND4x1_ASAP7_75t_L g1134 ( 
.A(n_1130),
.B(n_31),
.C(n_32),
.D(n_405),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_1131),
.B1(n_32),
.B2(n_550),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1133),
.Y(n_1136)
);

NAND4xp75_ASAP7_75t_L g1137 ( 
.A(n_1136),
.B(n_37),
.C(n_40),
.D(n_41),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1135),
.B(n_42),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1138),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1137),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_L g1141 ( 
.A(n_1139),
.B(n_548),
.C(n_44),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1140),
.B(n_46),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_1142),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1141),
.Y(n_1144)
);

NAND5xp2_ASAP7_75t_L g1145 ( 
.A(n_1143),
.B(n_50),
.C(n_51),
.D(n_52),
.E(n_53),
.Y(n_1145)
);

XNOR2x1_ASAP7_75t_L g1146 ( 
.A(n_1144),
.B(n_54),
.Y(n_1146)
);

NAND4xp25_ASAP7_75t_L g1147 ( 
.A(n_1143),
.B(n_55),
.C(n_57),
.D(n_58),
.Y(n_1147)
);

OA22x2_ASAP7_75t_L g1148 ( 
.A1(n_1145),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_1148)
);

XNOR2x1_ASAP7_75t_L g1149 ( 
.A(n_1146),
.B(n_63),
.Y(n_1149)
);

AOI211x1_ASAP7_75t_L g1150 ( 
.A1(n_1147),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1149),
.B(n_1148),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1150),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1151),
.B(n_520),
.C(n_517),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_L g1154 ( 
.A(n_1152),
.B(n_520),
.C(n_517),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1153),
.B(n_69),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1154),
.A2(n_537),
.B1(n_535),
.B2(n_541),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1155),
.A2(n_519),
.B(n_513),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1156),
.A2(n_537),
.B1(n_518),
.B2(n_543),
.Y(n_1158)
);

OAI22x1_ASAP7_75t_SL g1159 ( 
.A1(n_1157),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_SL g1160 ( 
.A1(n_1158),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_1160)
);

OAI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1159),
.A2(n_521),
.B(n_517),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1160),
.A2(n_537),
.B1(n_518),
.B2(n_543),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1159),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1163),
.A2(n_521),
.B(n_520),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1161),
.A2(n_77),
.B(n_78),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1162),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1163),
.B(n_79),
.Y(n_1167)
);

OAI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_1166),
.A2(n_1165),
.B(n_1167),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1164),
.Y(n_1169)
);

XNOR2xp5_ASAP7_75t_L g1170 ( 
.A(n_1166),
.B(n_81),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1166),
.A2(n_521),
.B(n_436),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1169),
.B(n_84),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1168),
.A2(n_436),
.B(n_86),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1170),
.A2(n_426),
.B(n_87),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1171),
.A2(n_547),
.B(n_543),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_1168),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_SL g1177 ( 
.A1(n_1169),
.A2(n_537),
.B1(n_543),
.B2(n_541),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1169),
.Y(n_1178)
);

AOI31xp33_ASAP7_75t_SL g1179 ( 
.A1(n_1169),
.A2(n_85),
.A3(n_92),
.B(n_93),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1169),
.A2(n_547),
.B1(n_541),
.B2(n_539),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_L g1181 ( 
.A(n_1169),
.B(n_94),
.Y(n_1181)
);

XNOR2xp5_ASAP7_75t_L g1182 ( 
.A(n_1169),
.B(n_97),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1168),
.A2(n_547),
.B(n_541),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1178),
.Y(n_1184)
);

OAI222xp33_ASAP7_75t_L g1185 ( 
.A1(n_1176),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.C1(n_101),
.C2(n_103),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1175),
.A2(n_1173),
.B1(n_1181),
.B2(n_1172),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1173),
.A2(n_547),
.B1(n_539),
.B2(n_529),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_1179),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1174),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1182),
.Y(n_1190)
);

OAI222xp33_ASAP7_75t_L g1191 ( 
.A1(n_1183),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.C1(n_109),
.C2(n_111),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1177),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1184),
.A2(n_1190),
.B1(n_1189),
.B2(n_1188),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1192),
.Y(n_1194)
);

NOR2xp67_ASAP7_75t_SL g1195 ( 
.A(n_1186),
.B(n_1187),
.Y(n_1195)
);

XNOR2xp5_ASAP7_75t_L g1196 ( 
.A(n_1191),
.B(n_1180),
.Y(n_1196)
);

AOI222xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1185),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.C1(n_115),
.C2(n_116),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1184),
.A2(n_539),
.B1(n_529),
.B2(n_426),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1184),
.B(n_529),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1193),
.A2(n_118),
.B(n_119),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1194),
.B(n_120),
.Y(n_1201)
);

OAI21xp33_ASAP7_75t_L g1202 ( 
.A1(n_1195),
.A2(n_539),
.B(n_529),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1196),
.A2(n_474),
.B1(n_479),
.B2(n_124),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1199),
.A2(n_479),
.B1(n_404),
.B2(n_546),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1201),
.A2(n_1197),
.B1(n_1198),
.B2(n_125),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1202),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1205),
.A2(n_1200),
.B1(n_1204),
.B2(n_1203),
.Y(n_1207)
);

AOI221xp5_ASAP7_75t_L g1208 ( 
.A1(n_1207),
.A2(n_1206),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_1208)
);

AOI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1208),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_1209)
);

AOI221xp5_ASAP7_75t_L g1210 ( 
.A1(n_1209),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.C(n_145),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1210),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_1211)
);

AOI211xp5_ASAP7_75t_L g1212 ( 
.A1(n_1211),
.A2(n_149),
.B(n_150),
.C(n_152),
.Y(n_1212)
);

AOI211xp5_ASAP7_75t_L g1213 ( 
.A1(n_1212),
.A2(n_154),
.B(n_155),
.C(n_160),
.Y(n_1213)
);


endmodule