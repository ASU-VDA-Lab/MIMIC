module real_jpeg_14587_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_311, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_311;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_3),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_95),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_44),
.B1(n_48),
.B2(n_95),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_95),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_4),
.A2(n_44),
.B1(n_48),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_4),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_141),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_141),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_141),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_7),
.A2(n_44),
.B1(n_48),
.B2(n_61),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_61),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_61),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_8),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_8),
.A2(n_36),
.B1(n_44),
.B2(n_48),
.Y(n_233)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_10),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_10),
.B(n_44),
.C(n_47),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_10),
.B(n_30),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_10),
.A2(n_139),
.B(n_142),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_10),
.A2(n_28),
.B(n_29),
.C(n_170),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_10),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_10),
.B(n_58),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_11),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_44),
.B1(n_48),
.B2(n_136),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_136),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_136),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_12),
.A2(n_39),
.B1(n_44),
.B2(n_48),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_13),
.B(n_27),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_44),
.B1(n_48),
.B2(n_53),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_53),
.Y(n_105)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_16),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_16),
.A2(n_27),
.B1(n_29),
.B2(n_67),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_16),
.A2(n_44),
.B1(n_48),
.B2(n_67),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_67),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_109),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_107),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_96),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_20),
.B(n_96),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_69),
.C(n_77),
.Y(n_20)
);

FAx1_ASAP7_75t_L g306 ( 
.A(n_21),
.B(n_69),
.CI(n_77),
.CON(n_306),
.SN(n_306)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_55),
.B1(n_56),
.B2(n_68),
.Y(n_21)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_40),
.B1(n_41),
.B2(n_54),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_23),
.B(n_41),
.C(n_56),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_23)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_24),
.B(n_177),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_26),
.A2(n_31),
.B(n_124),
.Y(n_170)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g228 ( 
.A1(n_29),
.A2(n_59),
.A3(n_64),
.B1(n_216),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_30),
.B(n_177),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_32),
.B1(n_46),
.B2(n_47),
.Y(n_50)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_32),
.B(n_128),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_35),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_38),
.A2(n_71),
.B1(n_73),
.B2(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_40),
.A2(n_41),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_49),
.B(n_51),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_49),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_42),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_42),
.A2(n_49),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_42),
.A2(n_49),
.B1(n_222),
.B2(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_42),
.A2(n_49),
.B1(n_88),
.B2(n_250),
.Y(n_256)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_52),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_43),
.A2(n_135),
.B(n_137),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_43),
.B(n_124),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_43),
.A2(n_137),
.B(n_221),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_48),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_49),
.B(n_126),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_56),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_63),
.B(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_59),
.A2(n_62),
.B(n_124),
.C(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_62),
.A2(n_63),
.B1(n_243),
.B2(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_62),
.A2(n_263),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_63),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_63),
.B(n_94),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_63),
.A2(n_91),
.B(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_69),
.A2(n_70),
.B(n_74),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_71),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_71),
.A2(n_73),
.B1(n_190),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_71),
.A2(n_176),
.B(n_219),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_265),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_73),
.A2(n_190),
.B(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_73),
.A2(n_191),
.B(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_75),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_75),
.A2(n_125),
.B(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_90),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_78),
.A2(n_79),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_80),
.A2(n_81),
.B1(n_90),
.B2(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_82),
.A2(n_83),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_82),
.B(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_82),
.A2(n_83),
.B1(n_233),
.B2(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_83),
.B(n_143),
.Y(n_142)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_85),
.A2(n_139),
.B1(n_156),
.B2(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_90),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_305),
.B(n_308),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_292),
.B(n_304),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_275),
.B(n_291),
.Y(n_113)
);

OAI321xp33_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_235),
.A3(n_268),
.B1(n_273),
.B2(n_274),
.C(n_311),
.Y(n_114)
);

AOI21x1_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_207),
.B(n_234),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_184),
.B(n_206),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_165),
.B(n_183),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_144),
.B(n_164),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_129),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_122),
.B1(n_127),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_156),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_134),
.C(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B(n_142),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_139),
.A2(n_156),
.B1(n_172),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_139),
.A2(n_156),
.B1(n_198),
.B2(n_232),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_140),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_152),
.B(n_163),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_150),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_148),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_158),
.B(n_162),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_155),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_157),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_178),
.C(n_182),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_171),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_173)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_186),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_199),
.B2(n_200),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_202),
.C(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_193),
.C(n_197),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_209),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_224),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_210),
.B(n_225),
.C(n_226),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_217),
.B2(n_223),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_218),
.C(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_231),
.Y(n_245)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_252),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_252),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_246),
.C(n_251),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_237),
.A2(n_238),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_244),
.C(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_249),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_248),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_267),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_260),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_260),
.C(n_267),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_258),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_266),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_290),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_290),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_288),
.B2(n_289),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_286),
.C(n_289),
.Y(n_303)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_298),
.C(n_303),
.Y(n_307)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_307),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_306),
.Y(n_310)
);


endmodule