module fake_jpeg_25215_n_238 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_238);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_23),
.B1(n_15),
.B2(n_11),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_29),
.B1(n_11),
.B2(n_27),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_22),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_49),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_50),
.B1(n_61),
.B2(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_56),
.B1(n_12),
.B2(n_16),
.Y(n_80)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_60),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_25),
.B1(n_24),
.B2(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_15),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_62),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_37),
.C(n_34),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_69),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_58),
.B1(n_42),
.B2(n_27),
.Y(n_67)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_47),
.B(n_61),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_37),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_74),
.B1(n_77),
.B2(n_80),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_34),
.C(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_61),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_33),
.B1(n_18),
.B2(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_81),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_16),
.Y(n_79)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_47),
.B(n_61),
.C(n_17),
.D(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_56),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_39),
.B1(n_20),
.B2(n_19),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_53),
.B1(n_39),
.B2(n_18),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_75),
.B(n_68),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_41),
.Y(n_126)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_79),
.B(n_22),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_99),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_83),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_59),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_61),
.B(n_10),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_102),
.A2(n_78),
.B(n_9),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_106),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_107),
.B1(n_51),
.B2(n_20),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_53),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_64),
.B(n_53),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_20),
.B1(n_19),
.B2(n_39),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_82),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_112),
.A2(n_119),
.B(n_128),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_66),
.C(n_73),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_125),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_93),
.B(n_95),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_22),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_85),
.A2(n_17),
.B(n_22),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_22),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_131),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_41),
.C(n_51),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_134),
.Y(n_137)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_19),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_94),
.C(n_89),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_99),
.B1(n_86),
.B2(n_106),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_142),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_161),
.B1(n_122),
.B2(n_120),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_84),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_144),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_100),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_84),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_149),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_101),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_89),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_111),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_97),
.B1(n_19),
.B2(n_17),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_112),
.B1(n_135),
.B2(n_120),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

BUFx4f_ASAP7_75t_SL g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_117),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_126),
.C(n_128),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_178),
.C(n_179),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_154),
.B1(n_139),
.B2(n_141),
.Y(n_185)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_113),
.CI(n_134),
.CON(n_167),
.SN(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_155),
.B(n_137),
.C(n_149),
.D(n_158),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_111),
.B1(n_113),
.B2(n_112),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_118),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_173),
.B(n_153),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_130),
.C(n_124),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_117),
.C(n_114),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_147),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_187),
.C(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_170),
.B1(n_168),
.B2(n_171),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_189),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_137),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_194),
.C(n_180),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_158),
.Y(n_190)
);

OA21x2_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_123),
.B(n_154),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_167),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_141),
.C(n_160),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_193),
.A2(n_189),
.B1(n_164),
.B2(n_187),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_181),
.B(n_190),
.C(n_188),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_169),
.B1(n_165),
.B2(n_170),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_202),
.B1(n_172),
.B2(n_51),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_199),
.C(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_201),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_166),
.B(n_163),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_203),
.B(n_206),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_161),
.B1(n_167),
.B2(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_211),
.Y(n_219)
);

BUFx4f_ASAP7_75t_SL g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_182),
.C(n_156),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_213),
.A2(n_198),
.B1(n_205),
.B2(n_200),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_17),
.C(n_10),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_215),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_9),
.C(n_1),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_217),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_9),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_0),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_227),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_0),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_0),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_229),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_222),
.A2(n_218),
.B(n_221),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_217),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_1),
.C2(n_6),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_230),
.A2(n_231),
.B(n_8),
.Y(n_235)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_3),
.C(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_232),
.B(n_235),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_8),
.Y(n_238)
);


endmodule